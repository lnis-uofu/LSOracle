module top(pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 , pi8 , pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 , pi16 , pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 , po0 , po1 , po2 , po3 , po4 , po5 , po6 , po7 , po8 , po9 , po10 , po11 , po12 , po13 , po14 , po15 , po16 , po17 , po18 , po19 , po20 , po21 , po22 , po23 , po24 );
  input pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 , pi8 , pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 , pi16 , pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 ;
  output po0 , po1 , po2 , po3 , po4 , po5 , po6 , po7 , po8 , po9 , po10 , po11 , po12 , po13 , po14 , po15 , po16 , po17 , po18 , po19 , po20 , po21 , po22 , po23 , po24 ;
  wire n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517;
  assign n25 = pi0 | pi1 ;
  assign n26 = ~pi22 & n25 ;
  assign n27 = ~pi2 & n26 ;
  assign n28 = pi2 & ~n26 ;
  assign n29 = n27 | n28 ;
  assign n30 = pi5 | pi8 ;
  assign n31 = pi7 | pi10 ;
  assign n32 = pi4 | pi6 ;
  assign n33 = n31 | n32 ;
  assign n34 = n30 | n33 ;
  assign n35 = pi2 | n25 ;
  assign n36 = pi3 | n35 ;
  assign n37 = pi9 | n36 ;
  assign n38 = pi11 | pi12 ;
  assign n39 = n37 | n38 ;
  assign n40 = n34 | n39 ;
  assign n41 = ~pi22 & n40 ;
  assign n42 = pi13 & ~n41 ;
  assign n43 = ~pi13 & n41 ;
  assign n44 = n42 | n43 ;
  assign n45 = pi13 | n40 ;
  assign n46 = pi14 | n45 ;
  assign n47 = ~pi22 & n46 ;
  assign n48 = ~pi15 & n47 ;
  assign n49 = pi15 & ~n47 ;
  assign n50 = n48 | n49 ;
  assign n51 = pi17 | n46 ;
  assign n52 = pi16 | n51 ;
  assign n53 = pi15 | pi18 ;
  assign n54 = pi19 | n53 ;
  assign n55 = n52 | n54 ;
  assign n56 = ~pi22 & n55 ;
  assign n57 = ~pi20 & n56 ;
  assign n58 = pi20 & ~n56 ;
  assign n59 = n57 | n58 ;
  assign n60 = pi16 | pi20 ;
  assign n61 = n51 | n60 ;
  assign n62 = n54 | n61 ;
  assign n63 = ~pi22 & n62 ;
  assign n64 = ~pi21 & n63 ;
  assign n65 = pi21 & ~n63 ;
  assign n66 = n64 | n65 ;
  assign n67 = n59 & n66 ;
  assign n68 = n50 & n67 ;
  assign n69 = ~n50 & n67 ;
  assign n70 = n68 | n69 ;
  assign n71 = pi16 | n46 ;
  assign n72 = pi15 | pi17 ;
  assign n73 = n71 | n72 ;
  assign n74 = ~pi22 & n73 ;
  assign n75 = ~pi18 & n74 ;
  assign n76 = pi18 & ~n74 ;
  assign n77 = n75 | n76 ;
  assign n78 = pi18 | n73 ;
  assign n79 = ~pi22 & n78 ;
  assign n80 = pi19 & ~n79 ;
  assign n81 = pi19 | pi22 ;
  assign n82 = n78 & ~n81 ;
  assign n83 = n80 | n82 ;
  assign n84 = n77 & n83 ;
  assign n85 = pi15 | n46 ;
  assign n86 = ~pi22 & n85 ;
  assign n87 = pi16 & ~n86 ;
  assign n88 = ~pi16 & n86 ;
  assign n89 = n87 | n88 ;
  assign n90 = pi16 | n85 ;
  assign n91 = ~pi22 & n90 ;
  assign n92 = pi17 & ~n91 ;
  assign n93 = ~pi17 & n91 ;
  assign n94 = n92 | n93 ;
  assign n95 = n89 & n94 ;
  assign n96 = n84 & n95 ;
  assign n97 = ~n89 & n94 ;
  assign n98 = n77 | n83 ;
  assign n99 = n97 & ~n98 ;
  assign n100 = n96 | n99 ;
  assign n101 = n70 & n100 ;
  assign n102 = n84 & n97 ;
  assign n103 = n69 & n102 ;
  assign n104 = n77 & ~n83 ;
  assign n105 = n95 & n104 ;
  assign n106 = n68 & n105 ;
  assign n107 = n89 | n94 ;
  assign n108 = ~n77 & n83 ;
  assign n109 = ~n107 & n108 ;
  assign n110 = ~n59 & n66 ;
  assign n111 = ~n50 & n110 ;
  assign n112 = n109 & n111 ;
  assign n113 = n50 & n110 ;
  assign n114 = n109 & n113 ;
  assign n115 = n112 | n114 ;
  assign n116 = n106 | n115 ;
  assign n117 = n104 & ~n107 ;
  assign n118 = n68 & n117 ;
  assign n119 = n69 & n105 ;
  assign n120 = n97 & n104 ;
  assign n121 = n68 & n120 ;
  assign n122 = n119 | n121 ;
  assign n123 = n89 & ~n94 ;
  assign n124 = n108 & n123 ;
  assign n125 = n111 & n124 ;
  assign n126 = n69 & n117 ;
  assign n127 = n125 | n126 ;
  assign n128 = n122 | n127 ;
  assign n129 = n118 | n128 ;
  assign n130 = n116 | n129 ;
  assign n131 = n103 | n130 ;
  assign n132 = n96 & n113 ;
  assign n133 = n98 | n107 ;
  assign n134 = n69 & ~n133 ;
  assign n135 = n132 | n134 ;
  assign n136 = n95 & ~n98 ;
  assign n137 = n68 & n136 ;
  assign n138 = n84 & n123 ;
  assign n139 = n113 & n138 ;
  assign n140 = n137 | n139 ;
  assign n141 = n97 & n108 ;
  assign n142 = n68 & n141 ;
  assign n143 = n69 & n141 ;
  assign n144 = n95 & n108 ;
  assign n145 = n69 & n144 ;
  assign n146 = n143 | n145 ;
  assign n147 = n84 & ~n107 ;
  assign n148 = n113 & n147 ;
  assign n149 = n69 & n136 ;
  assign n150 = n148 | n149 ;
  assign n151 = n146 | n150 ;
  assign n152 = n142 | n151 ;
  assign n153 = n140 | n152 ;
  assign n154 = n111 & n147 ;
  assign n155 = n111 & n138 ;
  assign n156 = n154 | n155 ;
  assign n157 = n153 | n156 ;
  assign n158 = n135 | n157 ;
  assign n159 = n131 | n158 ;
  assign n160 = n69 & n138 ;
  assign n161 = n113 & n124 ;
  assign n162 = n68 & n124 ;
  assign n163 = n161 | n162 ;
  assign n164 = n68 & ~n133 ;
  assign n165 = n68 & n138 ;
  assign n166 = ~n98 & n123 ;
  assign n167 = n69 & n166 ;
  assign n168 = n165 | n167 ;
  assign n169 = n164 | n168 ;
  assign n170 = n163 | n169 ;
  assign n171 = n160 | n170 ;
  assign n172 = n159 | n171 ;
  assign n173 = n68 & n102 ;
  assign n174 = n68 & n166 ;
  assign n175 = n173 | n174 ;
  assign n176 = n68 & n144 ;
  assign n177 = n102 & n113 ;
  assign n178 = n69 & n147 ;
  assign n179 = n177 | n178 ;
  assign n180 = n176 | n179 ;
  assign n181 = n96 & n111 ;
  assign n182 = n68 & n147 ;
  assign n183 = n102 & n111 ;
  assign n184 = n182 | n183 ;
  assign n185 = n181 | n184 ;
  assign n186 = n180 | n185 ;
  assign n187 = n113 & n144 ;
  assign n188 = n113 & n141 ;
  assign n189 = n111 & n141 ;
  assign n190 = n188 | n189 ;
  assign n191 = n68 & n109 ;
  assign n192 = n111 & n144 ;
  assign n193 = n69 & n109 ;
  assign n194 = n192 | n193 ;
  assign n195 = n191 | n194 ;
  assign n196 = n190 | n195 ;
  assign n197 = n113 & n120 ;
  assign n198 = n105 & n111 ;
  assign n199 = n197 | n198 ;
  assign n200 = n104 & n123 ;
  assign n201 = n68 & n200 ;
  assign n202 = n105 & n113 ;
  assign n203 = n201 | n202 ;
  assign n204 = n69 & n200 ;
  assign n205 = n69 & n124 ;
  assign n206 = n69 & n120 ;
  assign n207 = n205 | n206 ;
  assign n208 = n204 | n207 ;
  assign n209 = n203 | n208 ;
  assign n210 = n199 | n209 ;
  assign n211 = n196 | n210 ;
  assign n212 = n187 | n211 ;
  assign n213 = n186 | n212 ;
  assign n214 = n175 | n213 ;
  assign n215 = n172 | n214 ;
  assign n216 = n101 | n215 ;
  assign n217 = n44 & n216 ;
  assign n218 = ~pi22 & n45 ;
  assign n219 = ~pi14 & n218 ;
  assign n220 = pi14 & ~n218 ;
  assign n221 = n219 | n220 ;
  assign n222 = n59 | n66 ;
  assign n223 = n50 & ~n222 ;
  assign n224 = n124 & n223 ;
  assign n225 = n50 | n222 ;
  assign n226 = n144 & ~n225 ;
  assign n227 = n141 & n223 ;
  assign n228 = n226 | n227 ;
  assign n229 = n141 & ~n225 ;
  assign n230 = n144 & n223 ;
  assign n231 = n124 & ~n225 ;
  assign n232 = n230 | n231 ;
  assign n233 = n229 | n232 ;
  assign n234 = n228 | n233 ;
  assign n235 = n147 & ~n225 ;
  assign n236 = n96 & n223 ;
  assign n237 = n102 & n223 ;
  assign n238 = n59 & ~n66 ;
  assign n239 = ~n50 & n238 ;
  assign n240 = ~n133 & n239 ;
  assign n241 = n237 | n240 ;
  assign n242 = n50 & n238 ;
  assign n243 = ~n133 & n242 ;
  assign n244 = n113 & n117 ;
  assign n245 = n113 & n200 ;
  assign n246 = n244 | n245 ;
  assign n247 = n243 | n246 ;
  assign n248 = n147 & n223 ;
  assign n249 = n138 & n223 ;
  assign n250 = n248 | n249 ;
  assign n251 = n247 | n250 ;
  assign n252 = n102 & ~n225 ;
  assign n253 = n111 & n117 ;
  assign n254 = n111 & n200 ;
  assign n255 = n253 | n254 ;
  assign n256 = n252 | n255 ;
  assign n257 = n251 | n256 ;
  assign n258 = n241 | n257 ;
  assign n259 = n236 | n258 ;
  assign n260 = n96 & ~n225 ;
  assign n261 = n138 & ~n225 ;
  assign n262 = n260 | n261 ;
  assign n263 = n259 | n262 ;
  assign n264 = n235 | n263 ;
  assign n265 = n109 & n223 ;
  assign n266 = n147 & n239 ;
  assign n267 = n144 & n242 ;
  assign n268 = n144 & n239 ;
  assign n269 = n267 | n268 ;
  assign n270 = n102 & n242 ;
  assign n271 = n138 & n239 ;
  assign n272 = n147 & n242 ;
  assign n273 = n138 & n242 ;
  assign n274 = n272 | n273 ;
  assign n275 = n271 | n274 ;
  assign n276 = n270 | n275 ;
  assign n277 = n269 | n276 ;
  assign n278 = n141 & n242 ;
  assign n279 = n111 & n166 ;
  assign n280 = n278 | n279 ;
  assign n281 = n96 & n242 ;
  assign n282 = n102 & n239 ;
  assign n283 = n111 & n136 ;
  assign n284 = n282 | n283 ;
  assign n285 = n281 | n284 ;
  assign n286 = n280 | n285 ;
  assign n287 = n99 & n113 ;
  assign n288 = n113 & n166 ;
  assign n289 = n287 | n288 ;
  assign n290 = n96 & n239 ;
  assign n291 = n111 & n120 ;
  assign n292 = n290 | n291 ;
  assign n293 = n99 & n111 ;
  assign n294 = n113 & n136 ;
  assign n295 = n293 | n294 ;
  assign n296 = n292 | n295 ;
  assign n297 = n289 | n296 ;
  assign n298 = n286 | n297 ;
  assign n299 = n277 | n298 ;
  assign n300 = n266 | n299 ;
  assign n301 = n111 & ~n133 ;
  assign n302 = n113 & ~n133 ;
  assign n303 = n301 | n302 ;
  assign n304 = n300 | n303 ;
  assign n305 = n265 | n304 ;
  assign n306 = n264 | n305 ;
  assign n307 = n234 | n306 ;
  assign n308 = n224 | n307 ;
  assign n309 = n200 & n239 ;
  assign n310 = n136 & n242 ;
  assign n311 = n117 & n239 ;
  assign n312 = n310 | n311 ;
  assign n313 = n99 & n242 ;
  assign n314 = n166 & n242 ;
  assign n315 = n99 & n239 ;
  assign n316 = n136 & n239 ;
  assign n317 = n117 & n242 ;
  assign n318 = n166 & n239 ;
  assign n319 = n317 | n318 ;
  assign n320 = n316 | n319 ;
  assign n321 = n315 | n320 ;
  assign n322 = n314 | n321 ;
  assign n323 = n313 | n322 ;
  assign n324 = n312 | n323 ;
  assign n325 = n109 & n242 ;
  assign n326 = n200 & n242 ;
  assign n327 = n105 & n239 ;
  assign n328 = n120 & n239 ;
  assign n329 = n327 | n328 ;
  assign n330 = n326 | n329 ;
  assign n331 = n120 & n242 ;
  assign n332 = n105 & n242 ;
  assign n333 = n141 & n239 ;
  assign n334 = n332 | n333 ;
  assign n335 = n331 | n334 ;
  assign n336 = n330 | n335 ;
  assign n337 = n325 | n336 ;
  assign n338 = n124 & n242 ;
  assign n339 = n109 & n239 ;
  assign n340 = n124 & n239 ;
  assign n341 = n339 | n340 ;
  assign n342 = n338 | n341 ;
  assign n343 = n337 | n342 ;
  assign n344 = n246 | n343 ;
  assign n345 = n304 | n344 ;
  assign n346 = n255 | n345 ;
  assign n347 = n324 | n346 ;
  assign n348 = n309 | n347 ;
  assign n349 = n308 & n348 ;
  assign n350 = n216 & ~n349 ;
  assign n351 = n221 | n350 ;
  assign n352 = ~n308 & n348 ;
  assign n353 = n308 & ~n348 ;
  assign n354 = n352 | n353 ;
  assign n355 = ~n350 & n354 ;
  assign n356 = n308 | n348 ;
  assign n357 = ~n216 & n356 ;
  assign n358 = n354 | n357 ;
  assign n359 = n221 & ~n358 ;
  assign n360 = n355 | n359 ;
  assign n361 = n351 & ~n360 ;
  assign n362 = ~n217 & n361 ;
  assign n363 = pi8 | pi10 ;
  assign n364 = pi4 | pi5 ;
  assign n365 = n363 | n364 ;
  assign n366 = pi6 | pi7 ;
  assign n367 = n37 | n366 ;
  assign n368 = n365 | n367 ;
  assign n369 = ~pi22 & n368 ;
  assign n370 = pi11 & ~n369 ;
  assign n371 = ~pi11 & n369 ;
  assign n372 = n370 | n371 ;
  assign n373 = n216 & n372 ;
  assign n374 = n105 & ~n225 ;
  assign n375 = n294 | n326 ;
  assign n376 = n374 | n375 ;
  assign n377 = n178 | n253 ;
  assign n378 = n261 | n301 ;
  assign n379 = n200 & n223 ;
  assign n380 = n117 & ~n225 ;
  assign n381 = n302 | n380 ;
  assign n382 = n244 | n381 ;
  assign n383 = n164 | n204 ;
  assign n384 = n106 | n338 ;
  assign n385 = n383 | n384 ;
  assign n386 = n120 & ~n225 ;
  assign n387 = n325 | n386 ;
  assign n388 = n243 | n328 ;
  assign n389 = n117 & n223 ;
  assign n390 = n252 | n389 ;
  assign n391 = n207 | n390 ;
  assign n392 = n121 | n162 ;
  assign n393 = n391 | n392 ;
  assign n394 = n388 | n393 ;
  assign n395 = n387 | n394 ;
  assign n396 = n68 & n96 ;
  assign n397 = n109 & ~n225 ;
  assign n398 = n200 & ~n225 ;
  assign n399 = n146 | n334 ;
  assign n400 = n105 & n223 ;
  assign n401 = n241 | n254 ;
  assign n402 = n68 & n99 ;
  assign n403 = n118 | n402 ;
  assign n404 = n176 | n403 ;
  assign n405 = n401 | n404 ;
  assign n406 = n400 | n405 ;
  assign n407 = n291 | n406 ;
  assign n408 = n399 | n407 ;
  assign n409 = n245 | n408 ;
  assign n410 = n103 | n149 ;
  assign n411 = n126 | n410 ;
  assign n412 = n175 | n327 ;
  assign n413 = n411 | n412 ;
  assign n414 = n409 | n413 ;
  assign n415 = n398 | n414 ;
  assign n416 = n397 | n415 ;
  assign n417 = n396 | n416 ;
  assign n418 = n395 | n417 ;
  assign n419 = n248 | n283 ;
  assign n420 = n193 | n339 ;
  assign n421 = n167 | n420 ;
  assign n422 = n419 | n421 ;
  assign n423 = n418 | n422 ;
  assign n424 = n385 | n423 ;
  assign n425 = n382 | n424 ;
  assign n426 = n379 | n425 ;
  assign n427 = n378 | n426 ;
  assign n428 = n377 | n427 ;
  assign n429 = n182 | n287 ;
  assign n430 = n69 & n96 ;
  assign n431 = n134 | n181 ;
  assign n432 = n165 | n340 ;
  assign n433 = n431 | n432 ;
  assign n434 = n430 | n433 ;
  assign n435 = n331 | n434 ;
  assign n436 = n429 | n435 ;
  assign n437 = n137 | n288 ;
  assign n438 = n119 | n191 ;
  assign n439 = n249 | n438 ;
  assign n440 = n437 | n439 ;
  assign n441 = n132 | n279 ;
  assign n442 = n160 | n441 ;
  assign n443 = n236 | n442 ;
  assign n444 = n120 & n223 ;
  assign n445 = n69 & n99 ;
  assign n446 = n142 | n293 ;
  assign n447 = n445 | n446 ;
  assign n448 = n444 | n447 ;
  assign n449 = n201 | n448 ;
  assign n450 = n443 | n449 ;
  assign n451 = n440 | n450 ;
  assign n452 = n436 | n451 ;
  assign n453 = n428 | n452 ;
  assign n454 = n376 | n453 ;
  assign n455 = n260 | n454 ;
  assign n456 = n183 | n245 ;
  assign n457 = n188 | n397 ;
  assign n458 = n333 | n457 ;
  assign n459 = n456 | n458 ;
  assign n460 = n254 | n283 ;
  assign n461 = n154 | n273 ;
  assign n462 = n460 | n461 ;
  assign n463 = n270 | n309 ;
  assign n464 = n162 | n463 ;
  assign n465 = n207 | n444 ;
  assign n466 = n464 | n465 ;
  assign n467 = n146 | n160 ;
  assign n468 = n119 | n173 ;
  assign n469 = n467 | n468 ;
  assign n470 = n177 | n282 ;
  assign n471 = n106 | n400 ;
  assign n472 = n470 | n471 ;
  assign n473 = n469 | n472 ;
  assign n474 = n466 | n473 ;
  assign n475 = n311 | n474 ;
  assign n476 = n191 | n475 ;
  assign n477 = n290 | n325 ;
  assign n478 = n240 | n477 ;
  assign n479 = n476 | n478 ;
  assign n480 = n136 & ~n225 ;
  assign n481 = n148 | n480 ;
  assign n482 = n479 | n481 ;
  assign n483 = n317 | n430 ;
  assign n484 = n341 | n483 ;
  assign n485 = n227 | n484 ;
  assign n486 = n281 | n294 ;
  assign n487 = n121 | n187 ;
  assign n488 = n244 | n487 ;
  assign n489 = n193 | n488 ;
  assign n490 = n235 | n489 ;
  assign n491 = n486 | n490 ;
  assign n492 = n485 | n491 ;
  assign n493 = n482 | n492 ;
  assign n494 = n462 | n493 ;
  assign n495 = n459 | n494 ;
  assign n496 = n99 & ~n225 ;
  assign n497 = n139 | n230 ;
  assign n498 = n155 | n497 ;
  assign n499 = n201 | n260 ;
  assign n500 = n99 & n223 ;
  assign n501 = n386 | n500 ;
  assign n502 = n204 | n501 ;
  assign n503 = n499 | n502 ;
  assign n504 = n243 | n338 ;
  assign n505 = n165 | n182 ;
  assign n506 = n192 | n505 ;
  assign n507 = n377 | n506 ;
  assign n508 = n226 | n507 ;
  assign n509 = n504 | n508 ;
  assign n510 = n136 & n223 ;
  assign n511 = n236 | n310 ;
  assign n512 = n510 | n511 ;
  assign n513 = n142 | n396 ;
  assign n514 = n176 | n513 ;
  assign n515 = n512 | n514 ;
  assign n516 = n509 | n515 ;
  assign n517 = n503 | n516 ;
  assign n518 = n498 | n517 ;
  assign n519 = n496 | n518 ;
  assign n520 = n103 | n291 ;
  assign n521 = n519 | n520 ;
  assign n522 = n374 | n521 ;
  assign n523 = n495 | n522 ;
  assign n524 = n455 & n523 ;
  assign n525 = n308 & ~n524 ;
  assign n526 = n373 & ~n525 ;
  assign n527 = ~n373 & n525 ;
  assign n528 = n526 | n527 ;
  assign n529 = pi11 & ~pi22 ;
  assign n530 = n369 | n529 ;
  assign n531 = pi12 & n530 ;
  assign n532 = pi12 | n529 ;
  assign n533 = n369 | n532 ;
  assign n534 = ~n531 & n533 ;
  assign n535 = n216 & n534 ;
  assign n536 = ~n528 & n535 ;
  assign n537 = n526 | n536 ;
  assign n538 = n217 & ~n361 ;
  assign n539 = n362 | n538 ;
  assign n540 = n537 & ~n539 ;
  assign n541 = n362 | n540 ;
  assign n542 = n455 & ~n523 ;
  assign n543 = ~n455 & n523 ;
  assign n544 = n542 | n543 ;
  assign n545 = n221 & ~n544 ;
  assign n546 = n525 | n545 ;
  assign n547 = n455 | n523 ;
  assign n548 = ~n308 & n547 ;
  assign n549 = n545 & ~n548 ;
  assign n550 = n546 & ~n549 ;
  assign n551 = ~n373 & n550 ;
  assign n552 = n373 & ~n550 ;
  assign n553 = n551 | n552 ;
  assign n554 = n350 | n354 ;
  assign n555 = n534 | n554 ;
  assign n556 = ~n358 & n533 ;
  assign n557 = ~n531 & n556 ;
  assign n558 = n555 & ~n557 ;
  assign n559 = n354 & ~n357 ;
  assign n560 = n44 & n559 ;
  assign n561 = ~n44 & n355 ;
  assign n562 = n560 | n561 ;
  assign n563 = n558 & ~n562 ;
  assign n564 = ~n553 & n563 ;
  assign n565 = n551 | n564 ;
  assign n566 = n221 & n559 ;
  assign n567 = ~n220 & n355 ;
  assign n568 = ~n219 & n567 ;
  assign n569 = n44 & ~n358 ;
  assign n570 = n44 | n554 ;
  assign n571 = ~n569 & n570 ;
  assign n572 = ~n568 & n571 ;
  assign n573 = ~n566 & n572 ;
  assign n574 = n565 & n573 ;
  assign n575 = n565 | n573 ;
  assign n576 = ~n574 & n575 ;
  assign n577 = n528 & ~n535 ;
  assign n578 = n536 | n577 ;
  assign n579 = n576 & ~n578 ;
  assign n580 = n574 | n579 ;
  assign n581 = ~n537 & n539 ;
  assign n582 = n540 | n581 ;
  assign n583 = n580 & ~n582 ;
  assign n584 = n166 & n223 ;
  assign n585 = n230 | n584 ;
  assign n586 = n142 | n178 ;
  assign n587 = n165 | n235 ;
  assign n588 = n266 | n587 ;
  assign n589 = n586 | n588 ;
  assign n590 = n137 | n252 ;
  assign n591 = n148 | n590 ;
  assign n592 = n162 | n591 ;
  assign n593 = n589 | n592 ;
  assign n594 = n224 | n338 ;
  assign n595 = n155 | n594 ;
  assign n596 = n445 | n595 ;
  assign n597 = n281 | n290 ;
  assign n598 = n189 | n597 ;
  assign n599 = n293 | n598 ;
  assign n600 = n596 | n599 ;
  assign n601 = n593 | n600 ;
  assign n602 = n177 | n316 ;
  assign n603 = n601 | n602 ;
  assign n604 = n161 | n182 ;
  assign n605 = n603 | n604 ;
  assign n606 = n315 | n317 ;
  assign n607 = n430 | n606 ;
  assign n608 = n605 | n607 ;
  assign n609 = n271 | n510 ;
  assign n610 = n183 | n609 ;
  assign n611 = n249 | n610 ;
  assign n612 = n243 | n611 ;
  assign n613 = n114 | n160 ;
  assign n614 = n125 | n139 ;
  assign n615 = n613 | n614 ;
  assign n616 = n229 | n463 ;
  assign n617 = n287 | n379 ;
  assign n618 = n166 & ~n225 ;
  assign n619 = n288 | n480 ;
  assign n620 = n618 | n619 ;
  assign n621 = n617 | n620 ;
  assign n622 = n616 | n621 ;
  assign n623 = n313 | n622 ;
  assign n624 = n272 | n623 ;
  assign n625 = n417 | n624 ;
  assign n626 = n615 | n625 ;
  assign n627 = n612 | n626 ;
  assign n628 = n608 | n627 ;
  assign n629 = n585 | n628 ;
  assign n630 = n205 | n272 ;
  assign n631 = n332 | n630 ;
  assign n632 = n161 | n584 ;
  assign n633 = n187 | n632 ;
  assign n634 = n333 | n633 ;
  assign n635 = n247 | n634 ;
  assign n636 = n252 | n635 ;
  assign n637 = n237 | n636 ;
  assign n638 = n631 | n637 ;
  assign n639 = n193 | n314 ;
  assign n640 = n328 | n340 ;
  assign n641 = n639 | n640 ;
  assign n642 = n397 | n641 ;
  assign n643 = n313 | n500 ;
  assign n644 = n642 | n643 ;
  assign n645 = n638 | n644 ;
  assign n646 = n183 | n645 ;
  assign n647 = n139 | n287 ;
  assign n648 = n279 | n647 ;
  assign n649 = n646 | n648 ;
  assign n650 = ~n133 & n223 ;
  assign n651 = n137 | n311 ;
  assign n652 = n271 | n651 ;
  assign n653 = n134 | n167 ;
  assign n654 = n652 | n653 ;
  assign n655 = n229 | n654 ;
  assign n656 = n650 | n655 ;
  assign n657 = n235 | n656 ;
  assign n658 = n126 | n657 ;
  assign n659 = n261 | n281 ;
  assign n660 = n231 | n659 ;
  assign n661 = n309 | n325 ;
  assign n662 = n112 | n189 ;
  assign n663 = n661 | n662 ;
  assign n664 = n660 | n663 ;
  assign n665 = n374 | n664 ;
  assign n666 = n658 | n665 ;
  assign n667 = n379 | n389 ;
  assign n668 = n253 | n667 ;
  assign n669 = n149 | n668 ;
  assign n670 = n154 | n291 ;
  assign n671 = n438 | n670 ;
  assign n672 = n444 | n671 ;
  assign n673 = n669 | n672 ;
  assign n674 = n666 | n673 ;
  assign n675 = n106 | n226 ;
  assign n676 = n267 | n316 ;
  assign n677 = n202 | n676 ;
  assign n678 = n675 | n677 ;
  assign n679 = n236 | n678 ;
  assign n680 = n118 | n164 ;
  assign n681 = n331 | n680 ;
  assign n682 = n679 | n681 ;
  assign n683 = n470 | n682 ;
  assign n684 = n674 | n683 ;
  assign n685 = n649 | n684 ;
  assign n686 = n510 | n685 ;
  assign n687 = n629 & n686 ;
  assign n688 = n523 & ~n687 ;
  assign n689 = pi4 | n36 ;
  assign n690 = pi5 | n689 ;
  assign n691 = n366 | n690 ;
  assign n692 = pi8 | n691 ;
  assign n693 = ~pi22 & n692 ;
  assign n694 = pi9 & ~n693 ;
  assign n695 = ~pi9 & n693 ;
  assign n696 = n694 | n695 ;
  assign n697 = n216 & n696 ;
  assign n698 = ~n688 & n697 ;
  assign n699 = n688 & ~n697 ;
  assign n700 = n698 | n699 ;
  assign n701 = pi9 | n692 ;
  assign n702 = ~pi22 & n701 ;
  assign n703 = ~pi10 & n702 ;
  assign n704 = pi10 & ~n702 ;
  assign n705 = n703 | n704 ;
  assign n706 = n216 & n705 ;
  assign n707 = ~n700 & n706 ;
  assign n708 = n698 | n707 ;
  assign n709 = n355 & ~n534 ;
  assign n710 = n372 | n554 ;
  assign n711 = n534 & n559 ;
  assign n712 = ~n358 & n372 ;
  assign n713 = n711 | n712 ;
  assign n714 = n710 & ~n713 ;
  assign n715 = ~n709 & n714 ;
  assign n716 = n544 & ~n548 ;
  assign n717 = n221 & n716 ;
  assign n718 = n544 | n548 ;
  assign n719 = n44 & ~n718 ;
  assign n720 = n525 | n544 ;
  assign n721 = n44 | n720 ;
  assign n722 = ~n525 & n544 ;
  assign n723 = ~n221 & n722 ;
  assign n724 = n721 & ~n723 ;
  assign n725 = ~n719 & n724 ;
  assign n726 = ~n717 & n725 ;
  assign n727 = n715 & n726 ;
  assign n728 = n629 & ~n686 ;
  assign n729 = ~n629 & n686 ;
  assign n730 = n728 | n729 ;
  assign n731 = n221 & ~n730 ;
  assign n732 = n688 | n731 ;
  assign n733 = n629 | n686 ;
  assign n734 = ~n523 & n733 ;
  assign n735 = n731 & ~n734 ;
  assign n736 = n732 & ~n735 ;
  assign n737 = ~n697 & n736 ;
  assign n738 = n697 & ~n736 ;
  assign n739 = n737 | n738 ;
  assign n740 = n44 & n716 ;
  assign n741 = n534 & ~n718 ;
  assign n742 = n534 | n720 ;
  assign n743 = ~n44 & n722 ;
  assign n744 = n742 & ~n743 ;
  assign n745 = ~n741 & n744 ;
  assign n746 = ~n740 & n745 ;
  assign n747 = ~n739 & n746 ;
  assign n748 = n737 | n747 ;
  assign n749 = n715 | n726 ;
  assign n750 = ~n727 & n749 ;
  assign n751 = n748 & n750 ;
  assign n752 = n727 | n751 ;
  assign n753 = n708 & n752 ;
  assign n754 = n553 & ~n563 ;
  assign n755 = n564 | n754 ;
  assign n756 = n708 | n752 ;
  assign n757 = ~n753 & n756 ;
  assign n758 = ~n755 & n757 ;
  assign n759 = n753 | n758 ;
  assign n760 = ~n576 & n578 ;
  assign n761 = n579 | n760 ;
  assign n762 = n759 & ~n761 ;
  assign n763 = ~n759 & n761 ;
  assign n764 = n762 | n763 ;
  assign n765 = n755 & ~n757 ;
  assign n766 = n758 | n765 ;
  assign n767 = n372 & n559 ;
  assign n768 = n355 & ~n372 ;
  assign n769 = n554 | n705 ;
  assign n770 = ~n358 & n705 ;
  assign n771 = n769 & ~n770 ;
  assign n772 = ~n768 & n771 ;
  assign n773 = ~n767 & n772 ;
  assign n774 = ~pi22 & n690 ;
  assign n775 = pi6 & ~pi22 ;
  assign n776 = n774 | n775 ;
  assign n777 = ~pi7 & n776 ;
  assign n778 = pi7 & ~n776 ;
  assign n779 = n777 | n778 ;
  assign n780 = n216 & n779 ;
  assign n781 = n125 | n137 ;
  assign n782 = n260 | n480 ;
  assign n783 = n116 | n142 ;
  assign n784 = n333 | n783 ;
  assign n785 = n265 | n293 ;
  assign n786 = n231 | n290 ;
  assign n787 = n785 | n786 ;
  assign n788 = n784 | n787 ;
  assign n789 = n782 | n788 ;
  assign n790 = n198 | n205 ;
  assign n791 = n432 | n790 ;
  assign n792 = n512 | n791 ;
  assign n793 = n789 | n792 ;
  assign n794 = n309 | n793 ;
  assign n795 = n781 | n794 ;
  assign n796 = n496 | n618 ;
  assign n797 = n189 | n650 ;
  assign n798 = n192 | n235 ;
  assign n799 = n167 | n798 ;
  assign n800 = n797 | n799 ;
  assign n801 = n316 | n339 ;
  assign n802 = n103 | n402 ;
  assign n803 = n197 | n802 ;
  assign n804 = n181 | n803 ;
  assign n805 = n281 | n804 ;
  assign n806 = n203 | n805 ;
  assign n807 = n801 | n806 ;
  assign n808 = n374 | n500 ;
  assign n809 = n271 | n302 ;
  assign n810 = n160 | n282 ;
  assign n811 = n809 | n810 ;
  assign n812 = n230 | n811 ;
  assign n813 = n266 | n331 ;
  assign n814 = n812 | n813 ;
  assign n815 = n808 | n814 ;
  assign n816 = n807 | n815 ;
  assign n817 = n800 | n816 ;
  assign n818 = n400 | n817 ;
  assign n819 = n148 | n430 ;
  assign n820 = n332 | n819 ;
  assign n821 = n818 | n820 ;
  assign n822 = n145 | n821 ;
  assign n823 = n314 | n822 ;
  assign n824 = n133 | n225 ;
  assign n825 = ~n161 & n824 ;
  assign n826 = n268 | n396 ;
  assign n827 = n237 | n826 ;
  assign n828 = n319 | n488 ;
  assign n829 = n173 | n397 ;
  assign n830 = n118 | n829 ;
  assign n831 = n828 | n830 ;
  assign n832 = n827 | n831 ;
  assign n833 = n825 & ~n832 ;
  assign n834 = ~n287 & n833 ;
  assign n835 = n164 | n253 ;
  assign n836 = n154 | n835 ;
  assign n837 = n177 | n188 ;
  assign n838 = n584 | n837 ;
  assign n839 = n836 | n838 ;
  assign n840 = n248 | n839 ;
  assign n841 = n834 & ~n840 ;
  assign n842 = ~n823 & n841 ;
  assign n843 = ~n796 & n842 ;
  assign n844 = ~n795 & n843 ;
  assign n845 = ~n132 & n844 ;
  assign n846 = n294 | n338 ;
  assign n847 = n267 | n846 ;
  assign n848 = n311 | n327 ;
  assign n849 = n154 | n173 ;
  assign n850 = n189 | n310 ;
  assign n851 = n849 | n850 ;
  assign n852 = n848 | n851 ;
  assign n853 = n847 | n852 ;
  assign n854 = n340 | n407 ;
  assign n855 = n268 | n331 ;
  assign n856 = n192 | n855 ;
  assign n857 = n226 | n856 ;
  assign n858 = n244 | n857 ;
  assign n859 = n126 | n167 ;
  assign n860 = n396 | n859 ;
  assign n861 = n155 | n191 ;
  assign n862 = n860 | n861 ;
  assign n863 = n243 | n862 ;
  assign n864 = n858 | n863 ;
  assign n865 = n103 | n430 ;
  assign n866 = n178 | n273 ;
  assign n867 = n865 | n866 ;
  assign n868 = n193 | n867 ;
  assign n869 = n183 | n374 ;
  assign n870 = n868 | n869 ;
  assign n871 = n864 | n870 ;
  assign n872 = n182 | n445 ;
  assign n873 = n207 | n872 ;
  assign n874 = n397 | n441 ;
  assign n875 = n121 | n165 ;
  assign n876 = n224 | n271 ;
  assign n877 = n875 | n876 ;
  assign n878 = n787 | n877 ;
  assign n879 = n874 | n878 ;
  assign n880 = n873 | n879 ;
  assign n881 = n871 | n880 ;
  assign n882 = n227 | n236 ;
  assign n883 = n112 | n177 ;
  assign n884 = n229 | n883 ;
  assign n885 = n302 | n884 ;
  assign n886 = n160 | n198 ;
  assign n887 = n885 | n886 ;
  assign n888 = n882 | n887 ;
  assign n889 = n316 | n888 ;
  assign n890 = n881 | n889 ;
  assign n891 = n854 | n890 ;
  assign n892 = n125 | n260 ;
  assign n893 = n891 | n892 ;
  assign n894 = n853 | n893 ;
  assign n895 = ~n845 & n894 ;
  assign n896 = n686 & ~n895 ;
  assign n897 = n780 & ~n896 ;
  assign n898 = ~n780 & n896 ;
  assign n899 = n897 | n898 ;
  assign n900 = ~pi22 & n691 ;
  assign n901 = ~pi8 & n900 ;
  assign n902 = pi8 & ~n900 ;
  assign n903 = n901 | n902 ;
  assign n904 = n216 & n903 ;
  assign n905 = ~n899 & n904 ;
  assign n906 = n897 | n905 ;
  assign n907 = n773 & n906 ;
  assign n908 = n730 & ~n734 ;
  assign n909 = n221 & n908 ;
  assign n910 = ~n688 & n730 ;
  assign n911 = ~n221 & n910 ;
  assign n912 = n688 | n730 ;
  assign n913 = n44 | n912 ;
  assign n914 = n730 | n734 ;
  assign n915 = n44 & ~n914 ;
  assign n916 = n913 & ~n915 ;
  assign n917 = ~n911 & n916 ;
  assign n918 = ~n909 & n917 ;
  assign n919 = n372 | n720 ;
  assign n920 = n534 & n716 ;
  assign n921 = n372 & ~n718 ;
  assign n922 = ~n534 & n722 ;
  assign n923 = n921 | n922 ;
  assign n924 = n920 | n923 ;
  assign n925 = n919 & ~n924 ;
  assign n926 = n918 & n925 ;
  assign n927 = n559 & n705 ;
  assign n928 = n355 & ~n705 ;
  assign n929 = n554 | n696 ;
  assign n930 = ~n358 & n696 ;
  assign n931 = n929 & ~n930 ;
  assign n932 = ~n928 & n931 ;
  assign n933 = ~n927 & n932 ;
  assign n934 = n918 & ~n925 ;
  assign n935 = ~n918 & n925 ;
  assign n936 = n934 | n935 ;
  assign n937 = n933 & n936 ;
  assign n938 = n926 | n937 ;
  assign n939 = n773 | n906 ;
  assign n940 = ~n907 & n939 ;
  assign n941 = n938 & n940 ;
  assign n942 = n907 | n941 ;
  assign n943 = n700 & ~n706 ;
  assign n944 = n707 | n943 ;
  assign n945 = n942 & ~n944 ;
  assign n946 = ~n942 & n944 ;
  assign n947 = n945 | n946 ;
  assign n948 = n748 | n750 ;
  assign n949 = ~n751 & n948 ;
  assign n950 = ~n947 & n949 ;
  assign n951 = n945 | n950 ;
  assign n952 = ~n766 & n951 ;
  assign n953 = n766 & ~n951 ;
  assign n954 = n952 | n953 ;
  assign n955 = n559 & n696 ;
  assign n956 = n355 & ~n696 ;
  assign n957 = n554 | n903 ;
  assign n958 = ~n358 & n903 ;
  assign n959 = n957 & ~n958 ;
  assign n960 = ~n956 & n959 ;
  assign n961 = ~n955 & n960 ;
  assign n962 = n705 | n720 ;
  assign n963 = n372 & n716 ;
  assign n964 = n705 & ~n718 ;
  assign n965 = ~n372 & n722 ;
  assign n966 = n964 | n965 ;
  assign n967 = n963 | n966 ;
  assign n968 = n962 & ~n967 ;
  assign n969 = n961 & n968 ;
  assign n970 = n183 | n496 ;
  assign n971 = n302 | n970 ;
  assign n972 = n291 | n314 ;
  assign n973 = n318 | n972 ;
  assign n974 = n182 | n283 ;
  assign n975 = n261 | n974 ;
  assign n976 = n340 | n975 ;
  assign n977 = n973 | n976 ;
  assign n978 = n971 | n977 ;
  assign n979 = n862 | n978 ;
  assign n980 = n463 | n979 ;
  assign n981 = n430 | n980 ;
  assign n982 = n281 | n981 ;
  assign n983 = n198 | n982 ;
  assign n984 = n227 | n983 ;
  assign n985 = n272 | n325 ;
  assign n986 = n377 | n617 ;
  assign n987 = n813 | n986 ;
  assign n988 = n125 | n244 ;
  assign n989 = n106 | n988 ;
  assign n990 = n987 | n989 ;
  assign n991 = n985 | n990 ;
  assign n992 = n230 | n991 ;
  assign n993 = n154 | n165 ;
  assign n994 = n992 | n993 ;
  assign n995 = n237 | n268 ;
  assign n996 = n293 | n995 ;
  assign n997 = n278 | n332 ;
  assign n998 = n189 | n267 ;
  assign n999 = n997 | n998 ;
  assign n1000 = n996 | n999 ;
  assign n1001 = n188 | n317 ;
  assign n1002 = n315 | n386 ;
  assign n1003 = n1001 | n1002 ;
  assign n1004 = n204 | n260 ;
  assign n1005 = n201 | n500 ;
  assign n1006 = n1004 | n1005 ;
  assign n1007 = n1003 | n1006 ;
  assign n1008 = n1000 | n1007 ;
  assign n1009 = n994 | n1008 ;
  assign n1010 = n224 | n380 ;
  assign n1011 = n114 | n206 ;
  assign n1012 = n1010 | n1011 ;
  assign n1013 = n403 | n1012 ;
  assign n1014 = n825 & ~n1013 ;
  assign n1015 = n164 | n294 ;
  assign n1016 = n650 | n1015 ;
  assign n1017 = n265 | n1016 ;
  assign n1018 = n1014 & ~n1017 ;
  assign n1019 = ~n1009 & n1018 ;
  assign n1020 = ~n149 & n1019 ;
  assign n1021 = ~n984 & n1020 ;
  assign n1022 = ~n177 & n1021 ;
  assign n1023 = ~n271 & n1022 ;
  assign n1024 = ~n313 & n1023 ;
  assign n1025 = ~n374 & n1024 ;
  assign n1026 = n375 | n848 ;
  assign n1027 = n240 | n315 ;
  assign n1028 = n1026 | n1027 ;
  assign n1029 = n301 | n338 ;
  assign n1030 = n143 | n396 ;
  assign n1031 = n121 | n1010 ;
  assign n1032 = n604 | n1031 ;
  assign n1033 = n289 | n1032 ;
  assign n1034 = n1030 | n1033 ;
  assign n1035 = n237 | n317 ;
  assign n1036 = n190 | n1035 ;
  assign n1037 = n269 | n278 ;
  assign n1038 = n1036 | n1037 ;
  assign n1039 = n439 | n830 ;
  assign n1040 = n1038 | n1039 ;
  assign n1041 = n203 | n1040 ;
  assign n1042 = n1034 | n1041 ;
  assign n1043 = n865 | n1042 ;
  assign n1044 = n1029 | n1043 ;
  assign n1045 = n137 | n318 ;
  assign n1046 = n316 | n398 ;
  assign n1047 = n126 | n282 ;
  assign n1048 = n204 | n1047 ;
  assign n1049 = n266 | n1048 ;
  assign n1050 = n334 | n1049 ;
  assign n1051 = n275 | n1050 ;
  assign n1052 = n659 | n1051 ;
  assign n1053 = n1046 | n1052 ;
  assign n1054 = n291 | n431 ;
  assign n1055 = n164 | n1054 ;
  assign n1056 = n798 | n1055 ;
  assign n1057 = n125 | n374 ;
  assign n1058 = n174 | n1057 ;
  assign n1059 = n584 | n1058 ;
  assign n1060 = n1056 | n1059 ;
  assign n1061 = ~n498 & n824 ;
  assign n1062 = ~n884 & n1061 ;
  assign n1063 = ~n246 & n1062 ;
  assign n1064 = ~n1060 & n1063 ;
  assign n1065 = ~n187 & n1064 ;
  assign n1066 = ~n114 & n1065 ;
  assign n1067 = n400 | n618 ;
  assign n1068 = n650 | n1067 ;
  assign n1069 = n389 | n1068 ;
  assign n1070 = n1066 & ~n1069 ;
  assign n1071 = ~n145 & n1070 ;
  assign n1072 = ~n207 & n1071 ;
  assign n1073 = ~n1053 & n1072 ;
  assign n1074 = ~n1045 & n1073 ;
  assign n1075 = ~n1044 & n1074 ;
  assign n1076 = ~n1028 & n1075 ;
  assign n1077 = n1025 | n1076 ;
  assign n1078 = ~n845 & n1077 ;
  assign n1079 = n1025 & ~n1078 ;
  assign n1080 = ~pi6 & n774 ;
  assign n1081 = pi6 & ~n774 ;
  assign n1082 = n1080 | n1081 ;
  assign n1083 = n216 & n1082 ;
  assign n1084 = ~n1025 & n1078 ;
  assign n1085 = n1079 | n1084 ;
  assign n1086 = n1083 & ~n1085 ;
  assign n1087 = n1079 | n1086 ;
  assign n1088 = n961 | n968 ;
  assign n1089 = ~n969 & n1088 ;
  assign n1090 = n1087 & n1089 ;
  assign n1091 = n969 | n1090 ;
  assign n1092 = n221 | n896 ;
  assign n1093 = n845 & ~n894 ;
  assign n1094 = n686 | n1093 ;
  assign n1095 = n845 & n894 ;
  assign n1096 = n845 | n894 ;
  assign n1097 = ~n1095 & n1096 ;
  assign n1098 = n1094 & n1097 ;
  assign n1099 = n221 & n1098 ;
  assign n1100 = n896 | n1097 ;
  assign n1101 = ~n1099 & n1100 ;
  assign n1102 = n1092 & n1101 ;
  assign n1103 = ~n780 & n1102 ;
  assign n1104 = n780 & ~n1102 ;
  assign n1105 = n1103 | n1104 ;
  assign n1106 = ~n44 & n910 ;
  assign n1107 = n534 | n912 ;
  assign n1108 = n44 & n908 ;
  assign n1109 = n534 & ~n914 ;
  assign n1110 = n1108 | n1109 ;
  assign n1111 = n1107 & ~n1110 ;
  assign n1112 = ~n1106 & n1111 ;
  assign n1113 = ~n1105 & n1112 ;
  assign n1114 = n1103 | n1113 ;
  assign n1115 = n1091 & n1114 ;
  assign n1116 = n1091 | n1114 ;
  assign n1117 = ~n1115 & n1116 ;
  assign n1118 = n899 & ~n904 ;
  assign n1119 = n905 | n1118 ;
  assign n1120 = n1117 & ~n1119 ;
  assign n1121 = n1115 | n1120 ;
  assign n1122 = n739 & ~n746 ;
  assign n1123 = n747 | n1122 ;
  assign n1124 = n1121 & ~n1123 ;
  assign n1125 = ~n1121 & n1123 ;
  assign n1126 = n1124 | n1125 ;
  assign n1127 = n938 | n940 ;
  assign n1128 = ~n941 & n1127 ;
  assign n1129 = ~n1126 & n1128 ;
  assign n1130 = n1124 | n1129 ;
  assign n1131 = n947 & ~n949 ;
  assign n1132 = n950 | n1131 ;
  assign n1133 = n1130 & ~n1132 ;
  assign n1134 = n933 | n936 ;
  assign n1135 = ~n937 & n1134 ;
  assign n1136 = n1105 & ~n1112 ;
  assign n1137 = n1113 | n1136 ;
  assign n1138 = n559 & n903 ;
  assign n1139 = n355 & ~n903 ;
  assign n1140 = n554 | n779 ;
  assign n1141 = ~n358 & n779 ;
  assign n1142 = n1140 & ~n1141 ;
  assign n1143 = ~n1139 & n1142 ;
  assign n1144 = ~n1138 & n1143 ;
  assign n1145 = n696 | n720 ;
  assign n1146 = n705 & n716 ;
  assign n1147 = n1145 & ~n1146 ;
  assign n1148 = n696 & ~n718 ;
  assign n1149 = ~n705 & n722 ;
  assign n1150 = n1148 | n1149 ;
  assign n1151 = n1147 & ~n1150 ;
  assign n1152 = n1144 & n1151 ;
  assign n1153 = n1144 | n1151 ;
  assign n1154 = ~n1152 & n1153 ;
  assign n1155 = n221 | n1100 ;
  assign n1156 = ~n896 & n1097 ;
  assign n1157 = ~n44 & n1156 ;
  assign n1158 = n1094 & ~n1097 ;
  assign n1159 = n221 & n1158 ;
  assign n1160 = n44 & n1098 ;
  assign n1161 = n1159 | n1160 ;
  assign n1162 = n1157 | n1161 ;
  assign n1163 = n1155 & ~n1162 ;
  assign n1164 = n1154 & n1163 ;
  assign n1165 = n1152 | n1164 ;
  assign n1166 = ~n1137 & n1165 ;
  assign n1167 = n1087 | n1089 ;
  assign n1168 = ~n1090 & n1167 ;
  assign n1169 = n1137 & ~n1152 ;
  assign n1170 = ~n1164 & n1169 ;
  assign n1171 = n1168 & ~n1170 ;
  assign n1172 = ~n1166 & n1171 ;
  assign n1173 = n1166 | n1172 ;
  assign n1174 = n1135 & n1173 ;
  assign n1175 = n1135 | n1173 ;
  assign n1176 = ~n1174 & n1175 ;
  assign n1177 = ~n1117 & n1119 ;
  assign n1178 = n1120 | n1177 ;
  assign n1179 = n1176 & ~n1178 ;
  assign n1180 = n1174 | n1179 ;
  assign n1181 = n1126 & ~n1128 ;
  assign n1182 = n1129 | n1181 ;
  assign n1183 = n1180 & ~n1182 ;
  assign n1184 = ~n1083 & n1085 ;
  assign n1185 = n1086 | n1184 ;
  assign n1186 = ~n534 & n910 ;
  assign n1187 = n372 | n912 ;
  assign n1188 = n534 & n908 ;
  assign n1189 = n372 & ~n914 ;
  assign n1190 = n1188 | n1189 ;
  assign n1191 = n1187 & ~n1190 ;
  assign n1192 = ~n1186 & n1191 ;
  assign n1193 = ~n1185 & n1192 ;
  assign n1194 = n1185 & ~n1192 ;
  assign n1195 = n1193 | n1194 ;
  assign n1196 = ~pi22 & n689 ;
  assign n1197 = pi5 & ~n1196 ;
  assign n1198 = ~pi5 & n1196 ;
  assign n1199 = n1197 | n1198 ;
  assign n1200 = n216 & n1199 ;
  assign n1201 = n1025 & ~n1200 ;
  assign n1202 = n1025 & ~n1076 ;
  assign n1203 = ~n1025 & n1076 ;
  assign n1204 = n1202 | n1203 ;
  assign n1205 = n221 & ~n1204 ;
  assign n1206 = n1078 | n1205 ;
  assign n1207 = n1025 & n1076 ;
  assign n1208 = n845 & ~n1207 ;
  assign n1209 = n1205 & ~n1208 ;
  assign n1210 = n1206 & ~n1209 ;
  assign n1211 = ~n1201 & n1210 ;
  assign n1212 = ~n1025 & n1200 ;
  assign n1213 = n1211 | n1212 ;
  assign n1214 = ~n1195 & n1213 ;
  assign n1215 = n1193 | n1214 ;
  assign n1216 = ~n372 & n910 ;
  assign n1217 = n705 | n912 ;
  assign n1218 = n372 & n908 ;
  assign n1219 = n705 & ~n914 ;
  assign n1220 = n1218 | n1219 ;
  assign n1221 = n1217 & ~n1220 ;
  assign n1222 = ~n1216 & n1221 ;
  assign n1223 = n44 | n1100 ;
  assign n1224 = ~n534 & n1156 ;
  assign n1225 = n44 & n1158 ;
  assign n1226 = n534 & n1098 ;
  assign n1227 = n1225 | n1226 ;
  assign n1228 = n1224 | n1227 ;
  assign n1229 = n1223 & ~n1228 ;
  assign n1230 = n1222 & n1229 ;
  assign n1231 = n1222 | n1229 ;
  assign n1232 = ~n1230 & n1231 ;
  assign n1233 = n696 & n716 ;
  assign n1234 = ~n718 & n903 ;
  assign n1235 = n720 | n903 ;
  assign n1236 = ~n696 & n722 ;
  assign n1237 = n1235 & ~n1236 ;
  assign n1238 = ~n1234 & n1237 ;
  assign n1239 = ~n1233 & n1238 ;
  assign n1240 = n1232 & n1239 ;
  assign n1241 = n1230 | n1240 ;
  assign n1242 = n1154 | n1163 ;
  assign n1243 = ~n1164 & n1242 ;
  assign n1244 = n1241 & n1243 ;
  assign n1245 = ~pi22 & n36 ;
  assign n1246 = ~pi4 & n1245 ;
  assign n1247 = pi4 & ~n1245 ;
  assign n1248 = n1246 | n1247 ;
  assign n1249 = n216 & n1248 ;
  assign n1250 = ~n1025 & n1249 ;
  assign n1251 = n1025 & ~n1249 ;
  assign n1252 = n1204 & ~n1208 ;
  assign n1253 = n221 & n1252 ;
  assign n1254 = n1204 | n1208 ;
  assign n1255 = n44 & ~n1254 ;
  assign n1256 = n1078 | n1204 ;
  assign n1257 = n44 | n1256 ;
  assign n1258 = ~n1078 & n1204 ;
  assign n1259 = ~n221 & n1258 ;
  assign n1260 = n1257 & ~n1259 ;
  assign n1261 = ~n1255 & n1260 ;
  assign n1262 = ~n1253 & n1261 ;
  assign n1263 = ~n1251 & n1262 ;
  assign n1264 = ~n1250 & n1263 ;
  assign n1265 = n1250 | n1264 ;
  assign n1266 = n559 & n779 ;
  assign n1267 = n355 & ~n779 ;
  assign n1268 = n554 | n1082 ;
  assign n1269 = ~n358 & n1082 ;
  assign n1270 = n1268 & ~n1269 ;
  assign n1271 = ~n1267 & n1270 ;
  assign n1272 = ~n1266 & n1271 ;
  assign n1273 = n1265 & n1272 ;
  assign n1274 = n1265 | n1272 ;
  assign n1275 = ~n1273 & n1274 ;
  assign n1276 = n705 & n908 ;
  assign n1277 = ~n705 & n910 ;
  assign n1278 = n696 | n912 ;
  assign n1279 = n696 & ~n914 ;
  assign n1280 = n1278 & ~n1279 ;
  assign n1281 = ~n1277 & n1280 ;
  assign n1282 = ~n1276 & n1281 ;
  assign n1283 = n534 & n1158 ;
  assign n1284 = n534 | n1100 ;
  assign n1285 = ~n372 & n1156 ;
  assign n1286 = n372 & n1098 ;
  assign n1287 = n1285 | n1286 ;
  assign n1288 = n1284 & ~n1287 ;
  assign n1289 = ~n1283 & n1288 ;
  assign n1290 = n1282 & n1289 ;
  assign n1291 = n1282 | n1289 ;
  assign n1292 = ~n1290 & n1291 ;
  assign n1293 = n716 & n903 ;
  assign n1294 = ~n718 & n779 ;
  assign n1295 = n720 | n779 ;
  assign n1296 = n722 & ~n903 ;
  assign n1297 = n1295 & ~n1296 ;
  assign n1298 = ~n1294 & n1297 ;
  assign n1299 = ~n1293 & n1298 ;
  assign n1300 = n1292 & n1299 ;
  assign n1301 = n1290 | n1300 ;
  assign n1302 = n1275 & n1301 ;
  assign n1303 = n1273 | n1302 ;
  assign n1304 = n1241 | n1243 ;
  assign n1305 = ~n1244 & n1304 ;
  assign n1306 = n1303 & n1305 ;
  assign n1307 = n1244 | n1306 ;
  assign n1308 = n1215 & n1307 ;
  assign n1309 = n1215 | n1307 ;
  assign n1310 = ~n1308 & n1309 ;
  assign n1311 = n1166 | n1170 ;
  assign n1312 = ~n1168 & n1311 ;
  assign n1313 = n1172 | n1312 ;
  assign n1314 = n1310 & ~n1313 ;
  assign n1315 = n1308 | n1314 ;
  assign n1316 = ~n1176 & n1178 ;
  assign n1317 = n1179 | n1316 ;
  assign n1318 = n1315 & ~n1317 ;
  assign n1319 = n1201 | n1212 ;
  assign n1320 = n1210 | n1319 ;
  assign n1321 = n1210 & n1319 ;
  assign n1322 = n1320 & ~n1321 ;
  assign n1323 = n1232 | n1239 ;
  assign n1324 = ~n1240 & n1323 ;
  assign n1325 = ~n1322 & n1324 ;
  assign n1326 = n1322 & ~n1324 ;
  assign n1327 = n1325 | n1326 ;
  assign n1328 = n559 & n1082 ;
  assign n1329 = n355 & ~n1082 ;
  assign n1330 = n554 | n1199 ;
  assign n1331 = ~n358 & n1199 ;
  assign n1332 = n1330 & ~n1331 ;
  assign n1333 = ~n1329 & n1332 ;
  assign n1334 = ~n1328 & n1333 ;
  assign n1335 = ~pi22 & n35 ;
  assign n1336 = pi3 & ~n1335 ;
  assign n1337 = pi3 | pi22 ;
  assign n1338 = n35 & ~n1337 ;
  assign n1339 = n1336 | n1338 ;
  assign n1340 = n216 & n1339 ;
  assign n1341 = n178 | n317 ;
  assign n1342 = n204 | n374 ;
  assign n1343 = n1341 | n1342 ;
  assign n1344 = n380 | n496 ;
  assign n1345 = n326 | n618 ;
  assign n1346 = n121 | n316 ;
  assign n1347 = n189 | n1346 ;
  assign n1348 = n175 | n1347 ;
  assign n1349 = n462 | n1348 ;
  assign n1350 = n378 | n883 ;
  assign n1351 = n1349 | n1350 ;
  assign n1352 = n193 | n1351 ;
  assign n1353 = n164 | n1352 ;
  assign n1354 = n260 | n310 ;
  assign n1355 = n1353 | n1354 ;
  assign n1356 = n155 | n1355 ;
  assign n1357 = n294 | n340 ;
  assign n1358 = ~n302 & n824 ;
  assign n1359 = n240 | n333 ;
  assign n1360 = n243 | n1359 ;
  assign n1361 = n1358 & ~n1360 ;
  assign n1362 = ~n1357 & n1361 ;
  assign n1363 = ~n248 & n1362 ;
  assign n1364 = ~n400 & n1363 ;
  assign n1365 = ~n390 & n1364 ;
  assign n1366 = ~n1356 & n1365 ;
  assign n1367 = ~n153 & n1366 ;
  assign n1368 = n201 | n619 ;
  assign n1369 = n192 | n1368 ;
  assign n1370 = n597 | n1369 ;
  assign n1371 = n287 | n1370 ;
  assign n1372 = n161 | n1371 ;
  assign n1373 = n1367 & ~n1372 ;
  assign n1374 = ~n1345 & n1373 ;
  assign n1375 = ~n1344 & n1374 ;
  assign n1376 = ~n1343 & n1375 ;
  assign n1377 = ~n379 & n1376 ;
  assign n1378 = n221 & n1377 ;
  assign n1379 = n1025 | n1378 ;
  assign n1380 = n1340 & ~n1379 ;
  assign n1381 = ~n1340 & n1379 ;
  assign n1382 = n1380 | n1381 ;
  assign n1383 = n44 & n1252 ;
  assign n1384 = n534 & ~n1254 ;
  assign n1385 = n534 | n1256 ;
  assign n1386 = ~n44 & n1258 ;
  assign n1387 = n1385 & ~n1386 ;
  assign n1388 = ~n1384 & n1387 ;
  assign n1389 = ~n1383 & n1388 ;
  assign n1390 = ~n1382 & n1389 ;
  assign n1391 = n1380 | n1390 ;
  assign n1392 = n1334 & n1391 ;
  assign n1393 = n1334 | n1391 ;
  assign n1394 = ~n1392 & n1393 ;
  assign n1395 = n696 & n908 ;
  assign n1396 = ~n696 & n910 ;
  assign n1397 = n903 | n912 ;
  assign n1398 = n903 & ~n914 ;
  assign n1399 = n1397 & ~n1398 ;
  assign n1400 = ~n1396 & n1399 ;
  assign n1401 = ~n1395 & n1400 ;
  assign n1402 = n372 & n1158 ;
  assign n1403 = n372 | n1100 ;
  assign n1404 = ~n705 & n1156 ;
  assign n1405 = n705 & n1098 ;
  assign n1406 = n1404 | n1405 ;
  assign n1407 = n1403 & ~n1406 ;
  assign n1408 = ~n1402 & n1407 ;
  assign n1409 = n1401 & n1408 ;
  assign n1410 = n1401 | n1408 ;
  assign n1411 = ~n1409 & n1410 ;
  assign n1412 = n722 & ~n779 ;
  assign n1413 = n720 | n1082 ;
  assign n1414 = n716 & n779 ;
  assign n1415 = ~n718 & n1082 ;
  assign n1416 = n1414 | n1415 ;
  assign n1417 = n1413 & ~n1416 ;
  assign n1418 = ~n1412 & n1417 ;
  assign n1419 = n1411 & n1418 ;
  assign n1420 = n1409 | n1419 ;
  assign n1421 = n1394 & n1420 ;
  assign n1422 = n1392 | n1421 ;
  assign n1423 = ~n1327 & n1422 ;
  assign n1424 = n1325 | n1423 ;
  assign n1425 = n1195 & ~n1213 ;
  assign n1426 = n1214 | n1425 ;
  assign n1427 = n1424 & ~n1426 ;
  assign n1428 = n1303 | n1305 ;
  assign n1429 = ~n1306 & n1428 ;
  assign n1430 = ~n1325 & n1426 ;
  assign n1431 = ~n1423 & n1430 ;
  assign n1432 = n1429 & ~n1431 ;
  assign n1433 = ~n1427 & n1432 ;
  assign n1434 = n1427 | n1433 ;
  assign n1435 = ~n1310 & n1313 ;
  assign n1436 = n1314 | n1435 ;
  assign n1437 = n1434 & ~n1436 ;
  assign n1438 = n1427 | n1431 ;
  assign n1439 = ~n1429 & n1438 ;
  assign n1440 = n1275 | n1301 ;
  assign n1441 = ~n1302 & n1440 ;
  assign n1442 = n559 & n1339 ;
  assign n1443 = n350 & n554 ;
  assign n1444 = ~n1442 & n1443 ;
  assign n1445 = n221 & ~n1377 ;
  assign n1446 = n1025 & ~n1445 ;
  assign n1447 = ~n1025 & n1445 ;
  assign n1448 = n44 & n1377 ;
  assign n1449 = n1447 | n1448 ;
  assign n1450 = n1446 | n1449 ;
  assign n1451 = n1444 & ~n1450 ;
  assign n1452 = n559 & n1199 ;
  assign n1453 = n355 & ~n1199 ;
  assign n1454 = n554 | n1248 ;
  assign n1455 = ~n358 & n1248 ;
  assign n1456 = n1454 & ~n1455 ;
  assign n1457 = ~n1453 & n1456 ;
  assign n1458 = ~n1452 & n1457 ;
  assign n1459 = n1451 & n1458 ;
  assign n1460 = n1451 | n1458 ;
  assign n1461 = ~n1459 & n1460 ;
  assign n1462 = n722 & ~n1082 ;
  assign n1463 = n720 | n1199 ;
  assign n1464 = n716 & n1082 ;
  assign n1465 = ~n718 & n1199 ;
  assign n1466 = n1464 | n1465 ;
  assign n1467 = n1463 & ~n1466 ;
  assign n1468 = ~n1462 & n1467 ;
  assign n1469 = n903 & n908 ;
  assign n1470 = ~n903 & n910 ;
  assign n1471 = n779 | n912 ;
  assign n1472 = n779 & ~n914 ;
  assign n1473 = n1471 & ~n1472 ;
  assign n1474 = ~n1470 & n1473 ;
  assign n1475 = ~n1469 & n1474 ;
  assign n1476 = n1468 & n1475 ;
  assign n1477 = n1468 | n1475 ;
  assign n1478 = ~n1476 & n1477 ;
  assign n1479 = n705 & n1158 ;
  assign n1480 = n705 | n1100 ;
  assign n1481 = ~n696 & n1156 ;
  assign n1482 = n696 & n1098 ;
  assign n1483 = n1481 | n1482 ;
  assign n1484 = n1480 & ~n1483 ;
  assign n1485 = ~n1479 & n1484 ;
  assign n1486 = n1478 & n1485 ;
  assign n1487 = n1476 | n1486 ;
  assign n1488 = n1461 & n1487 ;
  assign n1489 = n1459 | n1488 ;
  assign n1490 = n1251 | n1265 ;
  assign n1491 = n1262 & ~n1264 ;
  assign n1492 = n1490 & ~n1491 ;
  assign n1493 = n1489 | n1492 ;
  assign n1494 = n1489 & n1492 ;
  assign n1495 = n1493 & ~n1494 ;
  assign n1496 = n1292 | n1299 ;
  assign n1497 = ~n1300 & n1496 ;
  assign n1498 = ~n1495 & n1497 ;
  assign n1499 = n1489 & ~n1492 ;
  assign n1500 = n1498 | n1499 ;
  assign n1501 = n1441 & n1500 ;
  assign n1502 = n1441 | n1500 ;
  assign n1503 = ~n1501 & n1502 ;
  assign n1504 = n1327 & ~n1422 ;
  assign n1505 = n1423 | n1504 ;
  assign n1506 = n1503 & ~n1505 ;
  assign n1507 = n1501 | n1506 ;
  assign n1508 = ~n1433 & n1507 ;
  assign n1509 = ~n1439 & n1508 ;
  assign n1510 = ~n1503 & n1505 ;
  assign n1511 = n1506 | n1510 ;
  assign n1512 = n559 & n1248 ;
  assign n1513 = n355 & ~n1248 ;
  assign n1514 = n1512 | n1513 ;
  assign n1515 = n554 | n1339 ;
  assign n1516 = ~n358 & n1339 ;
  assign n1517 = n1515 & ~n1516 ;
  assign n1518 = ~n1514 & n1517 ;
  assign n1519 = n534 & n1252 ;
  assign n1520 = n372 & ~n1254 ;
  assign n1521 = n372 | n1256 ;
  assign n1522 = ~n534 & n1258 ;
  assign n1523 = n1521 & ~n1522 ;
  assign n1524 = ~n1520 & n1523 ;
  assign n1525 = ~n1519 & n1524 ;
  assign n1526 = n1518 & n1525 ;
  assign n1527 = n1518 | n1525 ;
  assign n1528 = ~n1444 & n1450 ;
  assign n1529 = n1451 | n1528 ;
  assign n1530 = n1527 & ~n1529 ;
  assign n1531 = n1526 | n1530 ;
  assign n1532 = n1382 & ~n1389 ;
  assign n1533 = n1390 | n1532 ;
  assign n1534 = n1531 & ~n1533 ;
  assign n1535 = ~n1531 & n1533 ;
  assign n1536 = n1534 | n1535 ;
  assign n1537 = n1411 | n1418 ;
  assign n1538 = ~n1419 & n1537 ;
  assign n1539 = ~n1536 & n1538 ;
  assign n1540 = n1534 | n1539 ;
  assign n1541 = n1394 | n1420 ;
  assign n1542 = ~n1421 & n1541 ;
  assign n1543 = n1540 & n1542 ;
  assign n1544 = n1540 | n1542 ;
  assign n1545 = ~n1543 & n1544 ;
  assign n1546 = n1495 & ~n1497 ;
  assign n1547 = n1498 | n1546 ;
  assign n1548 = n1545 & ~n1547 ;
  assign n1549 = n1543 | n1548 ;
  assign n1550 = ~n1511 & n1549 ;
  assign n1551 = n1511 & ~n1549 ;
  assign n1552 = n1550 | n1551 ;
  assign n1553 = n372 & n1252 ;
  assign n1554 = n705 & ~n1254 ;
  assign n1555 = n705 | n1256 ;
  assign n1556 = ~n372 & n1258 ;
  assign n1557 = n1555 & ~n1556 ;
  assign n1558 = ~n1554 & n1557 ;
  assign n1559 = ~n1553 & n1558 ;
  assign n1560 = n44 & ~n1377 ;
  assign n1561 = n1025 & ~n1560 ;
  assign n1562 = n534 & n1377 ;
  assign n1563 = ~n1025 & n1560 ;
  assign n1564 = n1562 | n1563 ;
  assign n1565 = n1561 | n1564 ;
  assign n1566 = n1559 & ~n1565 ;
  assign n1567 = ~n1559 & n1565 ;
  assign n1568 = n1566 | n1567 ;
  assign n1569 = n722 & ~n1199 ;
  assign n1570 = n720 | n1248 ;
  assign n1571 = n716 & n1199 ;
  assign n1572 = ~n718 & n1248 ;
  assign n1573 = n1571 | n1572 ;
  assign n1574 = n1570 & ~n1573 ;
  assign n1575 = ~n1569 & n1574 ;
  assign n1576 = ~n1568 & n1575 ;
  assign n1577 = n1566 | n1576 ;
  assign n1578 = n696 & n1158 ;
  assign n1579 = n696 | n1100 ;
  assign n1580 = ~n903 & n1156 ;
  assign n1581 = n903 & n1098 ;
  assign n1582 = n1580 | n1581 ;
  assign n1583 = n1579 & ~n1582 ;
  assign n1584 = ~n1578 & n1583 ;
  assign n1585 = n779 & n908 ;
  assign n1586 = ~n779 & n910 ;
  assign n1587 = n912 | n1082 ;
  assign n1588 = ~n914 & n1082 ;
  assign n1589 = n1587 & ~n1588 ;
  assign n1590 = ~n1586 & n1589 ;
  assign n1591 = ~n1585 & n1590 ;
  assign n1592 = n1584 & n1591 ;
  assign n1593 = n1584 | n1591 ;
  assign n1594 = ~n1592 & n1593 ;
  assign n1595 = n372 & n1377 ;
  assign n1596 = n534 & ~n1377 ;
  assign n1597 = ~n1025 & n1596 ;
  assign n1598 = n1025 & ~n1596 ;
  assign n1599 = n1597 | n1598 ;
  assign n1600 = n1595 | n1599 ;
  assign n1601 = n547 & n1339 ;
  assign n1602 = n525 & ~n1601 ;
  assign n1603 = ~n1600 & n1602 ;
  assign n1604 = n1594 & n1603 ;
  assign n1605 = n1592 | n1604 ;
  assign n1606 = n1577 & n1605 ;
  assign n1607 = n1577 | n1605 ;
  assign n1608 = ~n1606 & n1607 ;
  assign n1609 = n1478 | n1485 ;
  assign n1610 = ~n1486 & n1609 ;
  assign n1611 = n1608 & n1610 ;
  assign n1612 = n1606 | n1611 ;
  assign n1613 = n1461 | n1487 ;
  assign n1614 = ~n1488 & n1613 ;
  assign n1615 = n1612 & n1614 ;
  assign n1616 = n1612 | n1614 ;
  assign n1617 = ~n1615 & n1616 ;
  assign n1618 = n1536 & ~n1538 ;
  assign n1619 = n1539 | n1618 ;
  assign n1620 = n1617 & ~n1619 ;
  assign n1621 = n1615 | n1620 ;
  assign n1622 = ~n1545 & n1547 ;
  assign n1623 = n1548 | n1622 ;
  assign n1624 = n1621 & ~n1623 ;
  assign n1625 = ~n1617 & n1619 ;
  assign n1626 = n1620 | n1625 ;
  assign n1627 = n554 & n1339 ;
  assign n1628 = ~n559 & n1627 ;
  assign n1629 = n350 | n1628 ;
  assign n1630 = ~n705 & n1258 ;
  assign n1631 = n696 | n1256 ;
  assign n1632 = n705 & n1252 ;
  assign n1633 = n696 & ~n1254 ;
  assign n1634 = n1632 | n1633 ;
  assign n1635 = n1631 & ~n1634 ;
  assign n1636 = ~n1630 & n1635 ;
  assign n1637 = n908 & n1082 ;
  assign n1638 = n910 & ~n1082 ;
  assign n1639 = n912 | n1199 ;
  assign n1640 = ~n914 & n1199 ;
  assign n1641 = n1639 & ~n1640 ;
  assign n1642 = ~n1638 & n1641 ;
  assign n1643 = ~n1637 & n1642 ;
  assign n1644 = n1636 & n1643 ;
  assign n1645 = n1636 | n1643 ;
  assign n1646 = ~n1644 & n1645 ;
  assign n1647 = n903 & n1158 ;
  assign n1648 = n903 | n1100 ;
  assign n1649 = ~n779 & n1156 ;
  assign n1650 = n779 & n1098 ;
  assign n1651 = n1649 | n1650 ;
  assign n1652 = n1648 & ~n1651 ;
  assign n1653 = ~n1647 & n1652 ;
  assign n1654 = n1646 & n1653 ;
  assign n1655 = n1644 | n1654 ;
  assign n1656 = ~n1444 & n1655 ;
  assign n1657 = n1629 & n1656 ;
  assign n1658 = ~n1444 & n1629 ;
  assign n1659 = n1655 | n1658 ;
  assign n1660 = n1594 | n1603 ;
  assign n1661 = ~n1604 & n1660 ;
  assign n1662 = ~n1657 & n1661 ;
  assign n1663 = n1659 & n1662 ;
  assign n1664 = n1657 | n1663 ;
  assign n1665 = ~n1526 & n1527 ;
  assign n1666 = n1529 | n1665 ;
  assign n1667 = n1529 & n1665 ;
  assign n1668 = n1666 & ~n1667 ;
  assign n1669 = n1664 & ~n1668 ;
  assign n1670 = n1608 | n1610 ;
  assign n1671 = ~n1611 & n1670 ;
  assign n1672 = ~n1664 & n1668 ;
  assign n1673 = n1669 | n1672 ;
  assign n1674 = n1671 & ~n1673 ;
  assign n1675 = n1669 | n1674 ;
  assign n1676 = ~n1626 & n1675 ;
  assign n1677 = n1626 & ~n1675 ;
  assign n1678 = n1676 | n1677 ;
  assign n1679 = n1568 & ~n1575 ;
  assign n1680 = n1576 | n1679 ;
  assign n1681 = n1600 & ~n1602 ;
  assign n1682 = n1603 | n1681 ;
  assign n1683 = n716 & n1248 ;
  assign n1684 = n722 & ~n1248 ;
  assign n1685 = n720 | n1339 ;
  assign n1686 = ~n718 & n1339 ;
  assign n1687 = n1685 & ~n1686 ;
  assign n1688 = ~n1684 & n1687 ;
  assign n1689 = ~n1683 & n1688 ;
  assign n1690 = ~n1682 & n1689 ;
  assign n1691 = ~n696 & n1258 ;
  assign n1692 = n903 | n1256 ;
  assign n1693 = n696 & n1252 ;
  assign n1694 = n903 & ~n1254 ;
  assign n1695 = n1693 | n1694 ;
  assign n1696 = n1692 & ~n1695 ;
  assign n1697 = ~n1691 & n1696 ;
  assign n1698 = n372 & ~n1377 ;
  assign n1699 = ~n1025 & n1698 ;
  assign n1700 = n1025 & ~n1698 ;
  assign n1701 = n705 & n1377 ;
  assign n1702 = n1700 | n1701 ;
  assign n1703 = n1699 | n1702 ;
  assign n1704 = n1697 & ~n1703 ;
  assign n1705 = ~n1697 & n1703 ;
  assign n1706 = n1704 | n1705 ;
  assign n1707 = n779 & n1158 ;
  assign n1708 = n779 | n1100 ;
  assign n1709 = ~n1082 & n1156 ;
  assign n1710 = n1082 & n1098 ;
  assign n1711 = n1709 | n1710 ;
  assign n1712 = n1708 & ~n1711 ;
  assign n1713 = ~n1707 & n1712 ;
  assign n1714 = ~n1706 & n1713 ;
  assign n1715 = n1704 | n1714 ;
  assign n1716 = n1682 & ~n1689 ;
  assign n1717 = n1690 | n1716 ;
  assign n1718 = n1715 & ~n1717 ;
  assign n1719 = n1690 | n1718 ;
  assign n1720 = ~n1680 & n1719 ;
  assign n1721 = ~n1657 & n1659 ;
  assign n1722 = n1661 | n1721 ;
  assign n1723 = n1680 & ~n1719 ;
  assign n1724 = n1720 | n1723 ;
  assign n1725 = n1663 | n1724 ;
  assign n1726 = n1722 & ~n1725 ;
  assign n1727 = n1720 | n1726 ;
  assign n1728 = ~n1671 & n1673 ;
  assign n1729 = n1674 | n1728 ;
  assign n1730 = n1727 & ~n1729 ;
  assign n1731 = ~n1727 & n1729 ;
  assign n1732 = ~n903 & n1258 ;
  assign n1733 = n779 | n1256 ;
  assign n1734 = n903 & n1252 ;
  assign n1735 = n779 & ~n1254 ;
  assign n1736 = n1734 | n1735 ;
  assign n1737 = n1733 & ~n1736 ;
  assign n1738 = ~n1732 & n1737 ;
  assign n1739 = n1082 & n1158 ;
  assign n1740 = n1082 | n1100 ;
  assign n1741 = n1156 & ~n1199 ;
  assign n1742 = n1098 & n1199 ;
  assign n1743 = n1741 | n1742 ;
  assign n1744 = n1740 & ~n1743 ;
  assign n1745 = ~n1739 & n1744 ;
  assign n1746 = n1738 & n1745 ;
  assign n1747 = n1738 | n1745 ;
  assign n1748 = ~n1746 & n1747 ;
  assign n1749 = n908 & n1248 ;
  assign n1750 = n910 & ~n1248 ;
  assign n1751 = n912 | n1339 ;
  assign n1752 = ~n914 & n1339 ;
  assign n1753 = n1751 & ~n1752 ;
  assign n1754 = ~n1750 & n1753 ;
  assign n1755 = ~n1749 & n1754 ;
  assign n1756 = n1748 & n1755 ;
  assign n1757 = n1746 | n1756 ;
  assign n1758 = n1706 & ~n1713 ;
  assign n1759 = n1714 | n1758 ;
  assign n1760 = n1757 & ~n1759 ;
  assign n1761 = n544 & n1339 ;
  assign n1762 = n688 | n1339 ;
  assign n1763 = n908 & n1339 ;
  assign n1764 = n912 & ~n1763 ;
  assign n1765 = n1762 & n1764 ;
  assign n1766 = n688 & n1765 ;
  assign n1767 = n705 & ~n1377 ;
  assign n1768 = ~n1025 & n1767 ;
  assign n1769 = n696 | n1025 ;
  assign n1770 = n1377 & n1769 ;
  assign n1771 = ~n705 & n1025 ;
  assign n1772 = n1770 | n1771 ;
  assign n1773 = n1768 | n1772 ;
  assign n1774 = n1766 & ~n1773 ;
  assign n1775 = n908 & n1199 ;
  assign n1776 = n910 & ~n1199 ;
  assign n1777 = n912 | n1248 ;
  assign n1778 = ~n914 & n1248 ;
  assign n1779 = n1777 & ~n1778 ;
  assign n1780 = ~n1776 & n1779 ;
  assign n1781 = ~n1775 & n1780 ;
  assign n1782 = n1774 & n1781 ;
  assign n1783 = n1774 | n1781 ;
  assign n1784 = ~n1782 & n1783 ;
  assign n1785 = n1761 & n1784 ;
  assign n1786 = n1761 | n1784 ;
  assign n1787 = ~n1785 & n1786 ;
  assign n1788 = ~n1757 & n1759 ;
  assign n1789 = n1760 | n1788 ;
  assign n1790 = n1787 & ~n1789 ;
  assign n1791 = n1760 | n1790 ;
  assign n1792 = n1782 | n1785 ;
  assign n1793 = n1646 | n1653 ;
  assign n1794 = ~n1654 & n1793 ;
  assign n1795 = n1792 & n1794 ;
  assign n1796 = n1792 | n1794 ;
  assign n1797 = ~n1795 & n1796 ;
  assign n1798 = ~n1715 & n1717 ;
  assign n1799 = n1718 | n1798 ;
  assign n1800 = ~n1797 & n1799 ;
  assign n1801 = n1797 & ~n1799 ;
  assign n1802 = n1800 | n1801 ;
  assign n1803 = ~n1791 & n1802 ;
  assign n1804 = n903 & n1377 ;
  assign n1805 = n696 & ~n1377 ;
  assign n1806 = ~n1025 & n1805 ;
  assign n1807 = n1025 & ~n1805 ;
  assign n1808 = n1806 | n1807 ;
  assign n1809 = n1804 | n1808 ;
  assign n1810 = n779 & n1252 ;
  assign n1811 = ~n779 & n1258 ;
  assign n1812 = n1082 | n1256 ;
  assign n1813 = n1082 & ~n1254 ;
  assign n1814 = n1812 & ~n1813 ;
  assign n1815 = ~n1811 & n1814 ;
  assign n1816 = ~n1810 & n1815 ;
  assign n1817 = ~n1809 & n1816 ;
  assign n1818 = n1809 & ~n1816 ;
  assign n1819 = n1817 | n1818 ;
  assign n1820 = n1158 & n1199 ;
  assign n1821 = n1100 | n1199 ;
  assign n1822 = n1156 & ~n1248 ;
  assign n1823 = n1098 & n1248 ;
  assign n1824 = n1822 | n1823 ;
  assign n1825 = n1821 & ~n1824 ;
  assign n1826 = ~n1820 & n1825 ;
  assign n1827 = ~n1819 & n1826 ;
  assign n1828 = n1817 | n1827 ;
  assign n1829 = ~n1766 & n1773 ;
  assign n1830 = n1774 | n1829 ;
  assign n1831 = n1828 & ~n1830 ;
  assign n1832 = ~n1828 & n1830 ;
  assign n1833 = n1831 | n1832 ;
  assign n1834 = n1748 | n1755 ;
  assign n1835 = ~n1756 & n1834 ;
  assign n1836 = ~n1833 & n1835 ;
  assign n1837 = n1831 | n1836 ;
  assign n1838 = ~n1787 & n1789 ;
  assign n1839 = n1790 | n1838 ;
  assign n1840 = ~n1837 & n1839 ;
  assign n1841 = n688 | n1765 ;
  assign n1842 = ~n1766 & n1841 ;
  assign n1843 = n779 | n1025 ;
  assign n1844 = n1377 & n1843 ;
  assign n1845 = n903 & n1025 ;
  assign n1846 = n903 | n1025 ;
  assign n1847 = ~n1377 & n1846 ;
  assign n1848 = ~n1845 & n1847 ;
  assign n1849 = n1844 | n1848 ;
  assign n1850 = n1158 & n1339 ;
  assign n1851 = n896 & ~n1850 ;
  assign n1852 = ~n1156 & n1851 ;
  assign n1853 = ~n1849 & n1852 ;
  assign n1854 = n1842 & n1853 ;
  assign n1855 = n1842 | n1853 ;
  assign n1856 = ~n1854 & n1855 ;
  assign n1857 = n1158 & n1248 ;
  assign n1858 = n1100 | n1248 ;
  assign n1859 = n1156 & ~n1339 ;
  assign n1860 = n1098 & n1339 ;
  assign n1861 = n1859 | n1860 ;
  assign n1862 = n1858 & ~n1861 ;
  assign n1863 = ~n1857 & n1862 ;
  assign n1864 = n1199 | n1256 ;
  assign n1865 = ~n1082 & n1258 ;
  assign n1866 = n1864 & ~n1865 ;
  assign n1867 = n1082 & n1252 ;
  assign n1868 = n1199 & ~n1254 ;
  assign n1869 = n1867 | n1868 ;
  assign n1870 = n1866 & ~n1869 ;
  assign n1871 = n1863 & n1870 ;
  assign n1872 = n1863 | n1870 ;
  assign n1873 = n1849 & ~n1852 ;
  assign n1874 = n1853 | n1873 ;
  assign n1875 = n1872 & ~n1874 ;
  assign n1876 = n1871 | n1875 ;
  assign n1877 = n1856 & n1876 ;
  assign n1878 = n1854 | n1877 ;
  assign n1879 = n1833 & ~n1835 ;
  assign n1880 = n1836 | n1879 ;
  assign n1881 = ~n1878 & n1880 ;
  assign n1882 = n1840 | n1881 ;
  assign n1883 = n1856 | n1876 ;
  assign n1884 = ~n1877 & n1883 ;
  assign n1885 = ~n1871 & n1872 ;
  assign n1886 = n1874 & n1885 ;
  assign n1887 = n1874 | n1885 ;
  assign n1888 = ~n1886 & n1887 ;
  assign n1889 = n1025 | n1082 ;
  assign n1890 = n1377 & n1889 ;
  assign n1891 = n779 & n1025 ;
  assign n1892 = n1843 & ~n1891 ;
  assign n1893 = ~n1377 & n1892 ;
  assign n1894 = n1890 | n1893 ;
  assign n1895 = n1248 | n1256 ;
  assign n1896 = n1248 & ~n1254 ;
  assign n1897 = n1895 & ~n1896 ;
  assign n1898 = n1199 & n1252 ;
  assign n1899 = ~n1199 & n1258 ;
  assign n1900 = n1898 | n1899 ;
  assign n1901 = n1897 & ~n1900 ;
  assign n1902 = ~n1894 & n1901 ;
  assign n1903 = n1204 & n1339 ;
  assign n1904 = n1078 & ~n1903 ;
  assign n1905 = n1025 | n1199 ;
  assign n1906 = n1377 & n1905 ;
  assign n1907 = n1025 & n1082 ;
  assign n1908 = n1377 | n1907 ;
  assign n1909 = n1889 & ~n1908 ;
  assign n1910 = n1906 | n1909 ;
  assign n1911 = n1904 & ~n1910 ;
  assign n1912 = n1894 & ~n1901 ;
  assign n1913 = n1902 | n1912 ;
  assign n1914 = n1911 & ~n1913 ;
  assign n1915 = n1902 | n1914 ;
  assign n1916 = n1888 & ~n1915 ;
  assign n1917 = ~n1888 & n1915 ;
  assign n1918 = ~n1904 & n1910 ;
  assign n1919 = n1911 | n1918 ;
  assign n1920 = n1199 & ~n1377 ;
  assign n1921 = n1025 & n1920 ;
  assign n1922 = n1248 & n1377 ;
  assign n1923 = n1025 | n1922 ;
  assign n1924 = n1920 | n1923 ;
  assign n1925 = ~n1921 & n1924 ;
  assign n1926 = n1248 & ~n1377 ;
  assign n1927 = n1339 | n1926 ;
  assign n1928 = n1920 | n1927 ;
  assign n1929 = ~n1903 & n1928 ;
  assign n1930 = n1925 | n1929 ;
  assign n1931 = n1919 & n1930 ;
  assign n1932 = n1919 | n1930 ;
  assign n1933 = n1256 | n1339 ;
  assign n1934 = ~n1248 & n1258 ;
  assign n1935 = n1248 & n1252 ;
  assign n1936 = ~n1254 & n1339 ;
  assign n1937 = n1935 | n1936 ;
  assign n1938 = n1934 | n1937 ;
  assign n1939 = n1933 & ~n1938 ;
  assign n1940 = n1932 & ~n1939 ;
  assign n1941 = n1931 | n1940 ;
  assign n1942 = ~n1097 & n1339 ;
  assign n1943 = ~n1941 & n1942 ;
  assign n1944 = n1917 | n1943 ;
  assign n1945 = n1941 & ~n1942 ;
  assign n1946 = ~n1911 & n1913 ;
  assign n1947 = n1914 | n1946 ;
  assign n1948 = n1945 | n1947 ;
  assign n1949 = ~n1944 & n1948 ;
  assign n1950 = n1916 | n1949 ;
  assign n1951 = n1884 & ~n1950 ;
  assign n1952 = n1878 & ~n1880 ;
  assign n1953 = ~n1884 & n1950 ;
  assign n1954 = n1819 & ~n1826 ;
  assign n1955 = n1827 | n1954 ;
  assign n1956 = n1953 | n1955 ;
  assign n1957 = ~n1952 & n1956 ;
  assign n1958 = ~n1951 & n1957 ;
  assign n1959 = n1882 | n1958 ;
  assign n1960 = n1791 & ~n1802 ;
  assign n1961 = n1837 & ~n1839 ;
  assign n1962 = n1960 | n1961 ;
  assign n1963 = n1959 & ~n1962 ;
  assign n1964 = n1803 | n1963 ;
  assign n1965 = n1795 | n1801 ;
  assign n1966 = n1964 & ~n1965 ;
  assign n1967 = ~n1964 & n1965 ;
  assign n1968 = ~n1663 & n1722 ;
  assign n1969 = n1724 & ~n1968 ;
  assign n1970 = n1726 | n1969 ;
  assign n1971 = ~n1967 & n1970 ;
  assign n1972 = n1966 | n1971 ;
  assign n1973 = n1731 | n1972 ;
  assign n1974 = ~n1730 & n1973 ;
  assign n1975 = n1678 | n1974 ;
  assign n1976 = ~n1676 & n1975 ;
  assign n1977 = ~n1621 & n1623 ;
  assign n1978 = n1624 | n1977 ;
  assign n1979 = n1976 | n1978 ;
  assign n1980 = ~n1624 & n1979 ;
  assign n1981 = n1552 | n1980 ;
  assign n1982 = ~n1550 & n1981 ;
  assign n1983 = n1433 | n1439 ;
  assign n1984 = ~n1507 & n1983 ;
  assign n1985 = n1509 | n1984 ;
  assign n1986 = n1982 | n1985 ;
  assign n1987 = ~n1509 & n1986 ;
  assign n1988 = ~n1434 & n1436 ;
  assign n1989 = n1437 | n1988 ;
  assign n1990 = n1987 | n1989 ;
  assign n1991 = ~n1437 & n1990 ;
  assign n1992 = ~n1315 & n1317 ;
  assign n1993 = n1318 | n1992 ;
  assign n1994 = n1991 | n1993 ;
  assign n1995 = ~n1318 & n1994 ;
  assign n1996 = ~n1180 & n1182 ;
  assign n1997 = n1183 | n1996 ;
  assign n1998 = n1995 | n1997 ;
  assign n1999 = ~n1183 & n1998 ;
  assign n2000 = ~n1130 & n1132 ;
  assign n2001 = n1133 | n2000 ;
  assign n2002 = n1999 | n2001 ;
  assign n2003 = ~n1133 & n2002 ;
  assign n2004 = n954 | n2003 ;
  assign n2005 = ~n952 & n2004 ;
  assign n2006 = n764 | n2005 ;
  assign n2007 = ~n762 & n2006 ;
  assign n2008 = ~n580 & n582 ;
  assign n2009 = n583 | n2008 ;
  assign n2010 = n2007 | n2009 ;
  assign n2011 = ~n583 & n2010 ;
  assign n2012 = n44 | n221 ;
  assign n2013 = n44 & n221 ;
  assign n2014 = n2012 & ~n2013 ;
  assign n2015 = n349 & ~n2014 ;
  assign n2016 = ~n349 & n2014 ;
  assign n2017 = n2015 | n2016 ;
  assign n2018 = n216 & ~n2017 ;
  assign n2019 = ~n2011 & n2018 ;
  assign n2020 = n583 | n2018 ;
  assign n2021 = n2010 & ~n2020 ;
  assign n2022 = n2019 | n2021 ;
  assign n2023 = ~n541 & n2022 ;
  assign n2024 = n541 & ~n2021 ;
  assign n2025 = ~n2019 & n2024 ;
  assign n2026 = n2023 | n2025 ;
  assign n2027 = n112 | n618 ;
  assign n2028 = n142 | n229 ;
  assign n2029 = n260 | n2028 ;
  assign n2030 = n390 | n1028 ;
  assign n2031 = n2029 | n2030 ;
  assign n2032 = n270 | n459 ;
  assign n2033 = n177 | n2032 ;
  assign n2034 = n192 | n2033 ;
  assign n2035 = n293 | n2034 ;
  assign n2036 = n2031 | n2035 ;
  assign n2037 = n224 | n2036 ;
  assign n2038 = n173 | n400 ;
  assign n2039 = n2037 | n2038 ;
  assign n2040 = n189 | n2039 ;
  assign n2041 = n292 | n2040 ;
  assign n2042 = n143 | n650 ;
  assign n2043 = n2041 | n2042 ;
  assign n2044 = n2027 | n2043 ;
  assign n2045 = n419 | n2044 ;
  assign n2046 = n198 | n398 ;
  assign n2047 = n132 | n254 ;
  assign n2048 = n445 | n2047 ;
  assign n2049 = n226 | n2048 ;
  assign n2050 = n2046 | n2049 ;
  assign n2051 = n182 | n193 ;
  assign n2052 = n149 | n2051 ;
  assign n2053 = n318 | n2052 ;
  assign n2054 = n114 | n2053 ;
  assign n2055 = n2050 | n2054 ;
  assign n2056 = n2045 | n2055 ;
  assign n2057 = ~n807 & n825 ;
  assign n2058 = n162 | n204 ;
  assign n2059 = n2057 & ~n2058 ;
  assign n2060 = ~n2056 & n2059 ;
  assign n2061 = ~n992 & n2060 ;
  assign n2062 = n2026 & n2061 ;
  assign n2063 = n2007 & n2009 ;
  assign n2064 = n2010 & ~n2063 ;
  assign n2065 = n162 | n265 ;
  assign n2066 = n137 | n2065 ;
  assign n2067 = n191 | n332 ;
  assign n2068 = n2066 | n2067 ;
  assign n2069 = n253 | n445 ;
  assign n2070 = n154 | n183 ;
  assign n2071 = n279 | n398 ;
  assign n2072 = n248 | n315 ;
  assign n2073 = n254 | n2072 ;
  assign n2074 = n2071 | n2073 ;
  assign n2075 = n187 | n2074 ;
  assign n2076 = n2070 | n2075 ;
  assign n2077 = n313 | n480 ;
  assign n2078 = n268 | n659 ;
  assign n2079 = n2077 | n2078 ;
  assign n2080 = n2076 | n2079 ;
  assign n2081 = n584 | n2080 ;
  assign n2082 = n325 | n444 ;
  assign n2083 = n400 | n2082 ;
  assign n2084 = n134 | n383 ;
  assign n2085 = n240 | n2084 ;
  assign n2086 = n272 | n2085 ;
  assign n2087 = n247 | n501 ;
  assign n2088 = n112 | n326 ;
  assign n2089 = n470 | n2088 ;
  assign n2090 = n867 | n973 ;
  assign n2091 = n2089 | n2090 ;
  assign n2092 = n2087 | n2091 ;
  assign n2093 = n2086 | n2092 ;
  assign n2094 = n2083 | n2093 ;
  assign n2095 = n2081 | n2094 ;
  assign n2096 = n309 | n327 ;
  assign n2097 = n125 | n288 ;
  assign n2098 = n2096 | n2097 ;
  assign n2099 = n206 | n594 ;
  assign n2100 = n290 | n2099 ;
  assign n2101 = n148 | n2100 ;
  assign n2102 = n2098 | n2101 ;
  assign n2103 = n496 | n2102 ;
  assign n2104 = n146 | n613 ;
  assign n2105 = n199 | n2104 ;
  assign n2106 = n2103 | n2105 ;
  assign n2107 = n679 | n2106 ;
  assign n2108 = n2095 | n2107 ;
  assign n2109 = n2069 | n2108 ;
  assign n2110 = n2068 | n2109 ;
  assign n2111 = n260 | n389 ;
  assign n2112 = n2110 | n2111 ;
  assign n2113 = ~n2064 & n2112 ;
  assign n2114 = n764 & n2005 ;
  assign n2115 = n2006 & ~n2114 ;
  assign n2116 = n510 | n984 ;
  assign n2117 = n272 | n315 ;
  assign n2118 = n2116 | n2117 ;
  assign n2119 = n431 | n634 ;
  assign n2120 = n588 | n810 ;
  assign n2121 = n803 | n2120 ;
  assign n2122 = n241 | n2121 ;
  assign n2123 = n2119 | n2122 ;
  assign n2124 = n853 | n2123 ;
  assign n2125 = n395 | n2124 ;
  assign n2126 = n226 | n2125 ;
  assign n2127 = n288 | n2126 ;
  assign n2128 = n2118 | n2127 ;
  assign n2129 = ~n2115 & n2128 ;
  assign n2130 = n954 & n2003 ;
  assign n2131 = n2004 & ~n2130 ;
  assign n2132 = n201 | n313 ;
  assign n2133 = n237 | n310 ;
  assign n2134 = n617 | n2133 ;
  assign n2135 = n139 | n396 ;
  assign n2136 = n459 | n2135 ;
  assign n2137 = n2134 | n2136 ;
  assign n2138 = n431 | n2066 ;
  assign n2139 = n2048 | n2089 ;
  assign n2140 = n2138 | n2139 ;
  assign n2141 = n2137 | n2140 ;
  assign n2142 = n2132 | n2141 ;
  assign n2143 = n236 | n328 ;
  assign n2144 = n178 | n2143 ;
  assign n2145 = n378 | n2144 ;
  assign n2146 = n250 | n2038 ;
  assign n2147 = n2145 | n2146 ;
  assign n2148 = n279 | n809 ;
  assign n2149 = n267 | n309 ;
  assign n2150 = n2148 | n2149 ;
  assign n2151 = n500 | n2150 ;
  assign n2152 = n266 | n2151 ;
  assign n2153 = n485 | n632 ;
  assign n2154 = n2152 | n2153 ;
  assign n2155 = n155 | n176 ;
  assign n2156 = n385 | n2155 ;
  assign n2157 = n2154 | n2156 ;
  assign n2158 = n114 | n386 ;
  assign n2159 = n402 | n2158 ;
  assign n2160 = n2157 | n2159 ;
  assign n2161 = n202 | n231 ;
  assign n2162 = n331 | n2161 ;
  assign n2163 = n491 | n2162 ;
  assign n2164 = n2160 | n2163 ;
  assign n2165 = n2147 | n2164 ;
  assign n2166 = n2142 | n2165 ;
  assign n2167 = ~n2131 & n2166 ;
  assign n2168 = n2131 & ~n2166 ;
  assign n2169 = n2167 | n2168 ;
  assign n2170 = n110 & n136 ;
  assign n2171 = n187 | n202 ;
  assign n2172 = n165 | n859 ;
  assign n2173 = n267 | n510 ;
  assign n2174 = n374 | n2173 ;
  assign n2175 = n2172 | n2174 ;
  assign n2176 = n194 | n275 ;
  assign n2177 = n2144 | n2176 ;
  assign n2178 = n410 | n2177 ;
  assign n2179 = n205 | n2178 ;
  assign n2180 = n311 | n318 ;
  assign n2181 = n260 | n2180 ;
  assign n2182 = n2179 | n2181 ;
  assign n2183 = n380 | n2182 ;
  assign n2184 = n2103 | n2183 ;
  assign n2185 = n230 | n389 ;
  assign n2186 = n145 | n2185 ;
  assign n2187 = n2142 | n2186 ;
  assign n2188 = n825 & ~n2187 ;
  assign n2189 = ~n1347 & n2188 ;
  assign n2190 = ~n2184 & n2189 ;
  assign n2191 = ~n2175 & n2190 ;
  assign n2192 = ~n2171 & n2191 ;
  assign n2193 = ~n2170 & n2192 ;
  assign n2194 = ~n1183 & n2001 ;
  assign n2195 = n1998 & n2194 ;
  assign n2196 = n2002 & ~n2195 ;
  assign n2197 = n2193 | n2196 ;
  assign n2198 = n174 | n274 ;
  assign n2199 = n231 | n2198 ;
  assign n2200 = n137 | n445 ;
  assign n2201 = n176 | n310 ;
  assign n2202 = n119 | n2201 ;
  assign n2203 = n161 | n327 ;
  assign n2204 = n2202 | n2203 ;
  assign n2205 = n243 | n2204 ;
  assign n2206 = n226 | n333 ;
  assign n2207 = n2205 | n2206 ;
  assign n2208 = n191 | n227 ;
  assign n2209 = n270 | n379 ;
  assign n2210 = n245 | n2209 ;
  assign n2211 = n2208 | n2210 ;
  assign n2212 = n252 | n823 ;
  assign n2213 = n398 | n2212 ;
  assign n2214 = n193 | n2028 ;
  assign n2215 = n207 | n378 ;
  assign n2216 = n1010 | n2215 ;
  assign n2217 = n2214 | n2216 ;
  assign n2218 = n840 | n2217 ;
  assign n2219 = n288 | n2218 ;
  assign n2220 = n267 | n290 ;
  assign n2221 = n2219 | n2220 ;
  assign n2222 = n2213 | n2221 ;
  assign n2223 = n2211 | n2222 ;
  assign n2224 = n2207 | n2223 ;
  assign n2225 = n126 | n2224 ;
  assign n2226 = n2200 | n2225 ;
  assign n2227 = n325 | n2226 ;
  assign n2228 = n2199 | n2227 ;
  assign n2229 = n1995 & n1997 ;
  assign n2230 = n1998 & ~n2229 ;
  assign n2231 = n2228 & ~n2230 ;
  assign n2232 = n145 | n165 ;
  assign n2233 = n183 | n650 ;
  assign n2234 = n2232 | n2233 ;
  assign n2235 = n339 | n398 ;
  assign n2236 = n227 | n338 ;
  assign n2237 = n790 | n813 ;
  assign n2238 = n668 | n2237 ;
  assign n2239 = n2236 | n2238 ;
  assign n2240 = n2235 | n2239 ;
  assign n2241 = n119 | n270 ;
  assign n2242 = n252 | n291 ;
  assign n2243 = n500 | n2242 ;
  assign n2244 = n175 | n2243 ;
  assign n2245 = n2241 | n2244 ;
  assign n2246 = n203 | n419 ;
  assign n2247 = n2245 | n2246 ;
  assign n2248 = n1036 | n2247 ;
  assign n2249 = n2240 | n2248 ;
  assign n2250 = n260 | n2249 ;
  assign n2251 = n243 | n787 ;
  assign n2252 = n2250 | n2251 ;
  assign n2253 = n2234 | n2252 ;
  assign n2254 = n301 | n584 ;
  assign n2255 = n271 | n862 ;
  assign n2256 = n121 | n2255 ;
  assign n2257 = n2254 | n2256 ;
  assign n2258 = n441 | n783 ;
  assign n2259 = n224 | n445 ;
  assign n2260 = n2258 | n2259 ;
  assign n2261 = n330 | n333 ;
  assign n2262 = n480 | n867 ;
  assign n2263 = n2261 | n2262 ;
  assign n2264 = n2260 | n2263 ;
  assign n2265 = n2257 | n2264 ;
  assign n2266 = n2253 | n2265 ;
  assign n2267 = n245 | n2266 ;
  assign n2268 = n314 | n2267 ;
  assign n2269 = n1991 & n1993 ;
  assign n2270 = n1994 & ~n2269 ;
  assign n2271 = n2268 & ~n2270 ;
  assign n2272 = n187 | n430 ;
  assign n2273 = n290 | n2272 ;
  assign n2274 = n198 | n386 ;
  assign n2275 = n174 | n510 ;
  assign n2276 = n500 | n2275 ;
  assign n2277 = n2274 | n2276 ;
  assign n2278 = n230 | n273 ;
  assign n2279 = n132 | n2278 ;
  assign n2280 = n374 | n2279 ;
  assign n2281 = n2277 | n2280 ;
  assign n2282 = n149 | n340 ;
  assign n2283 = n244 | n291 ;
  assign n2284 = n254 | n2283 ;
  assign n2285 = n811 | n2284 ;
  assign n2286 = n2282 | n2285 ;
  assign n2287 = n269 | n2082 ;
  assign n2288 = n2040 | n2287 ;
  assign n2289 = n2286 | n2288 ;
  assign n2290 = n2281 | n2289 ;
  assign n2291 = n181 | n207 ;
  assign n2292 = n155 | n2291 ;
  assign n2293 = n202 | n278 ;
  assign n2294 = n496 | n2293 ;
  assign n2295 = n2292 | n2294 ;
  assign n2296 = n237 | n2295 ;
  assign n2297 = n201 | n396 ;
  assign n2298 = n2296 | n2297 ;
  assign n2299 = n2290 | n2298 ;
  assign n2300 = n2273 | n2299 ;
  assign n2301 = n261 | n2300 ;
  assign n2302 = n1987 & n1989 ;
  assign n2303 = n1990 & ~n2302 ;
  assign n2304 = n2301 & ~n2303 ;
  assign n2305 = n386 | n618 ;
  assign n2306 = n248 | n2305 ;
  assign n2307 = n137 | n310 ;
  assign n2308 = n867 | n2307 ;
  assign n2309 = n463 | n2308 ;
  assign n2310 = n2306 | n2309 ;
  assign n2311 = n260 | n278 ;
  assign n2312 = n135 | n255 ;
  assign n2313 = n317 | n2312 ;
  assign n2314 = n325 | n2313 ;
  assign n2315 = n2311 | n2314 ;
  assign n2316 = n481 | n2315 ;
  assign n2317 = n809 | n2162 ;
  assign n2318 = n514 | n2317 ;
  assign n2319 = n128 | n2318 ;
  assign n2320 = n294 | n2319 ;
  assign n2321 = n224 | n2320 ;
  assign n2322 = n2235 | n2321 ;
  assign n2323 = n2316 | n2322 ;
  assign n2324 = n637 | n2323 ;
  assign n2325 = n183 | n644 ;
  assign n2326 = n114 | n631 ;
  assign n2327 = n2325 | n2326 ;
  assign n2328 = n2324 | n2327 ;
  assign n2329 = n2310 | n2328 ;
  assign n2330 = n230 | n2329 ;
  assign n2331 = n191 | n2330 ;
  assign n2332 = n1982 & n1985 ;
  assign n2333 = n1986 & ~n2332 ;
  assign n2334 = n2331 & ~n2333 ;
  assign n2335 = n390 | n2174 ;
  assign n2336 = n249 | n318 ;
  assign n2337 = n266 | n1344 ;
  assign n2338 = n2336 | n2337 ;
  assign n2339 = n882 | n2338 ;
  assign n2340 = n2278 | n2339 ;
  assign n2341 = n2335 | n2340 ;
  assign n2342 = n261 | n2341 ;
  assign n2343 = n301 | n330 ;
  assign n2344 = n584 | n650 ;
  assign n2345 = n2343 | n2344 ;
  assign n2346 = n2342 | n2345 ;
  assign n2347 = n315 | n787 ;
  assign n2348 = n224 | n2347 ;
  assign n2349 = n311 | n2348 ;
  assign n2350 = n2346 | n2349 ;
  assign n2351 = n332 | n397 ;
  assign n2352 = n194 | n2351 ;
  assign n2353 = n614 | n2352 ;
  assign n2354 = n2315 | n2353 ;
  assign n2355 = n2057 & ~n2354 ;
  assign n2356 = ~n474 & n2355 ;
  assign n2357 = ~n862 & n2356 ;
  assign n2358 = ~n2350 & n2357 ;
  assign n2359 = ~n445 & n2358 ;
  assign n2360 = ~n112 & n2359 ;
  assign n2361 = ~n1015 & n2360 ;
  assign n2362 = ~n500 & n2361 ;
  assign n2363 = n1552 & n1980 ;
  assign n2364 = n1981 & ~n2363 ;
  assign n2365 = n2362 | n2364 ;
  assign n2366 = n188 | n278 ;
  assign n2367 = n231 | n2366 ;
  assign n2368 = n374 | n400 ;
  assign n2369 = n441 | n2278 ;
  assign n2370 = n241 | n2369 ;
  assign n2371 = n181 | n326 ;
  assign n2372 = n293 | n2371 ;
  assign n2373 = n165 | n2372 ;
  assign n2374 = n444 | n2373 ;
  assign n2375 = n290 | n386 ;
  assign n2376 = n2374 | n2375 ;
  assign n2377 = n2370 | n2376 ;
  assign n2378 = n145 | n176 ;
  assign n2379 = n1011 | n2378 ;
  assign n2380 = n283 | n288 ;
  assign n2381 = n311 | n2380 ;
  assign n2382 = n2240 | n2381 ;
  assign n2383 = n2379 | n2382 ;
  assign n2384 = n2377 | n2383 ;
  assign n2385 = n2368 | n2384 ;
  assign n2386 = n163 | n2385 ;
  assign n2387 = n204 | n2386 ;
  assign n2388 = n611 | n2387 ;
  assign n2389 = n327 | n2388 ;
  assign n2390 = n2367 | n2389 ;
  assign n2391 = n193 | n2390 ;
  assign n2392 = n1976 & n1978 ;
  assign n2393 = n1979 & ~n2392 ;
  assign n2394 = n2391 & ~n2393 ;
  assign n2395 = n155 | n2094 ;
  assign n2396 = n390 | n800 ;
  assign n2397 = n648 | n976 ;
  assign n2398 = n2396 | n2397 ;
  assign n2399 = n2395 | n2398 ;
  assign n2400 = n634 | n2322 ;
  assign n2401 = n268 | n315 ;
  assign n2402 = n188 | n2401 ;
  assign n2403 = n2400 | n2402 ;
  assign n2404 = n2399 | n2403 ;
  assign n2405 = n380 | n2404 ;
  assign n2406 = n1678 & n1974 ;
  assign n2407 = n1975 & ~n2406 ;
  assign n2408 = ~n2405 & n2407 ;
  assign n2409 = ~n2391 & n2393 ;
  assign n2410 = n2394 | n2409 ;
  assign n2411 = n2408 | n2410 ;
  assign n2412 = ~n2394 & n2411 ;
  assign n2413 = n2362 & n2364 ;
  assign n2414 = n2365 & ~n2413 ;
  assign n2415 = ~n2412 & n2414 ;
  assign n2416 = n2365 & ~n2415 ;
  assign n2417 = ~n2331 & n2333 ;
  assign n2418 = n2334 | n2417 ;
  assign n2419 = n2416 | n2418 ;
  assign n2420 = ~n2334 & n2419 ;
  assign n2421 = ~n2301 & n2303 ;
  assign n2422 = n2304 | n2421 ;
  assign n2423 = n2420 | n2422 ;
  assign n2424 = ~n2304 & n2423 ;
  assign n2425 = ~n2268 & n2270 ;
  assign n2426 = n2271 | n2425 ;
  assign n2427 = n2424 | n2426 ;
  assign n2428 = ~n2271 & n2427 ;
  assign n2429 = ~n2228 & n2230 ;
  assign n2430 = n2231 | n2429 ;
  assign n2431 = n2428 | n2430 ;
  assign n2432 = ~n2231 & n2431 ;
  assign n2433 = n2193 & n2196 ;
  assign n2434 = n2197 & ~n2433 ;
  assign n2435 = ~n2432 & n2434 ;
  assign n2436 = n2197 & ~n2435 ;
  assign n2437 = n2169 | n2436 ;
  assign n2438 = ~n2167 & n2437 ;
  assign n2439 = n2115 & ~n2128 ;
  assign n2440 = n2129 | n2439 ;
  assign n2441 = n2438 | n2440 ;
  assign n2442 = ~n2129 & n2441 ;
  assign n2443 = n2064 & ~n2112 ;
  assign n2444 = n2113 | n2443 ;
  assign n2445 = n2442 | n2444 ;
  assign n2446 = ~n2113 & n2445 ;
  assign n2447 = n2025 | n2061 ;
  assign n2448 = n2023 | n2447 ;
  assign n2449 = ~n2446 & n2448 ;
  assign n2450 = ~n2062 & n2449 ;
  assign n2451 = n149 | n162 ;
  assign n2452 = n176 | n192 ;
  assign n2453 = n2451 | n2452 ;
  assign n2454 = n178 | n281 ;
  assign n2455 = n126 | n2454 ;
  assign n2456 = n229 | n2455 ;
  assign n2457 = n2453 | n2456 ;
  assign n2458 = n250 | n973 ;
  assign n2459 = n2240 | n2458 ;
  assign n2460 = n2457 | n2459 ;
  assign n2461 = n1356 | n2460 ;
  assign n2462 = n463 | n2461 ;
  assign n2463 = n450 | n2462 ;
  assign n2464 = n826 | n2463 ;
  assign n2465 = n386 | n2464 ;
  assign n2466 = n1057 | n2465 ;
  assign n2467 = n224 | n2466 ;
  assign n2468 = n2448 & ~n2467 ;
  assign n2469 = ~n2450 & n2468 ;
  assign n2470 = n148 | n165 ;
  assign n2471 = n374 | n660 ;
  assign n2472 = n667 | n2471 ;
  assign n2473 = n2470 | n2472 ;
  assign n2474 = n176 | n661 ;
  assign n2475 = n112 | n2474 ;
  assign n2476 = n315 | n339 ;
  assign n2477 = n293 | n2476 ;
  assign n2478 = n287 | n398 ;
  assign n2479 = n613 | n2478 ;
  assign n2480 = n134 | n183 ;
  assign n2481 = n188 | n2066 ;
  assign n2482 = n244 | n268 ;
  assign n2483 = n174 | n430 ;
  assign n2484 = n2482 | n2483 ;
  assign n2485 = n2481 | n2484 ;
  assign n2486 = n2480 | n2485 ;
  assign n2487 = n2479 | n2486 ;
  assign n2488 = n301 | n2487 ;
  assign n2489 = n318 | n2488 ;
  assign n2490 = n267 | n2489 ;
  assign n2491 = n2477 | n2490 ;
  assign n2492 = n204 | n313 ;
  assign n2493 = n642 | n2492 ;
  assign n2494 = n2491 | n2493 ;
  assign n2495 = n2475 | n2494 ;
  assign n2496 = n132 | n386 ;
  assign n2497 = n273 | n2496 ;
  assign n2498 = n189 | n2497 ;
  assign n2499 = n253 | n444 ;
  assign n2500 = n2498 | n2499 ;
  assign n2501 = n149 | n237 ;
  assign n2502 = n154 | n282 ;
  assign n2503 = n2501 | n2502 ;
  assign n2504 = n2500 | n2503 ;
  assign n2505 = n191 | n400 ;
  assign n2506 = n119 | n291 ;
  assign n2507 = n2505 | n2506 ;
  assign n2508 = n197 | n248 ;
  assign n2509 = n173 | n252 ;
  assign n2510 = n2508 | n2509 ;
  assign n2511 = n2507 | n2510 ;
  assign n2512 = n2504 | n2511 ;
  assign n2513 = n2495 | n2512 ;
  assign n2514 = n2473 | n2513 ;
  assign n2515 = n326 | n2514 ;
  assign n2516 = n121 | n143 ;
  assign n2517 = n249 | n302 ;
  assign n2518 = n2516 | n2517 ;
  assign n2519 = n2515 | n2518 ;
  assign n2520 = n2469 & ~n2519 ;
  assign n2521 = n855 | n1344 ;
  assign n2522 = ~n619 & n824 ;
  assign n2523 = n172 | n263 ;
  assign n2524 = n2522 & ~n2523 ;
  assign n2525 = ~n2152 & n2524 ;
  assign n2526 = ~n272 & n2525 ;
  assign n2527 = ~n332 & n2526 ;
  assign n2528 = ~n2521 & n2527 ;
  assign n2529 = ~n2345 & n2528 ;
  assign n2530 = ~n281 & n2529 ;
  assign n2531 = ~n510 & n2530 ;
  assign n2532 = ~n618 & n2531 ;
  assign n2533 = n2520 & n2532 ;
  assign n2534 = n118 | n162 ;
  assign n2535 = n277 | n2534 ;
  assign n2536 = n292 | n1049 ;
  assign n2537 = n157 | n2536 ;
  assign n2538 = n2535 | n2537 ;
  assign n2539 = n186 | n199 ;
  assign n2540 = n203 | n324 ;
  assign n2541 = n263 | n2540 ;
  assign n2542 = n2539 | n2541 ;
  assign n2543 = n2538 | n2542 ;
  assign n2544 = n206 | n2543 ;
  assign n2545 = n2533 | n2544 ;
  assign n2546 = n2533 & n2544 ;
  assign n2547 = n2545 & ~n2546 ;
  assign n2548 = n2520 | n2532 ;
  assign n2549 = ~n2533 & n2548 ;
  assign n2550 = n2547 & ~n2549 ;
  assign n2551 = n2469 | n2519 ;
  assign n2552 = n2469 & n2519 ;
  assign n2553 = n2551 & ~n2552 ;
  assign n2554 = ~n2549 & n2553 ;
  assign n2555 = n2448 & ~n2450 ;
  assign n2556 = n2467 & ~n2555 ;
  assign n2557 = n2469 | n2556 ;
  assign n2558 = n2553 & n2557 ;
  assign n2559 = ~n2062 & n2448 ;
  assign n2560 = n2446 & ~n2559 ;
  assign n2561 = n2450 | n2560 ;
  assign n2562 = n2557 & ~n2561 ;
  assign n2563 = n2442 & n2444 ;
  assign n2564 = n2445 & ~n2563 ;
  assign n2565 = ~n2561 & n2564 ;
  assign n2566 = n2561 & ~n2564 ;
  assign n2567 = n2565 | n2566 ;
  assign n2568 = n2438 & n2440 ;
  assign n2569 = n2441 & ~n2568 ;
  assign n2570 = n2564 & n2569 ;
  assign n2571 = n2169 & n2436 ;
  assign n2572 = n2437 & ~n2571 ;
  assign n2573 = n2569 & n2572 ;
  assign n2574 = n2432 & ~n2434 ;
  assign n2575 = n2435 | n2574 ;
  assign n2576 = n2572 & ~n2575 ;
  assign n2577 = n2428 & n2430 ;
  assign n2578 = n2431 & ~n2577 ;
  assign n2579 = ~n2575 & n2578 ;
  assign n2580 = n2424 & n2426 ;
  assign n2581 = n2427 & ~n2580 ;
  assign n2582 = n2578 & n2581 ;
  assign n2583 = n2420 & n2422 ;
  assign n2584 = n2423 & ~n2583 ;
  assign n2585 = n2581 & n2584 ;
  assign n2586 = n2416 & n2418 ;
  assign n2587 = n2419 & ~n2586 ;
  assign n2588 = n2584 & n2587 ;
  assign n2589 = n2412 & ~n2414 ;
  assign n2590 = n2415 | n2589 ;
  assign n2591 = n2587 & ~n2590 ;
  assign n2592 = n2408 & n2410 ;
  assign n2593 = n2411 & ~n2592 ;
  assign n2594 = n2405 & ~n2407 ;
  assign n2595 = n2408 | n2594 ;
  assign n2596 = n2590 & ~n2595 ;
  assign n2597 = n2593 & ~n2596 ;
  assign n2598 = ~n2587 & n2590 ;
  assign n2599 = n2591 | n2598 ;
  assign n2600 = n2597 & ~n2599 ;
  assign n2601 = n2591 | n2600 ;
  assign n2602 = n2584 | n2587 ;
  assign n2603 = ~n2588 & n2602 ;
  assign n2604 = n2601 & n2603 ;
  assign n2605 = n2588 | n2604 ;
  assign n2606 = n2581 | n2584 ;
  assign n2607 = ~n2585 & n2606 ;
  assign n2608 = n2605 & n2607 ;
  assign n2609 = n2585 | n2608 ;
  assign n2610 = n2578 | n2581 ;
  assign n2611 = ~n2582 & n2610 ;
  assign n2612 = n2609 & n2611 ;
  assign n2613 = n2582 | n2612 ;
  assign n2614 = n2575 & ~n2578 ;
  assign n2615 = n2579 | n2614 ;
  assign n2616 = n2613 & ~n2615 ;
  assign n2617 = n2579 | n2616 ;
  assign n2618 = ~n2572 & n2575 ;
  assign n2619 = n2576 | n2618 ;
  assign n2620 = n2617 & ~n2619 ;
  assign n2621 = n2576 | n2620 ;
  assign n2622 = n2569 | n2572 ;
  assign n2623 = ~n2573 & n2622 ;
  assign n2624 = n2621 & n2623 ;
  assign n2625 = n2573 | n2624 ;
  assign n2626 = n2564 | n2569 ;
  assign n2627 = ~n2570 & n2626 ;
  assign n2628 = n2625 & n2627 ;
  assign n2629 = n2570 | n2628 ;
  assign n2630 = ~n2567 & n2629 ;
  assign n2631 = n2565 | n2630 ;
  assign n2632 = ~n2557 & n2561 ;
  assign n2633 = n2562 | n2632 ;
  assign n2634 = n2631 & ~n2633 ;
  assign n2635 = n2562 | n2634 ;
  assign n2636 = n2553 | n2557 ;
  assign n2637 = ~n2558 & n2636 ;
  assign n2638 = n2635 & n2637 ;
  assign n2639 = n2558 | n2638 ;
  assign n2640 = n2549 & ~n2553 ;
  assign n2641 = n2554 | n2640 ;
  assign n2642 = n2639 & ~n2641 ;
  assign n2643 = n2554 | n2642 ;
  assign n2644 = ~n2547 & n2549 ;
  assign n2645 = n2550 | n2644 ;
  assign n2646 = n2643 & ~n2645 ;
  assign n2647 = n2550 | n2646 ;
  assign n2648 = n2533 & ~n2544 ;
  assign n2649 = n149 | n309 ;
  assign n2650 = n291 | n2649 ;
  assign n2651 = n343 | n2650 ;
  assign n2652 = n137 | n278 ;
  assign n2653 = n130 | n324 ;
  assign n2654 = n161 | n212 ;
  assign n2655 = n263 | n2654 ;
  assign n2656 = n2653 | n2655 ;
  assign n2657 = n2652 | n2656 ;
  assign n2658 = n2651 | n2657 ;
  assign n2659 = ~n2648 & n2658 ;
  assign n2660 = n2648 & ~n2658 ;
  assign n2661 = n2659 | n2660 ;
  assign n2662 = n2547 | n2661 ;
  assign n2663 = n2547 & n2661 ;
  assign n2664 = n2662 & ~n2663 ;
  assign n2665 = n2647 & n2664 ;
  assign n2666 = n2647 | n2664 ;
  assign n2667 = ~n2665 & n2666 ;
  assign n2668 = pi0 & ~pi22 ;
  assign n2669 = pi1 & ~n2668 ;
  assign n2670 = ~pi1 & n2668 ;
  assign n2671 = n2669 | n2670 ;
  assign n2672 = n29 & ~n2671 ;
  assign n2673 = ~n29 & n2671 ;
  assign n2674 = n2672 | n2673 ;
  assign n2675 = pi0 & n2674 ;
  assign n2676 = n2667 & n2675 ;
  assign n2677 = pi0 & ~n2674 ;
  assign n2678 = n2661 & n2677 ;
  assign n2679 = ~n25 & n2674 ;
  assign n2680 = ~n2549 & n2679 ;
  assign n2681 = ~pi0 & n2671 ;
  assign n2682 = n2547 & n2681 ;
  assign n2683 = n2680 | n2682 ;
  assign n2684 = n2678 | n2683 ;
  assign n2685 = n2676 | n2684 ;
  assign n2686 = n29 | n2685 ;
  assign n2687 = n29 & n2685 ;
  assign n2688 = n2686 & ~n2687 ;
  assign n2689 = ~n372 & n534 ;
  assign n2690 = n372 & ~n534 ;
  assign n2691 = n2689 | n2690 ;
  assign n2692 = ~n44 & n534 ;
  assign n2693 = n44 & ~n534 ;
  assign n2694 = n2692 | n2693 ;
  assign n2695 = ~n2691 & n2694 ;
  assign n2696 = n2595 & n2695 ;
  assign n2697 = ~n2014 & n2691 ;
  assign n2698 = n2593 & n2697 ;
  assign n2699 = ~n2593 & n2595 ;
  assign n2700 = n2593 & ~n2595 ;
  assign n2701 = n2699 | n2700 ;
  assign n2702 = n2014 & n2691 ;
  assign n2703 = n2701 & n2702 ;
  assign n2704 = n2698 | n2703 ;
  assign n2705 = n2696 | n2704 ;
  assign n2706 = n221 & ~n2705 ;
  assign n2707 = ~n221 & n2705 ;
  assign n2708 = n2706 | n2707 ;
  assign n2709 = n2595 & n2691 ;
  assign n2710 = n221 & ~n2709 ;
  assign n2711 = n2708 | n2710 ;
  assign n2712 = n221 & n2708 ;
  assign n2713 = ~n2709 & n2712 ;
  assign n2714 = n372 | n705 ;
  assign n2715 = n372 & n705 ;
  assign n2716 = n2714 & ~n2715 ;
  assign n2717 = ~n696 & n903 ;
  assign n2718 = n696 & ~n903 ;
  assign n2719 = n2717 | n2718 ;
  assign n2720 = n2716 & n2719 ;
  assign n2721 = n2601 | n2603 ;
  assign n2722 = ~n2604 & n2721 ;
  assign n2723 = n2720 & n2722 ;
  assign n2724 = ~n696 & n705 ;
  assign n2725 = n696 & ~n705 ;
  assign n2726 = n2724 | n2725 ;
  assign n2727 = n2719 | n2726 ;
  assign n2728 = n2716 & ~n2727 ;
  assign n2729 = ~n2590 & n2728 ;
  assign n2730 = ~n2719 & n2726 ;
  assign n2731 = n2587 & n2730 ;
  assign n2732 = ~n2716 & n2719 ;
  assign n2733 = n2584 & n2732 ;
  assign n2734 = n2731 | n2733 ;
  assign n2735 = n2729 | n2734 ;
  assign n2736 = n2723 | n2735 ;
  assign n2737 = n372 | n2736 ;
  assign n2738 = n372 & n2736 ;
  assign n2739 = n2737 & ~n2738 ;
  assign n2740 = ~n2713 & n2739 ;
  assign n2741 = n2711 & n2740 ;
  assign n2742 = n2595 & n2719 ;
  assign n2743 = n372 & ~n2742 ;
  assign n2744 = n2595 & n2730 ;
  assign n2745 = n2593 & n2732 ;
  assign n2746 = n2701 & n2720 ;
  assign n2747 = n2745 | n2746 ;
  assign n2748 = n2744 | n2747 ;
  assign n2749 = n372 & ~n2748 ;
  assign n2750 = ~n372 & n2748 ;
  assign n2751 = n2749 | n2750 ;
  assign n2752 = n2743 & n2751 ;
  assign n2753 = ~n2590 & n2732 ;
  assign n2754 = n2593 & n2730 ;
  assign n2755 = n2595 & n2728 ;
  assign n2756 = n2754 | n2755 ;
  assign n2757 = n2753 | n2756 ;
  assign n2758 = n2590 | n2700 ;
  assign n2759 = n2590 & n2700 ;
  assign n2760 = n2758 & ~n2759 ;
  assign n2761 = n2720 & ~n2760 ;
  assign n2762 = n2757 | n2761 ;
  assign n2763 = n372 | n2762 ;
  assign n2764 = n372 & n2762 ;
  assign n2765 = n2763 & ~n2764 ;
  assign n2766 = n2752 & n2765 ;
  assign n2767 = n2709 & n2766 ;
  assign n2768 = ~n2590 & n2730 ;
  assign n2769 = ~n2597 & n2599 ;
  assign n2770 = n2600 | n2769 ;
  assign n2771 = n2720 & ~n2770 ;
  assign n2772 = n2587 & n2732 ;
  assign n2773 = n2593 & n2728 ;
  assign n2774 = n2772 | n2773 ;
  assign n2775 = n2771 | n2774 ;
  assign n2776 = n2768 | n2775 ;
  assign n2777 = n372 & n2776 ;
  assign n2778 = n372 | n2776 ;
  assign n2779 = ~n2777 & n2778 ;
  assign n2780 = n2709 | n2766 ;
  assign n2781 = ~n2767 & n2780 ;
  assign n2782 = n2779 & n2781 ;
  assign n2783 = n2767 | n2782 ;
  assign n2784 = n2711 & ~n2713 ;
  assign n2785 = n2739 | n2784 ;
  assign n2786 = ~n2741 & n2785 ;
  assign n2787 = n2783 & n2786 ;
  assign n2788 = n2741 | n2787 ;
  assign n2789 = n2702 & ~n2760 ;
  assign n2790 = ~n2590 & n2697 ;
  assign n2791 = n2593 & n2695 ;
  assign n2792 = n2691 | n2694 ;
  assign n2793 = n2014 & ~n2792 ;
  assign n2794 = n2595 & n2793 ;
  assign n2795 = n2791 | n2794 ;
  assign n2796 = n2790 | n2795 ;
  assign n2797 = n2789 | n2796 ;
  assign n2798 = n221 | n2797 ;
  assign n2799 = n221 & n2797 ;
  assign n2800 = n2798 & ~n2799 ;
  assign n2801 = n2713 & n2800 ;
  assign n2802 = n2713 | n2800 ;
  assign n2803 = ~n2801 & n2802 ;
  assign n2804 = n2605 | n2607 ;
  assign n2805 = ~n2608 & n2804 ;
  assign n2806 = n2720 & n2805 ;
  assign n2807 = n2581 & n2732 ;
  assign n2808 = n2584 & n2730 ;
  assign n2809 = n2587 & n2728 ;
  assign n2810 = n2808 | n2809 ;
  assign n2811 = n2807 | n2810 ;
  assign n2812 = n2806 | n2811 ;
  assign n2813 = n372 & ~n2812 ;
  assign n2814 = ~n372 & n2812 ;
  assign n2815 = n2813 | n2814 ;
  assign n2816 = n2803 & n2815 ;
  assign n2817 = n2803 | n2815 ;
  assign n2818 = ~n2816 & n2817 ;
  assign n2819 = n2788 | n2818 ;
  assign n2820 = n2788 & n2818 ;
  assign n2821 = n2819 & ~n2820 ;
  assign n2822 = ~n2617 & n2619 ;
  assign n2823 = n2620 | n2822 ;
  assign n2824 = ~n779 & n903 ;
  assign n2825 = n779 & ~n903 ;
  assign n2826 = n2824 | n2825 ;
  assign n2827 = n1082 & ~n1199 ;
  assign n2828 = ~n1082 & n1199 ;
  assign n2829 = n2827 | n2828 ;
  assign n2830 = n2826 & n2829 ;
  assign n2831 = ~n2823 & n2830 ;
  assign n2832 = ~n2826 & n2829 ;
  assign n2833 = n2572 & n2832 ;
  assign n2834 = ~n779 & n1082 ;
  assign n2835 = n779 & ~n1082 ;
  assign n2836 = n2834 | n2835 ;
  assign n2837 = ~n2829 & n2836 ;
  assign n2838 = ~n2575 & n2837 ;
  assign n2839 = n2826 & ~n2829 ;
  assign n2840 = ~n2836 & n2839 ;
  assign n2841 = n2578 & n2840 ;
  assign n2842 = n2838 | n2841 ;
  assign n2843 = n2833 | n2842 ;
  assign n2844 = n2831 | n2843 ;
  assign n2845 = n903 | n2844 ;
  assign n2846 = n903 & n2844 ;
  assign n2847 = n2845 & ~n2846 ;
  assign n2848 = n2821 & n2847 ;
  assign n2849 = n2783 | n2786 ;
  assign n2850 = ~n2787 & n2849 ;
  assign n2851 = ~n2613 & n2615 ;
  assign n2852 = n2616 | n2851 ;
  assign n2853 = n2830 & ~n2852 ;
  assign n2854 = n2581 & n2840 ;
  assign n2855 = n2578 & n2837 ;
  assign n2856 = n2854 | n2855 ;
  assign n2857 = ~n2575 & n2832 ;
  assign n2858 = n2856 | n2857 ;
  assign n2859 = n2853 | n2858 ;
  assign n2860 = n903 & ~n2859 ;
  assign n2861 = ~n903 & n2859 ;
  assign n2862 = n2860 | n2861 ;
  assign n2863 = n2850 & n2862 ;
  assign n2864 = n2779 | n2781 ;
  assign n2865 = ~n2782 & n2864 ;
  assign n2866 = n2578 & n2832 ;
  assign n2867 = n2584 & n2840 ;
  assign n2868 = n2581 & n2837 ;
  assign n2869 = n2867 | n2868 ;
  assign n2870 = n2866 | n2869 ;
  assign n2871 = n2609 | n2611 ;
  assign n2872 = ~n2612 & n2871 ;
  assign n2873 = n2830 & n2872 ;
  assign n2874 = n2870 | n2873 ;
  assign n2875 = n903 | n2874 ;
  assign n2876 = n903 & n2874 ;
  assign n2877 = n2875 & ~n2876 ;
  assign n2878 = n2865 & n2877 ;
  assign n2879 = n2752 | n2765 ;
  assign n2880 = ~n2766 & n2879 ;
  assign n2881 = n2805 & n2830 ;
  assign n2882 = n2581 & n2832 ;
  assign n2883 = n2587 & n2840 ;
  assign n2884 = n2584 & n2837 ;
  assign n2885 = n2883 | n2884 ;
  assign n2886 = n2882 | n2885 ;
  assign n2887 = n2881 | n2886 ;
  assign n2888 = n903 & ~n2887 ;
  assign n2889 = ~n903 & n2887 ;
  assign n2890 = n2888 | n2889 ;
  assign n2891 = n2880 & n2890 ;
  assign n2892 = n2743 | n2751 ;
  assign n2893 = ~n2752 & n2892 ;
  assign n2894 = n2722 & n2830 ;
  assign n2895 = ~n2590 & n2840 ;
  assign n2896 = n2587 & n2837 ;
  assign n2897 = n2584 & n2832 ;
  assign n2898 = n2896 | n2897 ;
  assign n2899 = n2895 | n2898 ;
  assign n2900 = n2894 | n2899 ;
  assign n2901 = n903 | n2900 ;
  assign n2902 = n903 & n2900 ;
  assign n2903 = n2901 & ~n2902 ;
  assign n2904 = n2893 & n2903 ;
  assign n2905 = n2893 | n2903 ;
  assign n2906 = ~n2904 & n2905 ;
  assign n2907 = ~n2590 & n2832 ;
  assign n2908 = ~n2760 & n2830 ;
  assign n2909 = n2593 & n2837 ;
  assign n2910 = n2595 & n2840 ;
  assign n2911 = n2909 | n2910 ;
  assign n2912 = n2908 | n2911 ;
  assign n2913 = n2907 | n2912 ;
  assign n2914 = n903 | n2913 ;
  assign n2915 = n903 & n2913 ;
  assign n2916 = n2914 & ~n2915 ;
  assign n2917 = n2595 & n2829 ;
  assign n2918 = n903 & ~n2917 ;
  assign n2919 = n2595 & n2837 ;
  assign n2920 = n2701 & n2830 ;
  assign n2921 = n2593 & n2832 ;
  assign n2922 = n2920 | n2921 ;
  assign n2923 = n2919 | n2922 ;
  assign n2924 = n903 & ~n2923 ;
  assign n2925 = ~n903 & n2923 ;
  assign n2926 = n2924 | n2925 ;
  assign n2927 = n2918 & n2926 ;
  assign n2928 = n2916 & n2927 ;
  assign n2929 = n2742 & n2928 ;
  assign n2930 = ~n2590 & n2837 ;
  assign n2931 = ~n2770 & n2830 ;
  assign n2932 = n2587 & n2832 ;
  assign n2933 = n2593 & n2840 ;
  assign n2934 = n2932 | n2933 ;
  assign n2935 = n2931 | n2934 ;
  assign n2936 = n2930 | n2935 ;
  assign n2937 = n903 & ~n2936 ;
  assign n2938 = ~n903 & n2936 ;
  assign n2939 = n2937 | n2938 ;
  assign n2940 = n2742 | n2928 ;
  assign n2941 = ~n2929 & n2940 ;
  assign n2942 = n2939 & n2941 ;
  assign n2943 = n2929 | n2942 ;
  assign n2944 = n2906 & n2943 ;
  assign n2945 = n2904 | n2944 ;
  assign n2946 = n2880 | n2890 ;
  assign n2947 = ~n2891 & n2946 ;
  assign n2948 = n2945 & n2947 ;
  assign n2949 = n2891 | n2948 ;
  assign n2950 = n2865 | n2877 ;
  assign n2951 = ~n2878 & n2950 ;
  assign n2952 = n2949 & n2951 ;
  assign n2953 = n2878 | n2952 ;
  assign n2954 = n2850 | n2862 ;
  assign n2955 = ~n2863 & n2954 ;
  assign n2956 = n2953 & n2955 ;
  assign n2957 = n2863 | n2956 ;
  assign n2958 = n2821 | n2847 ;
  assign n2959 = ~n2848 & n2958 ;
  assign n2960 = n2957 & n2959 ;
  assign n2961 = n2848 | n2960 ;
  assign n2962 = n2816 | n2820 ;
  assign n2963 = n2578 & n2732 ;
  assign n2964 = n2720 & n2872 ;
  assign n2965 = n2581 & n2730 ;
  assign n2966 = n2584 & n2728 ;
  assign n2967 = n2965 | n2966 ;
  assign n2968 = n2964 | n2967 ;
  assign n2969 = n2963 | n2968 ;
  assign n2970 = n372 & n2969 ;
  assign n2971 = n372 | n2969 ;
  assign n2972 = ~n2970 & n2971 ;
  assign n2973 = n2702 & ~n2770 ;
  assign n2974 = ~n2590 & n2695 ;
  assign n2975 = n2587 & n2697 ;
  assign n2976 = n2593 & n2793 ;
  assign n2977 = n2975 | n2976 ;
  assign n2978 = n2974 | n2977 ;
  assign n2979 = n2973 | n2978 ;
  assign n2980 = n221 & ~n2979 ;
  assign n2981 = ~n221 & n2979 ;
  assign n2982 = n2980 | n2981 ;
  assign n2983 = n221 & n2595 ;
  assign n2984 = n2801 | n2983 ;
  assign n2985 = n2708 & n2983 ;
  assign n2986 = n2800 & n2985 ;
  assign n2987 = ~n2709 & n2986 ;
  assign n2988 = n2984 & ~n2987 ;
  assign n2989 = n2982 & n2988 ;
  assign n2990 = n2982 | n2988 ;
  assign n2991 = ~n2989 & n2990 ;
  assign n2992 = n2972 & n2991 ;
  assign n2993 = n2972 | n2991 ;
  assign n2994 = ~n2992 & n2993 ;
  assign n2995 = n2962 & n2994 ;
  assign n2996 = n2962 | n2994 ;
  assign n2997 = ~n2995 & n2996 ;
  assign n2998 = n2621 | n2623 ;
  assign n2999 = ~n2624 & n2998 ;
  assign n3000 = n2830 & n2999 ;
  assign n3001 = n2569 & n2832 ;
  assign n3002 = n2572 & n2837 ;
  assign n3003 = ~n2575 & n2840 ;
  assign n3004 = n3002 | n3003 ;
  assign n3005 = n3001 | n3004 ;
  assign n3006 = n3000 | n3005 ;
  assign n3007 = n903 | n3006 ;
  assign n3008 = n903 & n3006 ;
  assign n3009 = n3007 & ~n3008 ;
  assign n3010 = n2997 & n3009 ;
  assign n3011 = n2997 | n3009 ;
  assign n3012 = ~n3010 & n3011 ;
  assign n3013 = n2961 & n3012 ;
  assign n3014 = n2848 | n3012 ;
  assign n3015 = n2960 | n3014 ;
  assign n3016 = ~n1199 & n1248 ;
  assign n3017 = n1199 & ~n1248 ;
  assign n3018 = n3016 | n3017 ;
  assign n3019 = n29 & ~n1339 ;
  assign n3020 = ~n29 & n1339 ;
  assign n3021 = n3019 | n3020 ;
  assign n3022 = ~n3018 & n3021 ;
  assign n3023 = n2557 & n3022 ;
  assign n3024 = ~n2631 & n2633 ;
  assign n3025 = n2634 | n3024 ;
  assign n3026 = n3018 & n3021 ;
  assign n3027 = ~n3025 & n3026 ;
  assign n3028 = n1248 & ~n1339 ;
  assign n3029 = ~n1248 & n1339 ;
  assign n3030 = n3028 | n3029 ;
  assign n3031 = n3018 & ~n3021 ;
  assign n3032 = ~n3030 & n3031 ;
  assign n3033 = n2564 & n3032 ;
  assign n3034 = ~n3021 & n3030 ;
  assign n3035 = ~n2561 & n3034 ;
  assign n3036 = n3033 | n3035 ;
  assign n3037 = n3027 | n3036 ;
  assign n3038 = n3023 | n3037 ;
  assign n3039 = n1199 & n3038 ;
  assign n3040 = n1199 | n3038 ;
  assign n3041 = ~n3039 & n3040 ;
  assign n3042 = n3015 & n3041 ;
  assign n3043 = ~n3013 & n3042 ;
  assign n3044 = n2863 | n2959 ;
  assign n3045 = n2956 | n3044 ;
  assign n3046 = ~n2561 & n3022 ;
  assign n3047 = n2569 & n3032 ;
  assign n3048 = n2564 & n3034 ;
  assign n3049 = n3047 | n3048 ;
  assign n3050 = n3046 | n3049 ;
  assign n3051 = n2567 & ~n2629 ;
  assign n3052 = n2630 | n3051 ;
  assign n3053 = n3026 & ~n3052 ;
  assign n3054 = n3050 | n3053 ;
  assign n3055 = n1199 & n3054 ;
  assign n3056 = n1199 | n3054 ;
  assign n3057 = ~n3055 & n3056 ;
  assign n3058 = n3045 & n3057 ;
  assign n3059 = ~n2960 & n3058 ;
  assign n3060 = n2878 | n2955 ;
  assign n3061 = n2952 | n3060 ;
  assign n3062 = n2564 & n3022 ;
  assign n3063 = n2625 | n2627 ;
  assign n3064 = ~n2628 & n3063 ;
  assign n3065 = n3026 & n3064 ;
  assign n3066 = n2572 & n3032 ;
  assign n3067 = n2569 & n3034 ;
  assign n3068 = n3066 | n3067 ;
  assign n3069 = n3065 | n3068 ;
  assign n3070 = n3062 | n3069 ;
  assign n3071 = n1199 | n3070 ;
  assign n3072 = n1199 & n3070 ;
  assign n3073 = n3071 & ~n3072 ;
  assign n3074 = n3061 & n3073 ;
  assign n3075 = ~n2956 & n3074 ;
  assign n3076 = n2891 | n2951 ;
  assign n3077 = n2948 | n3076 ;
  assign n3078 = n2569 & n3022 ;
  assign n3079 = n2999 & n3026 ;
  assign n3080 = ~n2575 & n3032 ;
  assign n3081 = n2572 & n3034 ;
  assign n3082 = n3080 | n3081 ;
  assign n3083 = n3079 | n3082 ;
  assign n3084 = n3078 | n3083 ;
  assign n3085 = n1199 | n3084 ;
  assign n3086 = n1199 & n3084 ;
  assign n3087 = n3085 & ~n3086 ;
  assign n3088 = n3077 & n3087 ;
  assign n3089 = ~n2952 & n3088 ;
  assign n3090 = ~n2952 & n3077 ;
  assign n3091 = n3087 | n3090 ;
  assign n3092 = n2945 | n2947 ;
  assign n3093 = ~n2948 & n3092 ;
  assign n3094 = n2572 & n3022 ;
  assign n3095 = ~n2823 & n3026 ;
  assign n3096 = n2578 & n3032 ;
  assign n3097 = ~n2575 & n3034 ;
  assign n3098 = n3096 | n3097 ;
  assign n3099 = n3095 | n3098 ;
  assign n3100 = n3094 | n3099 ;
  assign n3101 = n1199 | n3100 ;
  assign n3102 = n1199 & n3100 ;
  assign n3103 = n3101 & ~n3102 ;
  assign n3104 = n3093 & n3103 ;
  assign n3105 = n2906 | n2943 ;
  assign n3106 = ~n2944 & n3105 ;
  assign n3107 = ~n2575 & n3022 ;
  assign n3108 = ~n2852 & n3026 ;
  assign n3109 = n2581 & n3032 ;
  assign n3110 = n2578 & n3034 ;
  assign n3111 = n3109 | n3110 ;
  assign n3112 = n3108 | n3111 ;
  assign n3113 = n3107 | n3112 ;
  assign n3114 = n1199 & n3113 ;
  assign n3115 = n1199 | n3113 ;
  assign n3116 = ~n3114 & n3115 ;
  assign n3117 = n3106 & n3116 ;
  assign n3118 = n2939 | n2941 ;
  assign n3119 = ~n2942 & n3118 ;
  assign n3120 = n2578 & n3022 ;
  assign n3121 = n2584 & n3032 ;
  assign n3122 = n2581 & n3034 ;
  assign n3123 = n3121 | n3122 ;
  assign n3124 = n3120 | n3123 ;
  assign n3125 = n2872 & n3026 ;
  assign n3126 = n3124 | n3125 ;
  assign n3127 = n1199 & n3126 ;
  assign n3128 = n1199 | n3126 ;
  assign n3129 = ~n3127 & n3128 ;
  assign n3130 = n3119 & n3129 ;
  assign n3131 = n2581 & n3022 ;
  assign n3132 = n2805 & n3026 ;
  assign n3133 = n2587 & n3032 ;
  assign n3134 = n2584 & n3034 ;
  assign n3135 = n3133 | n3134 ;
  assign n3136 = n3132 | n3135 ;
  assign n3137 = n3131 | n3136 ;
  assign n3138 = n1199 & n3137 ;
  assign n3139 = n1199 | n3137 ;
  assign n3140 = ~n3138 & n3139 ;
  assign n3141 = n2916 | n2927 ;
  assign n3142 = ~n2928 & n3141 ;
  assign n3143 = n3140 & n3142 ;
  assign n3144 = n2722 & n3026 ;
  assign n3145 = ~n2590 & n3032 ;
  assign n3146 = n2587 & n3034 ;
  assign n3147 = n2584 & n3022 ;
  assign n3148 = n3146 | n3147 ;
  assign n3149 = n3145 | n3148 ;
  assign n3150 = n3144 | n3149 ;
  assign n3151 = n1199 | n3150 ;
  assign n3152 = n1199 & n3150 ;
  assign n3153 = n3151 & ~n3152 ;
  assign n3154 = n2918 | n2926 ;
  assign n3155 = ~n2927 & n3154 ;
  assign n3156 = n3153 & n3155 ;
  assign n3157 = n2595 & n3034 ;
  assign n3158 = n2701 & n3026 ;
  assign n3159 = n2593 & n3022 ;
  assign n3160 = n3158 | n3159 ;
  assign n3161 = n3157 | n3160 ;
  assign n3162 = n1199 & n3161 ;
  assign n3163 = ~n2760 & n3026 ;
  assign n3164 = n2593 & n3034 ;
  assign n3165 = n3163 | n3164 ;
  assign n3166 = n2595 & n3032 ;
  assign n3167 = ~n2590 & n3022 ;
  assign n3168 = n1199 | n3167 ;
  assign n3169 = n3166 | n3168 ;
  assign n3170 = n3165 | n3169 ;
  assign n3171 = ~n3162 & n3170 ;
  assign n3172 = n3164 | n3167 ;
  assign n3173 = n3163 | n3172 ;
  assign n3174 = n3166 | n3173 ;
  assign n3175 = n1199 & n3174 ;
  assign n3176 = n1199 | n3157 ;
  assign n3177 = n3160 | n3176 ;
  assign n3178 = n2595 & n3021 ;
  assign n3179 = n1199 & n2917 ;
  assign n3180 = ~n3178 & n3179 ;
  assign n3181 = n3177 & n3180 ;
  assign n3182 = ~n3175 & n3181 ;
  assign n3183 = n3171 & n3182 ;
  assign n3184 = n3170 & ~n3175 ;
  assign n3185 = n1199 & ~n3178 ;
  assign n3186 = n3177 & n3185 ;
  assign n3187 = ~n3162 & n3186 ;
  assign n3188 = n3184 & n3187 ;
  assign n3189 = n2917 | n3188 ;
  assign n3190 = ~n2590 & n3034 ;
  assign n3191 = ~n2770 & n3026 ;
  assign n3192 = n2587 & n3022 ;
  assign n3193 = n2593 & n3032 ;
  assign n3194 = n3192 | n3193 ;
  assign n3195 = n3191 | n3194 ;
  assign n3196 = n3190 | n3195 ;
  assign n3197 = n1199 & n3196 ;
  assign n3198 = n1199 | n3196 ;
  assign n3199 = ~n3197 & n3198 ;
  assign n3200 = ~n3183 & n3199 ;
  assign n3201 = n3189 & n3200 ;
  assign n3202 = n3183 | n3201 ;
  assign n3203 = n3153 | n3155 ;
  assign n3204 = ~n3156 & n3203 ;
  assign n3205 = n3202 & n3204 ;
  assign n3206 = n3156 | n3205 ;
  assign n3207 = n3140 | n3142 ;
  assign n3208 = ~n3143 & n3207 ;
  assign n3209 = n3206 & n3208 ;
  assign n3210 = n3143 | n3209 ;
  assign n3211 = n3119 | n3129 ;
  assign n3212 = ~n3130 & n3211 ;
  assign n3213 = n3210 & n3212 ;
  assign n3214 = n3130 | n3213 ;
  assign n3215 = n3106 | n3116 ;
  assign n3216 = ~n3117 & n3215 ;
  assign n3217 = n3214 & n3216 ;
  assign n3218 = n3117 | n3217 ;
  assign n3219 = n3093 | n3103 ;
  assign n3220 = ~n3104 & n3219 ;
  assign n3221 = n3218 & n3220 ;
  assign n3222 = n3104 | n3221 ;
  assign n3223 = ~n3089 & n3222 ;
  assign n3224 = n3091 & n3223 ;
  assign n3225 = n3089 | n3224 ;
  assign n3226 = ~n2956 & n3061 ;
  assign n3227 = n3073 | n3226 ;
  assign n3228 = ~n3075 & n3227 ;
  assign n3229 = n3225 & n3228 ;
  assign n3230 = n3075 | n3229 ;
  assign n3231 = ~n2960 & n3045 ;
  assign n3232 = n3057 | n3231 ;
  assign n3233 = ~n3059 & n3232 ;
  assign n3234 = n3230 & n3233 ;
  assign n3235 = n3059 | n3234 ;
  assign n3236 = ~n3013 & n3015 ;
  assign n3237 = n3041 | n3236 ;
  assign n3238 = ~n3043 & n3237 ;
  assign n3239 = n3235 & n3238 ;
  assign n3240 = n3043 | n3239 ;
  assign n3241 = n3010 | n3013 ;
  assign n3242 = n2992 | n2995 ;
  assign n3243 = ~n2575 & n2732 ;
  assign n3244 = n2720 & ~n2852 ;
  assign n3245 = n2578 & n2730 ;
  assign n3246 = n2581 & n2728 ;
  assign n3247 = n3245 | n3246 ;
  assign n3248 = n3244 | n3247 ;
  assign n3249 = n3243 | n3248 ;
  assign n3250 = n372 & n3249 ;
  assign n3251 = n372 | n3249 ;
  assign n3252 = ~n3250 & n3251 ;
  assign n3253 = n2987 | n2989 ;
  assign n3254 = n2702 & n2722 ;
  assign n3255 = ~n2590 & n2793 ;
  assign n3256 = n2587 & n2695 ;
  assign n3257 = n2584 & n2697 ;
  assign n3258 = n3256 | n3257 ;
  assign n3259 = n3255 | n3258 ;
  assign n3260 = n3254 | n3259 ;
  assign n3261 = n221 & ~n2593 ;
  assign n3262 = n3260 | n3261 ;
  assign n3263 = n3260 & n3261 ;
  assign n3264 = n3262 & ~n3263 ;
  assign n3265 = n3253 & n3264 ;
  assign n3266 = n3253 | n3264 ;
  assign n3267 = ~n3265 & n3266 ;
  assign n3268 = n3252 & n3267 ;
  assign n3269 = n3252 | n3267 ;
  assign n3270 = ~n3268 & n3269 ;
  assign n3271 = n3242 & n3270 ;
  assign n3272 = n3242 | n3270 ;
  assign n3273 = ~n3271 & n3272 ;
  assign n3274 = n2830 & n3064 ;
  assign n3275 = n2564 & n2832 ;
  assign n3276 = n2569 & n2837 ;
  assign n3277 = n2572 & n2840 ;
  assign n3278 = n3276 | n3277 ;
  assign n3279 = n3275 | n3278 ;
  assign n3280 = n3274 | n3279 ;
  assign n3281 = n903 | n3280 ;
  assign n3282 = n903 & n3280 ;
  assign n3283 = n3281 & ~n3282 ;
  assign n3284 = n3273 & n3283 ;
  assign n3285 = n3273 | n3283 ;
  assign n3286 = ~n3284 & n3285 ;
  assign n3287 = n3241 & n3286 ;
  assign n3288 = n3010 | n3286 ;
  assign n3289 = n3013 | n3288 ;
  assign n3290 = ~n3287 & n3289 ;
  assign n3291 = n2553 & n3022 ;
  assign n3292 = n2635 | n2637 ;
  assign n3293 = ~n2638 & n3292 ;
  assign n3294 = n3026 & n3293 ;
  assign n3295 = ~n2561 & n3032 ;
  assign n3296 = n2557 & n3034 ;
  assign n3297 = n3295 | n3296 ;
  assign n3298 = n3294 | n3297 ;
  assign n3299 = n3291 | n3298 ;
  assign n3300 = n1199 & n3299 ;
  assign n3301 = n1199 | n3299 ;
  assign n3302 = ~n3300 & n3301 ;
  assign n3303 = n3290 | n3302 ;
  assign n3304 = n3289 & n3302 ;
  assign n3305 = ~n3287 & n3304 ;
  assign n3306 = n3303 & ~n3305 ;
  assign n3307 = n3240 & n3306 ;
  assign n3308 = n3240 | n3306 ;
  assign n3309 = ~n3307 & n3308 ;
  assign n3310 = n2688 & n3309 ;
  assign n3311 = n2688 | n3309 ;
  assign n3312 = ~n3310 & n3311 ;
  assign n3313 = ~n2643 & n2645 ;
  assign n3314 = n2646 | n3313 ;
  assign n3315 = n2675 & ~n3314 ;
  assign n3316 = n2547 & n2677 ;
  assign n3317 = n2553 & n2679 ;
  assign n3318 = ~n2549 & n2681 ;
  assign n3319 = n3317 | n3318 ;
  assign n3320 = n3316 | n3319 ;
  assign n3321 = n3315 | n3320 ;
  assign n3322 = n29 | n3321 ;
  assign n3323 = n29 & n3321 ;
  assign n3324 = n3322 & ~n3323 ;
  assign n3325 = n3235 | n3238 ;
  assign n3326 = ~n3239 & n3325 ;
  assign n3327 = n3324 & n3326 ;
  assign n3328 = ~n2639 & n2641 ;
  assign n3329 = n2642 | n3328 ;
  assign n3330 = n2675 & ~n3329 ;
  assign n3331 = ~n2549 & n2677 ;
  assign n3332 = n2557 & n2679 ;
  assign n3333 = n2553 & n2681 ;
  assign n3334 = n3332 | n3333 ;
  assign n3335 = n3331 | n3334 ;
  assign n3336 = n3330 | n3335 ;
  assign n3337 = n29 | n3336 ;
  assign n3338 = n29 & n3336 ;
  assign n3339 = n3337 & ~n3338 ;
  assign n3340 = n3230 | n3233 ;
  assign n3341 = ~n3234 & n3340 ;
  assign n3342 = n3339 & n3341 ;
  assign n3343 = n3339 | n3341 ;
  assign n3344 = ~n3342 & n3343 ;
  assign n3345 = n2675 & n3293 ;
  assign n3346 = n2553 & n2677 ;
  assign n3347 = ~n2561 & n2679 ;
  assign n3348 = n2557 & n2681 ;
  assign n3349 = n3347 | n3348 ;
  assign n3350 = n3346 | n3349 ;
  assign n3351 = n3345 | n3350 ;
  assign n3352 = n29 & ~n3351 ;
  assign n3353 = ~n29 & n3351 ;
  assign n3354 = n3352 | n3353 ;
  assign n3355 = n3218 | n3220 ;
  assign n3356 = ~n3221 & n3355 ;
  assign n3357 = n3130 | n3216 ;
  assign n3358 = n3213 | n3357 ;
  assign n3359 = ~n3217 & n3358 ;
  assign n3360 = n2569 & n2681 ;
  assign n3361 = n2675 & n3064 ;
  assign n3362 = n2564 & n2677 ;
  assign n3363 = n3361 | n3362 ;
  assign n3364 = n2572 & n2679 ;
  assign n3365 = n3363 | n3364 ;
  assign n3366 = n3360 | n3365 ;
  assign n3367 = n29 & ~n3366 ;
  assign n3368 = ~n29 & n3366 ;
  assign n3369 = n3367 | n3368 ;
  assign n3370 = n3359 | n3369 ;
  assign n3371 = n3210 | n3212 ;
  assign n3372 = ~n3213 & n3371 ;
  assign n3373 = ~n2575 & n2679 ;
  assign n3374 = n2572 & n2681 ;
  assign n3375 = n3373 | n3374 ;
  assign n3376 = n2675 & n2999 ;
  assign n3377 = n2569 & n2677 ;
  assign n3378 = n3376 | n3377 ;
  assign n3379 = n3375 | n3378 ;
  assign n3380 = n29 & ~n3379 ;
  assign n3381 = ~n29 & n3379 ;
  assign n3382 = n3380 | n3381 ;
  assign n3383 = n3372 & n3382 ;
  assign n3384 = n3358 & n3369 ;
  assign n3385 = ~n3217 & n3384 ;
  assign n3386 = n3383 | n3385 ;
  assign n3387 = n3206 | n3208 ;
  assign n3388 = ~n3209 & n3387 ;
  assign n3389 = n2578 & n2679 ;
  assign n3390 = ~n2575 & n2681 ;
  assign n3391 = n3389 | n3390 ;
  assign n3392 = n2675 & ~n2823 ;
  assign n3393 = n2572 & n2677 ;
  assign n3394 = n3392 | n3393 ;
  assign n3395 = n3391 | n3394 ;
  assign n3396 = n29 & ~n3395 ;
  assign n3397 = ~n29 & n3395 ;
  assign n3398 = n3396 | n3397 ;
  assign n3399 = n3388 & n3398 ;
  assign n3400 = n2578 & n2681 ;
  assign n3401 = n2675 & ~n2852 ;
  assign n3402 = ~n2575 & n2677 ;
  assign n3403 = n3401 | n3402 ;
  assign n3404 = n2581 & n2679 ;
  assign n3405 = n3403 | n3404 ;
  assign n3406 = n3400 | n3405 ;
  assign n3407 = n29 & ~n3406 ;
  assign n3408 = ~n29 & n3406 ;
  assign n3409 = n3407 | n3408 ;
  assign n3410 = ~n3183 & n3189 ;
  assign n3411 = n3199 | n3410 ;
  assign n3412 = ~n3201 & n3411 ;
  assign n3413 = n2578 & n2677 ;
  assign n3414 = n2584 & n2679 ;
  assign n3415 = n2581 & n2681 ;
  assign n3416 = n3414 | n3415 ;
  assign n3417 = n2675 & n2872 ;
  assign n3418 = n3416 | n3417 ;
  assign n3419 = n3413 | n3418 ;
  assign n3420 = n29 & ~n3419 ;
  assign n3421 = ~n29 & n3419 ;
  assign n3422 = n3420 | n3421 ;
  assign n3423 = n3412 | n3422 ;
  assign n3424 = n2675 & n2805 ;
  assign n3425 = n2581 & n2677 ;
  assign n3426 = n2587 & n2679 ;
  assign n3427 = n2584 & n2681 ;
  assign n3428 = n3426 | n3427 ;
  assign n3429 = n3425 | n3428 ;
  assign n3430 = n3424 | n3429 ;
  assign n3431 = n29 & ~n3430 ;
  assign n3432 = ~n29 & n3430 ;
  assign n3433 = n3431 | n3432 ;
  assign n3434 = n3184 | n3187 ;
  assign n3435 = ~n3188 & n3434 ;
  assign n3436 = n3433 & n3435 ;
  assign n3437 = ~n3162 & n3177 ;
  assign n3438 = n3185 | n3437 ;
  assign n3439 = ~n3187 & n3438 ;
  assign n3440 = n2584 & n2677 ;
  assign n3441 = n2675 & n2722 ;
  assign n3442 = ~n2590 & n2679 ;
  assign n3443 = n3441 | n3442 ;
  assign n3444 = n2587 & n2681 ;
  assign n3445 = n3443 | n3444 ;
  assign n3446 = n3440 | n3445 ;
  assign n3447 = n29 & ~n3446 ;
  assign n3448 = ~n29 & n3446 ;
  assign n3449 = n3447 | n3448 ;
  assign n3450 = n3439 | n3449 ;
  assign n3451 = n3433 | n3435 ;
  assign n3452 = n3450 & n3451 ;
  assign n3453 = n3439 & n3449 ;
  assign n3454 = n2593 & n2677 ;
  assign n3455 = ~n2701 & n2760 ;
  assign n3456 = n2675 & ~n3455 ;
  assign n3457 = n3454 | n3456 ;
  assign n3458 = ~n2590 & n2677 ;
  assign n3459 = n2595 & n2679 ;
  assign n3460 = n2593 & n2681 ;
  assign n3461 = n3459 | n3460 ;
  assign n3462 = n3458 | n3461 ;
  assign n3463 = pi0 | n2671 ;
  assign n3464 = n2595 & n3463 ;
  assign n3465 = n29 & ~n3464 ;
  assign n3466 = ~n3462 & n3465 ;
  assign n3467 = ~n3457 & n3466 ;
  assign n3468 = n3178 & n3467 ;
  assign n3469 = n3178 | n3467 ;
  assign n3470 = n2675 & ~n2770 ;
  assign n3471 = ~n2590 & n2681 ;
  assign n3472 = n2587 & n2677 ;
  assign n3473 = n2593 & n2679 ;
  assign n3474 = n3472 | n3473 ;
  assign n3475 = n3471 | n3474 ;
  assign n3476 = n3470 | n3475 ;
  assign n3477 = n29 & ~n3476 ;
  assign n3478 = ~n29 & n3476 ;
  assign n3479 = n3477 | n3478 ;
  assign n3480 = n3469 & n3479 ;
  assign n3481 = n3468 | n3480 ;
  assign n3482 = n3453 | n3481 ;
  assign n3483 = n3452 & n3482 ;
  assign n3484 = ~n3201 & n3422 ;
  assign n3485 = n3411 & n3484 ;
  assign n3486 = n3483 | n3485 ;
  assign n3487 = n3436 | n3486 ;
  assign n3488 = n3423 & n3487 ;
  assign n3489 = n3409 & n3488 ;
  assign n3490 = n3399 | n3489 ;
  assign n3491 = n3409 | n3488 ;
  assign n3492 = n3202 | n3204 ;
  assign n3493 = ~n3205 & n3492 ;
  assign n3494 = n3491 & n3493 ;
  assign n3495 = n3490 | n3494 ;
  assign n3496 = n3372 | n3382 ;
  assign n3497 = n3388 | n3398 ;
  assign n3498 = n3496 & n3497 ;
  assign n3499 = n3495 & n3498 ;
  assign n3500 = n3386 | n3499 ;
  assign n3501 = n3370 & n3500 ;
  assign n3502 = n3356 | n3501 ;
  assign n3503 = n3356 & n3501 ;
  assign n3504 = n2564 & n2681 ;
  assign n3505 = n2675 & ~n3052 ;
  assign n3506 = n3504 | n3505 ;
  assign n3507 = n2569 & n2679 ;
  assign n3508 = ~n2561 & n2677 ;
  assign n3509 = n3507 | n3508 ;
  assign n3510 = n3506 | n3509 ;
  assign n3511 = n29 & ~n3510 ;
  assign n3512 = ~n29 & n3510 ;
  assign n3513 = n3511 | n3512 ;
  assign n3514 = n3503 | n3513 ;
  assign n3515 = n3502 & n3514 ;
  assign n3516 = n2675 & ~n3025 ;
  assign n3517 = n2557 & n2677 ;
  assign n3518 = n2564 & n2679 ;
  assign n3519 = ~n2561 & n2681 ;
  assign n3520 = n3518 | n3519 ;
  assign n3521 = n3517 | n3520 ;
  assign n3522 = n3516 | n3521 ;
  assign n3523 = n29 & ~n3522 ;
  assign n3524 = ~n29 & n3522 ;
  assign n3525 = n3523 | n3524 ;
  assign n3526 = n3515 & n3525 ;
  assign n3527 = n3515 | n3525 ;
  assign n3528 = ~n3089 & n3091 ;
  assign n3529 = n3222 | n3528 ;
  assign n3530 = ~n3224 & n3529 ;
  assign n3531 = n3527 & n3530 ;
  assign n3532 = n3526 | n3531 ;
  assign n3533 = n3354 & n3532 ;
  assign n3534 = n3225 | n3228 ;
  assign n3535 = n3354 | n3532 ;
  assign n3536 = ~n3229 & n3535 ;
  assign n3537 = n3534 & n3536 ;
  assign n3538 = n3533 | n3537 ;
  assign n3539 = n3344 & n3538 ;
  assign n3540 = n3342 | n3539 ;
  assign n3541 = n3324 | n3326 ;
  assign n3542 = ~n3327 & n3541 ;
  assign n3543 = n3540 & n3542 ;
  assign n3544 = n3327 | n3543 ;
  assign n3545 = n3312 & n3544 ;
  assign n3546 = n3312 | n3544 ;
  assign n3547 = ~n3545 & n3546 ;
  assign n3548 = n317 | n339 ;
  assign n3549 = n197 | n2492 ;
  assign n3550 = n474 | n3549 ;
  assign n3551 = n174 | n188 ;
  assign n3552 = n244 | n3551 ;
  assign n3553 = n430 | n3552 ;
  assign n3554 = n268 | n3553 ;
  assign n3555 = n150 | n509 ;
  assign n3556 = n187 | n3555 ;
  assign n3557 = n3554 | n3556 ;
  assign n3558 = n271 | n3557 ;
  assign n3559 = n441 | n3558 ;
  assign n3560 = n3550 | n3559 ;
  assign n3561 = n137 | n245 ;
  assign n3562 = n121 | n3561 ;
  assign n3563 = n154 | n333 ;
  assign n3564 = n500 | n510 ;
  assign n3565 = n167 | n2133 ;
  assign n3566 = n176 | n278 ;
  assign n3567 = n139 | n183 ;
  assign n3568 = n191 | n3567 ;
  assign n3569 = n3566 | n3568 ;
  assign n3570 = n224 | n3569 ;
  assign n3571 = n201 | n3570 ;
  assign n3572 = n3565 | n3571 ;
  assign n3573 = n3564 | n3572 ;
  assign n3574 = n3563 | n3573 ;
  assign n3575 = n3562 | n3574 ;
  assign n3576 = n389 | n3575 ;
  assign n3577 = n281 | n301 ;
  assign n3578 = n164 | n3577 ;
  assign n3579 = n3576 | n3578 ;
  assign n3580 = n379 | n3579 ;
  assign n3581 = n103 | n3580 ;
  assign n3582 = n2027 | n3581 ;
  assign n3583 = n3560 | n3582 ;
  assign n3584 = n3548 | n3583 ;
  assign n3585 = n142 | n161 ;
  assign n3586 = n252 | n3585 ;
  assign n3587 = n3584 | n3586 ;
  assign n3588 = n266 | n3587 ;
  assign n3589 = n3547 & n3588 ;
  assign n3590 = n3547 | n3588 ;
  assign n3591 = ~n3589 & n3590 ;
  assign n3592 = n248 | n279 ;
  assign n3593 = n235 | n3592 ;
  assign n3594 = n155 | n611 ;
  assign n3595 = n236 | n260 ;
  assign n3596 = n334 | n389 ;
  assign n3597 = n293 | n1033 ;
  assign n3598 = n3596 | n3597 ;
  assign n3599 = n3595 | n3598 ;
  assign n3600 = n245 | n314 ;
  assign n3601 = n229 | n231 ;
  assign n3602 = n3600 | n3601 ;
  assign n3603 = n132 | n142 ;
  assign n3604 = n396 | n496 ;
  assign n3605 = n3603 | n3604 ;
  assign n3606 = n3602 | n3605 ;
  assign n3607 = n3599 | n3606 ;
  assign n3608 = n325 | n3607 ;
  assign n3609 = n3594 | n3608 ;
  assign n3610 = n176 | n318 ;
  assign n3611 = n3609 | n3610 ;
  assign n3612 = n145 | n167 ;
  assign n3613 = n106 | n3612 ;
  assign n3614 = n3611 | n3613 ;
  assign n3615 = n206 | n302 ;
  assign n3616 = n205 | n614 ;
  assign n3617 = n328 | n339 ;
  assign n3618 = n400 | n585 ;
  assign n3619 = n3617 | n3618 ;
  assign n3620 = n143 | n148 ;
  assign n3621 = n3619 | n3620 ;
  assign n3622 = n3616 | n3621 ;
  assign n3623 = n252 | n3622 ;
  assign n3624 = n290 | n3623 ;
  assign n3625 = n3615 | n3624 ;
  assign n3626 = n177 | n198 ;
  assign n3627 = n270 | n2158 ;
  assign n3628 = n3626 | n3627 ;
  assign n3629 = n202 | n311 ;
  assign n3630 = n1047 | n3629 ;
  assign n3631 = n272 | n3630 ;
  assign n3632 = n3628 | n3631 ;
  assign n3633 = n3625 | n3632 ;
  assign n3634 = n3614 | n3633 ;
  assign n3635 = n3593 | n3634 ;
  assign n3636 = n3540 | n3542 ;
  assign n3637 = ~n3543 & n3636 ;
  assign n3638 = n3635 & n3637 ;
  assign n3639 = n3344 | n3538 ;
  assign n3640 = ~n3539 & n3639 ;
  assign n3641 = n134 | n143 ;
  assign n3642 = n402 | n3641 ;
  assign n3643 = n137 | n192 ;
  assign n3644 = n173 | n2054 ;
  assign n3645 = n106 | n3644 ;
  assign n3646 = n622 | n3645 ;
  assign n3647 = n295 | n3646 ;
  assign n3648 = n2278 | n3647 ;
  assign n3649 = n240 | n340 ;
  assign n3650 = n249 | n3649 ;
  assign n3651 = n199 | n2207 ;
  assign n3652 = n160 | n3651 ;
  assign n3653 = n2174 | n3652 ;
  assign n3654 = n3650 | n3653 ;
  assign n3655 = n2296 | n2351 ;
  assign n3656 = n419 | n3655 ;
  assign n3657 = n3654 | n3656 ;
  assign n3658 = n3648 | n3657 ;
  assign n3659 = n3643 | n3658 ;
  assign n3660 = n3642 | n3659 ;
  assign n3661 = n154 | n3660 ;
  assign n3662 = n331 | n3661 ;
  assign n3663 = n3635 | n3637 ;
  assign n3664 = n3662 & n3663 ;
  assign n3665 = n3640 & n3664 ;
  assign n3666 = n3638 | n3665 ;
  assign n3667 = n3591 & n3666 ;
  assign n3668 = n3591 | n3666 ;
  assign n3669 = ~n3667 & n3668 ;
  assign n3670 = n3589 | n3667 ;
  assign n3671 = n3310 | n3545 ;
  assign n3672 = n197 | n231 ;
  assign n3673 = n189 | n481 ;
  assign n3674 = n3672 | n3673 ;
  assign n3675 = n161 | n202 ;
  assign n3676 = n227 | n3564 ;
  assign n3677 = n3675 | n3676 ;
  assign n3678 = n3674 | n3677 ;
  assign n3679 = n668 | n3678 ;
  assign n3680 = n265 | n457 ;
  assign n3681 = n183 | n3680 ;
  assign n3682 = n2050 | n3681 ;
  assign n3683 = n1068 | n3682 ;
  assign n3684 = n3679 | n3683 ;
  assign n3685 = n167 | n1344 ;
  assign n3686 = n1065 & ~n2159 ;
  assign n3687 = ~n154 & n3686 ;
  assign n3688 = ~n3685 & n3687 ;
  assign n3689 = ~n3684 & n3688 ;
  assign n3690 = ~n224 & n3689 ;
  assign n3691 = ~n444 & n3690 ;
  assign n3692 = n2660 & n3691 ;
  assign n3693 = n2660 | n3691 ;
  assign n3694 = ~n3692 & n3693 ;
  assign n3695 = ~n2661 & n3694 ;
  assign n3696 = n2661 & ~n3694 ;
  assign n3697 = n3695 | n3696 ;
  assign n3698 = n2663 | n2665 ;
  assign n3699 = ~n3697 & n3698 ;
  assign n3700 = n3697 & ~n3698 ;
  assign n3701 = n3699 | n3700 ;
  assign n3702 = n2675 & ~n3701 ;
  assign n3703 = n2677 & ~n3694 ;
  assign n3704 = n2547 & n2679 ;
  assign n3705 = n2661 & n2681 ;
  assign n3706 = n3704 | n3705 ;
  assign n3707 = n3703 | n3706 ;
  assign n3708 = n3702 | n3707 ;
  assign n3709 = n29 & ~n3708 ;
  assign n3710 = ~n29 & n3708 ;
  assign n3711 = n3709 | n3710 ;
  assign n3712 = n3305 | n3307 ;
  assign n3713 = n3284 | n3287 ;
  assign n3714 = n2572 & n2732 ;
  assign n3715 = n2720 & ~n2823 ;
  assign n3716 = ~n2575 & n2730 ;
  assign n3717 = n2578 & n2728 ;
  assign n3718 = n3716 | n3717 ;
  assign n3719 = n3715 | n3718 ;
  assign n3720 = n3714 | n3719 ;
  assign n3721 = n372 | n3720 ;
  assign n3722 = n372 & n3720 ;
  assign n3723 = n3721 & ~n3722 ;
  assign n3724 = n221 & n2590 ;
  assign n3725 = n2702 & n2805 ;
  assign n3726 = n2581 & n2697 ;
  assign n3727 = n2584 & n2695 ;
  assign n3728 = n2587 & n2793 ;
  assign n3729 = n3727 | n3728 ;
  assign n3730 = n3726 | n3729 ;
  assign n3731 = n3725 | n3730 ;
  assign n3732 = n3724 & n3731 ;
  assign n3733 = n3724 | n3731 ;
  assign n3734 = ~n3732 & n3733 ;
  assign n3735 = n221 & ~n3260 ;
  assign n3736 = n2593 & n3735 ;
  assign n3737 = n3265 | n3736 ;
  assign n3738 = n3734 & n3737 ;
  assign n3739 = n3734 | n3737 ;
  assign n3740 = ~n3738 & n3739 ;
  assign n3741 = n3723 & n3740 ;
  assign n3742 = n3723 | n3740 ;
  assign n3743 = ~n3741 & n3742 ;
  assign n3744 = n3268 | n3271 ;
  assign n3745 = n3743 & n3744 ;
  assign n3746 = n3743 | n3744 ;
  assign n3747 = ~n3745 & n3746 ;
  assign n3748 = n2830 & ~n3052 ;
  assign n3749 = ~n2561 & n2832 ;
  assign n3750 = n2564 & n2837 ;
  assign n3751 = n2569 & n2840 ;
  assign n3752 = n3750 | n3751 ;
  assign n3753 = n3749 | n3752 ;
  assign n3754 = n3748 | n3753 ;
  assign n3755 = n903 & ~n3754 ;
  assign n3756 = ~n903 & n3754 ;
  assign n3757 = n3755 | n3756 ;
  assign n3758 = n3747 & n3757 ;
  assign n3759 = n3747 | n3757 ;
  assign n3760 = ~n3758 & n3759 ;
  assign n3761 = n3713 & n3760 ;
  assign n3762 = n3284 | n3760 ;
  assign n3763 = n3287 | n3762 ;
  assign n3764 = ~n3761 & n3763 ;
  assign n3765 = ~n2549 & n3022 ;
  assign n3766 = n3026 & ~n3329 ;
  assign n3767 = n2557 & n3032 ;
  assign n3768 = n2553 & n3034 ;
  assign n3769 = n3767 | n3768 ;
  assign n3770 = n3766 | n3769 ;
  assign n3771 = n3765 | n3770 ;
  assign n3772 = n1199 | n3771 ;
  assign n3773 = n1199 & n3771 ;
  assign n3774 = n3772 & ~n3773 ;
  assign n3775 = n3764 | n3774 ;
  assign n3776 = n3763 & n3774 ;
  assign n3777 = ~n3761 & n3776 ;
  assign n3778 = n3775 & ~n3777 ;
  assign n3779 = n3712 & n3778 ;
  assign n3780 = n3712 | n3778 ;
  assign n3781 = ~n3779 & n3780 ;
  assign n3782 = n3711 & n3781 ;
  assign n3783 = n3711 | n3781 ;
  assign n3784 = ~n3782 & n3783 ;
  assign n3785 = n3671 & n3784 ;
  assign n3786 = n3310 | n3784 ;
  assign n3787 = n3545 | n3786 ;
  assign n3788 = ~n3785 & n3787 ;
  assign n3789 = n614 | n1347 ;
  assign n3790 = n971 | n3564 ;
  assign n3791 = n3789 | n3790 ;
  assign n3792 = n2221 | n3791 ;
  assign n3793 = n3549 | n3792 ;
  assign n3794 = n415 | n3793 ;
  assign n3795 = n436 | n3794 ;
  assign n3796 = n132 | n650 ;
  assign n3797 = n309 | n3796 ;
  assign n3798 = n3795 | n3797 ;
  assign n3799 = n3788 | n3798 ;
  assign n3800 = n3787 & n3798 ;
  assign n3801 = ~n3785 & n3800 ;
  assign n3802 = n3799 & ~n3801 ;
  assign n3803 = n3670 & n3802 ;
  assign n3804 = n3670 | n3802 ;
  assign n3805 = ~n3803 & n3804 ;
  assign n3806 = n3669 & n3805 ;
  assign n3807 = n3669 | n3805 ;
  assign n3808 = ~n3806 & n3807 ;
  assign n3809 = pi22 & ~pi23 ;
  assign n3810 = ~pi22 & pi23 ;
  assign n3811 = n3809 | n3810 ;
  assign n3812 = n3808 & n3811 ;
  assign n3813 = n3801 | n3803 ;
  assign n3814 = n3782 | n3785 ;
  assign n3815 = n3696 | n3699 ;
  assign n3816 = n226 | n271 ;
  assign n3817 = n2082 | n2133 ;
  assign n3818 = n286 | n338 ;
  assign n3819 = n2351 | n3818 ;
  assign n3820 = n3817 | n3819 ;
  assign n3821 = n317 | n3820 ;
  assign n3822 = n3816 | n3821 ;
  assign n3823 = n501 | n801 ;
  assign n3824 = n624 | n3823 ;
  assign n3825 = n1364 & ~n3824 ;
  assign n3826 = ~n3822 & n3825 ;
  assign n3827 = n855 | n2350 ;
  assign n3828 = n3826 & ~n3827 ;
  assign n3829 = ~n314 & n3828 ;
  assign n3830 = n235 | n398 ;
  assign n3831 = n260 | n3830 ;
  assign n3832 = n3829 & ~n3831 ;
  assign n3833 = n3692 | n3832 ;
  assign n3834 = n3692 & n3832 ;
  assign n3835 = n3833 & ~n3834 ;
  assign n3836 = n3694 | n3835 ;
  assign n3837 = n3694 & n3835 ;
  assign n3838 = n3836 & ~n3837 ;
  assign n3839 = n3815 & n3838 ;
  assign n3840 = n3696 | n3838 ;
  assign n3841 = n3699 | n3840 ;
  assign n3842 = ~n3839 & n3841 ;
  assign n3843 = n2675 & n3842 ;
  assign n3844 = n2677 & ~n3835 ;
  assign n3845 = n2661 & n2679 ;
  assign n3846 = n2681 & ~n3694 ;
  assign n3847 = n3845 | n3846 ;
  assign n3848 = n3844 | n3847 ;
  assign n3849 = n3843 | n3848 ;
  assign n3850 = n29 & ~n3849 ;
  assign n3851 = ~n29 & n3849 ;
  assign n3852 = n3850 | n3851 ;
  assign n3853 = n3777 | n3779 ;
  assign n3854 = n3758 | n3761 ;
  assign n3855 = n3741 | n3745 ;
  assign n3856 = n2569 & n2732 ;
  assign n3857 = n2720 & n2999 ;
  assign n3858 = n2572 & n2730 ;
  assign n3859 = ~n2575 & n2728 ;
  assign n3860 = n3858 | n3859 ;
  assign n3861 = n3857 | n3860 ;
  assign n3862 = n3856 | n3861 ;
  assign n3863 = n372 | n3862 ;
  assign n3864 = n372 & n3862 ;
  assign n3865 = n3863 & ~n3864 ;
  assign n3866 = n2702 & n2872 ;
  assign n3867 = n2578 & n2697 ;
  assign n3868 = n2581 & n2695 ;
  assign n3869 = n2584 & n2793 ;
  assign n3870 = n3868 | n3869 ;
  assign n3871 = n3867 | n3870 ;
  assign n3872 = n3866 | n3871 ;
  assign n3873 = n221 & ~n2587 ;
  assign n3874 = n3872 & n3873 ;
  assign n3875 = n3872 | n3873 ;
  assign n3876 = ~n3874 & n3875 ;
  assign n3877 = n221 & ~n3731 ;
  assign n3878 = ~n2590 & n3877 ;
  assign n3879 = n3738 | n3878 ;
  assign n3880 = n3876 & n3879 ;
  assign n3881 = n3876 | n3879 ;
  assign n3882 = ~n3880 & n3881 ;
  assign n3883 = n3865 & n3882 ;
  assign n3884 = n3865 | n3882 ;
  assign n3885 = ~n3883 & n3884 ;
  assign n3886 = n3855 & n3885 ;
  assign n3887 = n3855 | n3885 ;
  assign n3888 = ~n3886 & n3887 ;
  assign n3889 = n2830 & ~n3025 ;
  assign n3890 = n2557 & n2832 ;
  assign n3891 = n2564 & n2840 ;
  assign n3892 = ~n2561 & n2837 ;
  assign n3893 = n3891 | n3892 ;
  assign n3894 = n3890 | n3893 ;
  assign n3895 = n3889 | n3894 ;
  assign n3896 = n903 & ~n3895 ;
  assign n3897 = ~n903 & n3895 ;
  assign n3898 = n3896 | n3897 ;
  assign n3899 = n3888 & n3898 ;
  assign n3900 = n3888 | n3898 ;
  assign n3901 = ~n3899 & n3900 ;
  assign n3902 = n3854 & n3901 ;
  assign n3903 = n3758 | n3901 ;
  assign n3904 = n3761 | n3903 ;
  assign n3905 = ~n3902 & n3904 ;
  assign n3906 = n2547 & n3022 ;
  assign n3907 = n3026 & ~n3314 ;
  assign n3908 = n2553 & n3032 ;
  assign n3909 = ~n2549 & n3034 ;
  assign n3910 = n3908 | n3909 ;
  assign n3911 = n3907 | n3910 ;
  assign n3912 = n3906 | n3911 ;
  assign n3913 = n1199 | n3912 ;
  assign n3914 = n1199 & n3912 ;
  assign n3915 = n3913 & ~n3914 ;
  assign n3916 = n3905 | n3915 ;
  assign n3917 = n3904 & n3915 ;
  assign n3918 = ~n3902 & n3917 ;
  assign n3919 = n3916 & ~n3918 ;
  assign n3920 = n3853 & n3919 ;
  assign n3921 = n3853 | n3919 ;
  assign n3922 = ~n3920 & n3921 ;
  assign n3923 = n3852 & n3922 ;
  assign n3924 = n3852 | n3922 ;
  assign n3925 = ~n3923 & n3924 ;
  assign n3926 = n3814 & n3925 ;
  assign n3927 = n3782 | n3925 ;
  assign n3928 = n3785 | n3927 ;
  assign n3929 = ~n3926 & n3928 ;
  assign n3930 = n2183 | n2241 ;
  assign n3931 = n431 | n3930 ;
  assign n3932 = n2082 | n3931 ;
  assign n3933 = n118 | n206 ;
  assign n3934 = n1345 | n3933 ;
  assign n3935 = n3932 | n3934 ;
  assign n3936 = n2479 | n3549 ;
  assign n3937 = n3576 | n3936 ;
  assign n3938 = n3935 | n3937 ;
  assign n3939 = n182 | n3938 ;
  assign n3940 = n173 | n3939 ;
  assign n3941 = n198 | n3940 ;
  assign n3942 = n231 | n317 ;
  assign n3943 = n244 | n3942 ;
  assign n3944 = n3941 | n3943 ;
  assign n3945 = n3929 | n3944 ;
  assign n3946 = n3928 & n3944 ;
  assign n3947 = ~n3926 & n3946 ;
  assign n3948 = n3945 & ~n3947 ;
  assign n3949 = n3813 & n3948 ;
  assign n3950 = n3813 | n3948 ;
  assign n3951 = ~n3949 & n3950 ;
  assign n3952 = n3806 & n3951 ;
  assign n3953 = n3806 | n3951 ;
  assign n3954 = ~n3952 & n3953 ;
  assign n3955 = n3812 & ~n3954 ;
  assign n3956 = ~n3812 & n3954 ;
  assign n3957 = n3955 | n3956 ;
  assign n3958 = n3808 | n3954 ;
  assign n3959 = n3811 & n3958 ;
  assign n3960 = n3947 | n3949 ;
  assign n3961 = n270 | n328 ;
  assign n3962 = n135 | n603 ;
  assign n3963 = n3654 | n3962 ;
  assign n3964 = n126 | n191 ;
  assign n3965 = n103 | n3964 ;
  assign n3966 = n282 | n444 ;
  assign n3967 = n2042 | n3966 ;
  assign n3968 = n3965 | n3967 ;
  assign n3969 = n421 | n3968 ;
  assign n3970 = n3963 | n3969 ;
  assign n3971 = n202 | n3970 ;
  assign n3972 = n288 | n3971 ;
  assign n3973 = n325 | n398 ;
  assign n3974 = n3972 | n3973 ;
  assign n3975 = n332 | n3974 ;
  assign n3976 = n3961 | n3975 ;
  assign n3977 = n3923 | n3926 ;
  assign n3978 = n2679 & ~n3694 ;
  assign n3979 = n2681 & ~n3835 ;
  assign n3980 = n3694 & ~n3699 ;
  assign n3981 = n3835 | n3980 ;
  assign n3982 = n3835 & ~n3839 ;
  assign n3983 = n3981 & ~n3982 ;
  assign n3984 = n2675 & n3983 ;
  assign n3985 = n3979 | n3984 ;
  assign n3986 = n3978 | n3985 ;
  assign n3987 = n29 & ~n3986 ;
  assign n3988 = ~n29 & n3986 ;
  assign n3989 = n3987 | n3988 ;
  assign n3990 = n3918 | n3920 ;
  assign n3991 = n3899 | n3902 ;
  assign n3992 = n3883 | n3886 ;
  assign n3993 = n2564 & n2732 ;
  assign n3994 = n2720 & n3064 ;
  assign n3995 = n2569 & n2730 ;
  assign n3996 = n2572 & n2728 ;
  assign n3997 = n3995 | n3996 ;
  assign n3998 = n3994 | n3997 ;
  assign n3999 = n3993 | n3998 ;
  assign n4000 = n372 | n3999 ;
  assign n4001 = n372 & n3999 ;
  assign n4002 = n4000 & ~n4001 ;
  assign n4003 = n2702 & ~n2852 ;
  assign n4004 = ~n2575 & n2697 ;
  assign n4005 = n2578 & n2695 ;
  assign n4006 = n2581 & n2793 ;
  assign n4007 = n4005 | n4006 ;
  assign n4008 = n4004 | n4007 ;
  assign n4009 = n4003 | n4008 ;
  assign n4010 = n221 & ~n2584 ;
  assign n4011 = n4009 & n4010 ;
  assign n4012 = n4009 | n4010 ;
  assign n4013 = ~n4011 & n4012 ;
  assign n4014 = n221 & ~n3872 ;
  assign n4015 = n2587 & n4014 ;
  assign n4016 = n3880 | n4015 ;
  assign n4017 = n4013 & n4016 ;
  assign n4018 = n4013 | n4016 ;
  assign n4019 = ~n4017 & n4018 ;
  assign n4020 = n4002 & n4019 ;
  assign n4021 = n4002 | n4019 ;
  assign n4022 = ~n4020 & n4021 ;
  assign n4023 = n3992 & n4022 ;
  assign n4024 = n3992 | n4022 ;
  assign n4025 = ~n4023 & n4024 ;
  assign n4026 = n2830 & n3293 ;
  assign n4027 = n2553 & n2832 ;
  assign n4028 = ~n2561 & n2840 ;
  assign n4029 = n2557 & n2837 ;
  assign n4030 = n4028 | n4029 ;
  assign n4031 = n4027 | n4030 ;
  assign n4032 = n4026 | n4031 ;
  assign n4033 = n903 & ~n4032 ;
  assign n4034 = ~n903 & n4032 ;
  assign n4035 = n4033 | n4034 ;
  assign n4036 = n4025 & n4035 ;
  assign n4037 = n4025 | n4035 ;
  assign n4038 = ~n4036 & n4037 ;
  assign n4039 = n3991 & n4038 ;
  assign n4040 = n3899 | n4038 ;
  assign n4041 = n3902 | n4040 ;
  assign n4042 = ~n4039 & n4041 ;
  assign n4043 = n2661 & n3022 ;
  assign n4044 = n2667 & n3026 ;
  assign n4045 = ~n2549 & n3032 ;
  assign n4046 = n2547 & n3034 ;
  assign n4047 = n4045 | n4046 ;
  assign n4048 = n4044 | n4047 ;
  assign n4049 = n4043 | n4048 ;
  assign n4050 = n1199 | n4049 ;
  assign n4051 = n1199 & n4049 ;
  assign n4052 = n4050 & ~n4051 ;
  assign n4053 = n4042 | n4052 ;
  assign n4054 = n4041 & n4052 ;
  assign n4055 = ~n4039 & n4054 ;
  assign n4056 = n4053 & ~n4055 ;
  assign n4057 = n3990 & n4056 ;
  assign n4058 = n3990 | n4056 ;
  assign n4059 = ~n4057 & n4058 ;
  assign n4060 = n3989 & n4059 ;
  assign n4061 = n3989 | n4059 ;
  assign n4062 = ~n4060 & n4061 ;
  assign n4063 = n3977 & n4062 ;
  assign n4064 = n3977 | n4062 ;
  assign n4065 = ~n4063 & n4064 ;
  assign n4066 = n3976 | n4065 ;
  assign n4067 = n3976 & n4065 ;
  assign n4068 = n4066 & ~n4067 ;
  assign n4069 = n3960 & n4068 ;
  assign n4070 = n3960 | n4068 ;
  assign n4071 = ~n4069 & n4070 ;
  assign n4072 = n3952 & n4071 ;
  assign n4073 = n3952 | n4071 ;
  assign n4074 = ~n4072 & n4073 ;
  assign n4075 = n3959 & ~n4074 ;
  assign n4076 = ~n3959 & n4074 ;
  assign n4077 = n4075 | n4076 ;
  assign n4078 = n3958 | n4074 ;
  assign n4079 = n3811 & n4078 ;
  assign n4080 = n4067 | n4069 ;
  assign n4081 = n182 | n293 ;
  assign n4082 = n2241 | n3619 ;
  assign n4083 = n827 | n4082 ;
  assign n4084 = n657 | n1356 ;
  assign n4085 = n4083 | n4084 ;
  assign n4086 = n459 | n2103 ;
  assign n4087 = n199 | n4086 ;
  assign n4088 = n4085 | n4087 ;
  assign n4089 = n4081 | n4088 ;
  assign n4090 = n402 | n4089 ;
  assign n4091 = n266 | n4090 ;
  assign n4092 = n500 | n4091 ;
  assign n4093 = n618 | n4092 ;
  assign n4094 = n4060 | n4063 ;
  assign n4095 = n4055 | n4057 ;
  assign n4096 = n4036 | n4039 ;
  assign n4097 = n4020 | n4023 ;
  assign n4098 = ~n2561 & n2732 ;
  assign n4099 = n2720 & ~n3052 ;
  assign n4100 = n2564 & n2730 ;
  assign n4101 = n2569 & n2728 ;
  assign n4102 = n4100 | n4101 ;
  assign n4103 = n4099 | n4102 ;
  assign n4104 = n4098 | n4103 ;
  assign n4105 = n372 | n4104 ;
  assign n4106 = n372 & n4104 ;
  assign n4107 = n4105 & ~n4106 ;
  assign n4108 = n221 & ~n2581 ;
  assign n4109 = n2702 & ~n2823 ;
  assign n4110 = n2572 & n2697 ;
  assign n4111 = ~n2575 & n2695 ;
  assign n4112 = n2578 & n2793 ;
  assign n4113 = n4111 | n4112 ;
  assign n4114 = n4110 | n4113 ;
  assign n4115 = n4109 | n4114 ;
  assign n4116 = n4108 & n4115 ;
  assign n4117 = n4108 | n4115 ;
  assign n4118 = ~n4116 & n4117 ;
  assign n4119 = n221 & ~n4009 ;
  assign n4120 = n2584 & n4119 ;
  assign n4121 = n4017 | n4120 ;
  assign n4122 = n4118 & n4121 ;
  assign n4123 = n4118 | n4121 ;
  assign n4124 = ~n4122 & n4123 ;
  assign n4125 = n4107 & n4124 ;
  assign n4126 = n4107 | n4124 ;
  assign n4127 = ~n4125 & n4126 ;
  assign n4128 = n4097 & n4127 ;
  assign n4129 = n4097 | n4127 ;
  assign n4130 = ~n4128 & n4129 ;
  assign n4131 = n2830 & ~n3329 ;
  assign n4132 = ~n2549 & n2832 ;
  assign n4133 = n2557 & n2840 ;
  assign n4134 = n2553 & n2837 ;
  assign n4135 = n4133 | n4134 ;
  assign n4136 = n4132 | n4135 ;
  assign n4137 = n4131 | n4136 ;
  assign n4138 = n903 & ~n4137 ;
  assign n4139 = ~n903 & n4137 ;
  assign n4140 = n4138 | n4139 ;
  assign n4141 = n4130 & n4140 ;
  assign n4142 = n4130 | n4140 ;
  assign n4143 = ~n4141 & n4142 ;
  assign n4144 = n4096 & n4143 ;
  assign n4145 = n4036 | n4143 ;
  assign n4146 = n4039 | n4145 ;
  assign n4147 = ~n4144 & n4146 ;
  assign n4148 = n3022 & ~n3694 ;
  assign n4149 = n3026 & ~n3701 ;
  assign n4150 = n2547 & n3032 ;
  assign n4151 = n2661 & n3034 ;
  assign n4152 = n4150 | n4151 ;
  assign n4153 = n4149 | n4152 ;
  assign n4154 = n4148 | n4153 ;
  assign n4155 = n1199 | n4154 ;
  assign n4156 = n1199 & n4154 ;
  assign n4157 = n4155 & ~n4156 ;
  assign n4158 = n4147 | n4157 ;
  assign n4159 = n4146 & n4157 ;
  assign n4160 = ~n4144 & n4159 ;
  assign n4161 = n4158 & ~n4160 ;
  assign n4162 = n2679 & ~n3835 ;
  assign n4163 = n2675 & ~n3981 ;
  assign n4164 = n4162 | n4163 ;
  assign n4165 = n29 & ~n4164 ;
  assign n4166 = ~n29 & n4164 ;
  assign n4167 = n4165 | n4166 ;
  assign n4168 = n4161 | n4167 ;
  assign n4169 = ~n4160 & n4167 ;
  assign n4170 = n4158 & n4169 ;
  assign n4171 = n4168 & ~n4170 ;
  assign n4172 = n4095 | n4171 ;
  assign n4173 = n4095 & ~n4170 ;
  assign n4174 = n4168 & n4173 ;
  assign n4175 = n4172 & ~n4174 ;
  assign n4176 = n4094 & n4175 ;
  assign n4177 = n4094 | n4175 ;
  assign n4178 = ~n4176 & n4177 ;
  assign n4179 = n4093 | n4178 ;
  assign n4180 = n4093 & n4178 ;
  assign n4181 = n4179 & ~n4180 ;
  assign n4182 = n4080 & n4181 ;
  assign n4183 = n4080 | n4181 ;
  assign n4184 = ~n4182 & n4183 ;
  assign n4185 = n4072 & n4184 ;
  assign n4186 = n4072 | n4184 ;
  assign n4187 = ~n4185 & n4186 ;
  assign n4188 = n4079 & ~n4187 ;
  assign n4189 = ~n4079 & n4187 ;
  assign n4190 = n4188 | n4189 ;
  assign n4191 = n4180 | n4182 ;
  assign n4192 = n319 | n379 ;
  assign n4193 = n650 | n2158 ;
  assign n4194 = n2378 | n4193 ;
  assign n4195 = n4192 | n4194 ;
  assign n4196 = n143 | n2373 ;
  assign n4197 = n290 | n4196 ;
  assign n4198 = n206 | n2368 ;
  assign n4199 = n4197 | n4198 ;
  assign n4200 = n287 | n2381 ;
  assign n4201 = n444 | n4200 ;
  assign n4202 = n4199 | n4201 ;
  assign n4203 = n4195 | n4202 ;
  assign n4204 = n378 | n4203 ;
  assign n4205 = n889 | n1344 ;
  assign n4206 = n178 | n4205 ;
  assign n4207 = n645 | n4206 ;
  assign n4208 = n4204 | n4207 ;
  assign n4209 = n174 | n4208 ;
  assign n4210 = n480 | n4209 ;
  assign n4211 = n4174 | n4176 ;
  assign n4212 = n4160 | n4170 ;
  assign n4213 = n4125 | n4128 ;
  assign n4214 = n2557 & n2732 ;
  assign n4215 = n2720 & ~n3025 ;
  assign n4216 = ~n2561 & n2730 ;
  assign n4217 = n2564 & n2728 ;
  assign n4218 = n4216 | n4217 ;
  assign n4219 = n4215 | n4218 ;
  assign n4220 = n4214 | n4219 ;
  assign n4221 = n372 & n4220 ;
  assign n4222 = n372 | n4220 ;
  assign n4223 = ~n4221 & n4222 ;
  assign n4224 = n2569 & n2697 ;
  assign n4225 = n2702 & n2999 ;
  assign n4226 = n2572 & n2695 ;
  assign n4227 = ~n2575 & n2793 ;
  assign n4228 = n4226 | n4227 ;
  assign n4229 = n4225 | n4228 ;
  assign n4230 = n4224 | n4229 ;
  assign n4231 = n221 & ~n4230 ;
  assign n4232 = ~n221 & n4230 ;
  assign n4233 = n4231 | n4232 ;
  assign n4234 = n29 & n221 ;
  assign n4235 = n2578 & n4234 ;
  assign n4236 = n221 & n2578 ;
  assign n4237 = n29 | n4236 ;
  assign n4238 = ~n4235 & n4237 ;
  assign n4239 = n4233 & n4238 ;
  assign n4240 = n4233 | n4238 ;
  assign n4241 = ~n4239 & n4240 ;
  assign n4242 = n221 & ~n4115 ;
  assign n4243 = n2581 & n4242 ;
  assign n4244 = n4122 | n4243 ;
  assign n4245 = ~n4241 & n4244 ;
  assign n4246 = n4241 & ~n4244 ;
  assign n4247 = n4245 | n4246 ;
  assign n4248 = n4223 & n4247 ;
  assign n4249 = n4223 | n4247 ;
  assign n4250 = ~n4248 & n4249 ;
  assign n4251 = n4213 & n4250 ;
  assign n4252 = n4213 | n4250 ;
  assign n4253 = ~n4251 & n4252 ;
  assign n4254 = n2547 & n2832 ;
  assign n4255 = n2830 & ~n3314 ;
  assign n4256 = n2553 & n2840 ;
  assign n4257 = ~n2549 & n2837 ;
  assign n4258 = n4256 | n4257 ;
  assign n4259 = n4255 | n4258 ;
  assign n4260 = n4254 | n4259 ;
  assign n4261 = n903 & ~n4260 ;
  assign n4262 = ~n903 & n4260 ;
  assign n4263 = n4261 | n4262 ;
  assign n4264 = n4253 & n4263 ;
  assign n4265 = n4253 | n4263 ;
  assign n4266 = ~n4264 & n4265 ;
  assign n4267 = n4141 | n4144 ;
  assign n4268 = n4266 & n4267 ;
  assign n4269 = n4266 | n4267 ;
  assign n4270 = ~n4268 & n4269 ;
  assign n4271 = n3022 & ~n3835 ;
  assign n4272 = n2661 & n3032 ;
  assign n4273 = n3034 & ~n3694 ;
  assign n4274 = n4272 | n4273 ;
  assign n4275 = n3026 & n3841 ;
  assign n4276 = ~n3839 & n4275 ;
  assign n4277 = n4274 | n4276 ;
  assign n4278 = n4271 | n4277 ;
  assign n4279 = n1199 & n4278 ;
  assign n4280 = n1199 | n4278 ;
  assign n4281 = ~n4279 & n4280 ;
  assign n4282 = n4270 & n4281 ;
  assign n4283 = n4270 | n4281 ;
  assign n4284 = ~n4282 & n4283 ;
  assign n4285 = n4212 & n4284 ;
  assign n4286 = n4212 | n4284 ;
  assign n4287 = ~n4285 & n4286 ;
  assign n4288 = n4211 & n4287 ;
  assign n4289 = n4174 | n4287 ;
  assign n4290 = n4176 | n4289 ;
  assign n4291 = ~n4288 & n4290 ;
  assign n4292 = n4210 | n4291 ;
  assign n4293 = n4210 & n4291 ;
  assign n4294 = n4292 & ~n4293 ;
  assign n4295 = n4191 & n4294 ;
  assign n4296 = n4191 | n4294 ;
  assign n4297 = ~n4295 & n4296 ;
  assign n4298 = n4185 | n4297 ;
  assign n4299 = n4185 & n4297 ;
  assign n4300 = n4298 & ~n4299 ;
  assign n4301 = n4078 | n4187 ;
  assign n4302 = n3811 & n4301 ;
  assign n4303 = ~n4300 & n4302 ;
  assign n4304 = n4300 & ~n4302 ;
  assign n4305 = n4303 | n4304 ;
  assign n4306 = n4293 | n4295 ;
  assign n4307 = n155 | n178 ;
  assign n4308 = n248 | n2491 ;
  assign n4309 = n252 | n4308 ;
  assign n4310 = n150 | n604 ;
  assign n4311 = n203 | n4310 ;
  assign n4312 = n261 | n402 ;
  assign n4313 = n311 | n4312 ;
  assign n4314 = n2211 | n4313 ;
  assign n4315 = n3822 | n4314 ;
  assign n4316 = n4311 | n4315 ;
  assign n4317 = n3934 | n4316 ;
  assign n4318 = n4309 | n4317 ;
  assign n4319 = n125 | n4318 ;
  assign n4320 = n4307 | n4319 ;
  assign n4321 = n2028 | n4320 ;
  assign n4322 = n510 | n4321 ;
  assign n4323 = n4285 | n4288 ;
  assign n4324 = n4268 | n4282 ;
  assign n4325 = n4251 | n4264 ;
  assign n4326 = n2661 & n2832 ;
  assign n4327 = n2667 & n2830 ;
  assign n4328 = ~n2549 & n2840 ;
  assign n4329 = n2547 & n2837 ;
  assign n4330 = n4328 | n4329 ;
  assign n4331 = n4327 | n4330 ;
  assign n4332 = n4326 | n4331 ;
  assign n4333 = n903 & ~n4332 ;
  assign n4334 = ~n903 & n4332 ;
  assign n4335 = n4333 | n4334 ;
  assign n4336 = n4241 & n4244 ;
  assign n4337 = n4248 | n4336 ;
  assign n4338 = n4235 | n4239 ;
  assign n4339 = ~n2575 & n4234 ;
  assign n4340 = n221 & ~n2575 ;
  assign n4341 = n29 | n4340 ;
  assign n4342 = ~n4339 & n4341 ;
  assign n4343 = n4338 & n4342 ;
  assign n4344 = n4338 | n4342 ;
  assign n4345 = ~n4343 & n4344 ;
  assign n4346 = n2564 & n2697 ;
  assign n4347 = n2702 & n3064 ;
  assign n4348 = n2569 & n2695 ;
  assign n4349 = n2572 & n2793 ;
  assign n4350 = n4348 | n4349 ;
  assign n4351 = n4347 | n4350 ;
  assign n4352 = n4346 | n4351 ;
  assign n4353 = n221 | n4352 ;
  assign n4354 = n221 & n4352 ;
  assign n4355 = n4353 & ~n4354 ;
  assign n4356 = n4345 & n4355 ;
  assign n4357 = n4345 | n4355 ;
  assign n4358 = ~n4356 & n4357 ;
  assign n4359 = n2720 & n3293 ;
  assign n4360 = n2553 & n2732 ;
  assign n4361 = n2557 & n2730 ;
  assign n4362 = ~n2561 & n2728 ;
  assign n4363 = n4361 | n4362 ;
  assign n4364 = n4360 | n4363 ;
  assign n4365 = n4359 | n4364 ;
  assign n4366 = n372 & ~n4365 ;
  assign n4367 = ~n372 & n4365 ;
  assign n4368 = n4366 | n4367 ;
  assign n4369 = n4358 & n4368 ;
  assign n4370 = n4358 | n4368 ;
  assign n4371 = ~n4369 & n4370 ;
  assign n4372 = n4337 & n4371 ;
  assign n4373 = n4337 | n4371 ;
  assign n4374 = ~n4372 & n4373 ;
  assign n4375 = n4335 & n4374 ;
  assign n4376 = n4335 | n4374 ;
  assign n4377 = ~n4375 & n4376 ;
  assign n4378 = n4325 & n4377 ;
  assign n4379 = n4325 | n4377 ;
  assign n4380 = ~n4378 & n4379 ;
  assign n4381 = n3032 & ~n3694 ;
  assign n4382 = n3034 & ~n3835 ;
  assign n4383 = n3026 & n3983 ;
  assign n4384 = n4382 | n4383 ;
  assign n4385 = n4381 | n4384 ;
  assign n4386 = n1199 & ~n4385 ;
  assign n4387 = ~n1199 & n4385 ;
  assign n4388 = n4386 | n4387 ;
  assign n4389 = n4380 & n4388 ;
  assign n4390 = n4380 | n4388 ;
  assign n4391 = ~n4389 & n4390 ;
  assign n4392 = n4324 & n4391 ;
  assign n4393 = n4324 | n4391 ;
  assign n4394 = ~n4392 & n4393 ;
  assign n4395 = n4323 & n4394 ;
  assign n4396 = n4323 | n4394 ;
  assign n4397 = ~n4395 & n4396 ;
  assign n4398 = n4322 | n4397 ;
  assign n4399 = n4322 & n4397 ;
  assign n4400 = n4398 & ~n4399 ;
  assign n4401 = n4306 & n4400 ;
  assign n4402 = n4293 | n4400 ;
  assign n4403 = n4295 | n4402 ;
  assign n4404 = ~n4401 & n4403 ;
  assign n4405 = n4299 | n4404 ;
  assign n4406 = n4299 & n4404 ;
  assign n4407 = n4405 & ~n4406 ;
  assign n4408 = n4300 | n4301 ;
  assign n4409 = n3811 & n4408 ;
  assign n4410 = ~n4407 & n4409 ;
  assign n4411 = n4407 & ~n4409 ;
  assign n4412 = n4410 | n4411 ;
  assign n4413 = n4399 | n4401 ;
  assign n4414 = n882 | n2374 ;
  assign n4415 = n3580 | n4414 ;
  assign n4416 = n2534 | n4415 ;
  assign n4417 = n143 | n4416 ;
  assign n4418 = n504 | n4417 ;
  assign n4419 = n855 | n2028 ;
  assign n4420 = n2038 | n2241 ;
  assign n4421 = n801 | n2338 ;
  assign n4422 = n1011 | n4421 ;
  assign n4423 = n478 | n4422 ;
  assign n4424 = n4420 | n4423 ;
  assign n4425 = n4419 | n4424 ;
  assign n4426 = n327 | n4425 ;
  assign n4427 = n193 | n4426 ;
  assign n4428 = n2149 | n4427 ;
  assign n4429 = n4418 | n4428 ;
  assign n4430 = n4392 | n4395 ;
  assign n4431 = n4378 | n4389 ;
  assign n4432 = n3032 & ~n3835 ;
  assign n4433 = n3026 & ~n3981 ;
  assign n4434 = n4432 | n4433 ;
  assign n4435 = ~n1199 & n4434 ;
  assign n4436 = n1199 & ~n4434 ;
  assign n4437 = n4435 | n4436 ;
  assign n4438 = n4372 | n4375 ;
  assign n4439 = n4437 & n4438 ;
  assign n4440 = n4437 | n4438 ;
  assign n4441 = ~n4439 & n4440 ;
  assign n4442 = n2832 & ~n3694 ;
  assign n4443 = n2830 & ~n3701 ;
  assign n4444 = n2547 & n2840 ;
  assign n4445 = n2661 & n2837 ;
  assign n4446 = n4444 | n4445 ;
  assign n4447 = n4443 | n4446 ;
  assign n4448 = n4442 | n4447 ;
  assign n4449 = n903 & ~n4448 ;
  assign n4450 = ~n903 & n4448 ;
  assign n4451 = n4449 | n4450 ;
  assign n4452 = n4356 | n4369 ;
  assign n4453 = n4339 | n4343 ;
  assign n4454 = n2572 & n4234 ;
  assign n4455 = n221 & n2572 ;
  assign n4456 = n29 | n4455 ;
  assign n4457 = ~n4454 & n4456 ;
  assign n4458 = n4453 & n4457 ;
  assign n4459 = n4453 | n4457 ;
  assign n4460 = ~n4458 & n4459 ;
  assign n4461 = ~n2561 & n2697 ;
  assign n4462 = n2702 & ~n3052 ;
  assign n4463 = n2564 & n2695 ;
  assign n4464 = n2569 & n2793 ;
  assign n4465 = n4463 | n4464 ;
  assign n4466 = n4462 | n4465 ;
  assign n4467 = n4461 | n4466 ;
  assign n4468 = n221 | n4467 ;
  assign n4469 = n221 & n4467 ;
  assign n4470 = n4468 & ~n4469 ;
  assign n4471 = n4460 & n4470 ;
  assign n4472 = n4460 | n4470 ;
  assign n4473 = ~n4471 & n4472 ;
  assign n4474 = n2720 & ~n3329 ;
  assign n4475 = ~n2549 & n2732 ;
  assign n4476 = n2553 & n2730 ;
  assign n4477 = n2557 & n2728 ;
  assign n4478 = n4476 | n4477 ;
  assign n4479 = n4475 | n4478 ;
  assign n4480 = n4474 | n4479 ;
  assign n4481 = n372 & ~n4480 ;
  assign n4482 = ~n372 & n4480 ;
  assign n4483 = n4481 | n4482 ;
  assign n4484 = n4473 & n4483 ;
  assign n4485 = n4473 | n4483 ;
  assign n4486 = ~n4484 & n4485 ;
  assign n4487 = n4452 & n4486 ;
  assign n4488 = n4452 | n4486 ;
  assign n4489 = ~n4487 & n4488 ;
  assign n4490 = n4451 & n4489 ;
  assign n4491 = n4451 | n4489 ;
  assign n4492 = ~n4490 & n4491 ;
  assign n4493 = n4441 & n4492 ;
  assign n4494 = n4441 | n4492 ;
  assign n4495 = ~n4493 & n4494 ;
  assign n4496 = n4431 & n4495 ;
  assign n4497 = n4431 | n4495 ;
  assign n4498 = ~n4496 & n4497 ;
  assign n4499 = n4430 & n4498 ;
  assign n4500 = n4430 | n4498 ;
  assign n4501 = ~n4499 & n4500 ;
  assign n4502 = n4429 | n4501 ;
  assign n4503 = n4429 & n4501 ;
  assign n4504 = n4502 & ~n4503 ;
  assign n4505 = n4413 & n4504 ;
  assign n4506 = n4399 | n4504 ;
  assign n4507 = n4401 | n4506 ;
  assign n4508 = ~n4505 & n4507 ;
  assign n4509 = n4406 & n4508 ;
  assign n4510 = n4406 | n4508 ;
  assign n4511 = ~n4509 & n4510 ;
  assign n4512 = n4407 | n4408 ;
  assign n4513 = n3811 & n4512 ;
  assign n4514 = ~n4511 & n4513 ;
  assign n4515 = n4511 & ~n4513 ;
  assign n4516 = n4514 | n4515 ;
  assign n4517 = n154 | n226 ;
  assign n4518 = n619 | n4313 ;
  assign n4519 = n103 | n4518 ;
  assign n4520 = n205 | n2135 ;
  assign n4521 = n230 | n4520 ;
  assign n4522 = n237 | n282 ;
  assign n4523 = n2065 | n4522 ;
  assign n4524 = n112 | n287 ;
  assign n4525 = n2048 | n4524 ;
  assign n4526 = n4523 | n4525 ;
  assign n4527 = n4521 | n4526 ;
  assign n4528 = n2132 | n3626 ;
  assign n4529 = n326 | n459 ;
  assign n4530 = n145 | n431 ;
  assign n4531 = n4529 | n4530 ;
  assign n4532 = n4528 | n4531 ;
  assign n4533 = n4527 | n4532 ;
  assign n4534 = n667 | n4533 ;
  assign n4535 = n2307 | n4534 ;
  assign n4536 = n4519 | n4535 ;
  assign n4537 = n4517 | n4536 ;
  assign n4538 = n174 | n4426 ;
  assign n4539 = n106 | n972 ;
  assign n4540 = n4538 | n4539 ;
  assign n4541 = n4537 | n4540 ;
  assign n4542 = n231 | n4541 ;
  assign n4543 = n4496 | n4499 ;
  assign n4544 = n4439 | n4493 ;
  assign n4545 = n2832 & ~n3835 ;
  assign n4546 = n2661 & n2840 ;
  assign n4547 = n2837 & ~n3694 ;
  assign n4548 = n4546 | n4547 ;
  assign n4549 = n2830 & n3841 ;
  assign n4550 = ~n3839 & n4549 ;
  assign n4551 = n4548 | n4550 ;
  assign n4552 = n4545 | n4551 ;
  assign n4553 = n903 | n4552 ;
  assign n4554 = n903 & n4552 ;
  assign n4555 = n4553 & ~n4554 ;
  assign n4556 = n4487 | n4490 ;
  assign n4557 = n4555 & n4556 ;
  assign n4558 = n4555 | n4556 ;
  assign n4559 = ~n4557 & n4558 ;
  assign n4560 = n4471 | n4484 ;
  assign n4561 = n2720 & ~n3314 ;
  assign n4562 = n2547 & n2732 ;
  assign n4563 = ~n2549 & n2730 ;
  assign n4564 = n2553 & n2728 ;
  assign n4565 = n4563 | n4564 ;
  assign n4566 = n4562 | n4565 ;
  assign n4567 = n4561 | n4566 ;
  assign n4568 = n372 | n4567 ;
  assign n4569 = n372 & n4567 ;
  assign n4570 = n4568 & ~n4569 ;
  assign n4571 = n4454 | n4458 ;
  assign n4572 = n221 & n2569 ;
  assign n4573 = n29 | n1199 ;
  assign n4574 = n29 & n1199 ;
  assign n4575 = n4573 & ~n4574 ;
  assign n4576 = n4572 & n4575 ;
  assign n4577 = n4572 | n4575 ;
  assign n4578 = ~n4576 & n4577 ;
  assign n4579 = n2702 & ~n3025 ;
  assign n4580 = n2557 & n2697 ;
  assign n4581 = ~n2561 & n2695 ;
  assign n4582 = n2564 & n2793 ;
  assign n4583 = n4581 | n4582 ;
  assign n4584 = n4580 | n4583 ;
  assign n4585 = n4579 | n4584 ;
  assign n4586 = n221 & ~n4585 ;
  assign n4587 = ~n221 & n4585 ;
  assign n4588 = n4586 | n4587 ;
  assign n4589 = n4578 & n4588 ;
  assign n4590 = n4578 | n4588 ;
  assign n4591 = ~n4589 & n4590 ;
  assign n4592 = n4571 & n4591 ;
  assign n4593 = n4571 | n4591 ;
  assign n4594 = ~n4592 & n4593 ;
  assign n4595 = n4570 & n4594 ;
  assign n4596 = n4570 | n4594 ;
  assign n4597 = ~n4595 & n4596 ;
  assign n4598 = n4560 & n4597 ;
  assign n4599 = n4560 | n4597 ;
  assign n4600 = ~n4598 & n4599 ;
  assign n4601 = n4559 & n4600 ;
  assign n4602 = n4559 | n4600 ;
  assign n4603 = ~n4601 & n4602 ;
  assign n4604 = n4544 & n4603 ;
  assign n4605 = n4544 | n4603 ;
  assign n4606 = ~n4604 & n4605 ;
  assign n4607 = n4543 & n4606 ;
  assign n4608 = n4543 | n4606 ;
  assign n4609 = ~n4607 & n4608 ;
  assign n4610 = n4542 & n4609 ;
  assign n4611 = n4542 | n4609 ;
  assign n4612 = ~n4610 & n4611 ;
  assign n4613 = n4503 | n4505 ;
  assign n4614 = n4612 & n4613 ;
  assign n4615 = n4612 | n4613 ;
  assign n4616 = ~n4614 & n4615 ;
  assign n4617 = n4509 & n4616 ;
  assign n4618 = n4509 | n4616 ;
  assign n4619 = ~n4617 & n4618 ;
  assign n4620 = n4511 | n4512 ;
  assign n4621 = n3811 & n4620 ;
  assign n4622 = ~n4619 & n4621 ;
  assign n4623 = n4619 & ~n4621 ;
  assign n4624 = n4622 | n4623 ;
  assign n4625 = n4610 | n4614 ;
  assign n4626 = n187 | n302 ;
  assign n4627 = n139 | n4626 ;
  assign n4628 = n474 | n2086 ;
  assign n4629 = n403 | n4628 ;
  assign n4630 = n201 | n4629 ;
  assign n4631 = n137 | n4630 ;
  assign n4632 = n4627 | n4631 ;
  assign n4633 = n266 | n4632 ;
  assign n4634 = n379 | n4633 ;
  assign n4635 = n3609 | n4634 ;
  assign n4636 = n858 | n2243 ;
  assign n4637 = n847 | n4636 ;
  assign n4638 = n4635 | n4637 ;
  assign n4639 = n197 | n398 ;
  assign n4640 = n126 | n4639 ;
  assign n4641 = n278 | n4640 ;
  assign n4642 = n2088 | n4641 ;
  assign n4643 = n4638 | n4642 ;
  assign n4644 = n227 | n4643 ;
  assign n4645 = n4557 | n4601 ;
  assign n4646 = n2840 & ~n3694 ;
  assign n4647 = n2837 & ~n3835 ;
  assign n4648 = n4646 | n4647 ;
  assign n4649 = n2830 & n3981 ;
  assign n4650 = ~n3982 & n4649 ;
  assign n4651 = n4648 | n4650 ;
  assign n4652 = ~n903 & n4651 ;
  assign n4653 = n903 & ~n4646 ;
  assign n4654 = ~n4647 & n4653 ;
  assign n4655 = ~n4650 & n4654 ;
  assign n4656 = n4652 | n4655 ;
  assign n4657 = n4595 | n4598 ;
  assign n4658 = n2661 & n2732 ;
  assign n4659 = n2667 & n2720 ;
  assign n4660 = n2547 & n2730 ;
  assign n4661 = ~n2549 & n2728 ;
  assign n4662 = n4660 | n4661 ;
  assign n4663 = n4659 | n4662 ;
  assign n4664 = n4658 | n4663 ;
  assign n4665 = n372 & n4664 ;
  assign n4666 = n372 | n4664 ;
  assign n4667 = ~n4665 & n4666 ;
  assign n4668 = n4589 | n4592 ;
  assign n4669 = n2702 & n3293 ;
  assign n4670 = n2553 & n2697 ;
  assign n4671 = n2557 & n2695 ;
  assign n4672 = ~n2561 & n2793 ;
  assign n4673 = n4671 | n4672 ;
  assign n4674 = n4670 | n4673 ;
  assign n4675 = n4669 | n4674 ;
  assign n4676 = n221 | n4675 ;
  assign n4677 = n221 & n4675 ;
  assign n4678 = n4676 & ~n4677 ;
  assign n4679 = n221 & n2564 ;
  assign n4680 = n4573 & ~n4576 ;
  assign n4681 = n4679 | n4680 ;
  assign n4682 = n4679 & n4680 ;
  assign n4683 = n4681 & ~n4682 ;
  assign n4684 = n4678 & n4683 ;
  assign n4685 = n4678 | n4683 ;
  assign n4686 = ~n4684 & n4685 ;
  assign n4687 = n4668 & n4686 ;
  assign n4688 = n4668 | n4686 ;
  assign n4689 = ~n4687 & n4688 ;
  assign n4690 = n4667 & n4689 ;
  assign n4691 = n4667 | n4689 ;
  assign n4692 = ~n4690 & n4691 ;
  assign n4693 = n4657 & n4692 ;
  assign n4694 = n4657 | n4692 ;
  assign n4695 = ~n4693 & n4694 ;
  assign n4696 = n4656 & n4695 ;
  assign n4697 = n4656 | n4695 ;
  assign n4698 = ~n4696 & n4697 ;
  assign n4699 = n4645 & n4698 ;
  assign n4700 = n4645 | n4698 ;
  assign n4701 = ~n4699 & n4700 ;
  assign n4702 = n4604 | n4607 ;
  assign n4703 = n4701 & n4702 ;
  assign n4704 = n4701 | n4702 ;
  assign n4705 = ~n4703 & n4704 ;
  assign n4706 = n4644 | n4705 ;
  assign n4707 = n4644 & n4705 ;
  assign n4708 = n4706 & ~n4707 ;
  assign n4709 = n4625 & n4708 ;
  assign n4710 = n4625 | n4708 ;
  assign n4711 = ~n4709 & n4710 ;
  assign n4712 = n4617 | n4711 ;
  assign n4713 = n4617 & n4711 ;
  assign n4714 = n4712 & ~n4713 ;
  assign n4715 = n4619 | n4620 ;
  assign n4716 = n3811 & n4715 ;
  assign n4717 = ~n4714 & n4716 ;
  assign n4718 = n4714 & ~n4716 ;
  assign n4719 = n4717 | n4718 ;
  assign n4720 = n4707 | n4709 ;
  assign n4721 = n193 | n2350 ;
  assign n4722 = n309 | n619 ;
  assign n4723 = n189 | n4722 ;
  assign n4724 = n671 | n4723 ;
  assign n4725 = n3558 | n4724 ;
  assign n4726 = n2534 | n4725 ;
  assign n4727 = n2479 | n4726 ;
  assign n4728 = n4721 | n4727 ;
  assign n4729 = n310 | n4728 ;
  assign n4730 = n139 | n4729 ;
  assign n4731 = n3626 | n4730 ;
  assign n4732 = n240 | n4731 ;
  assign n4733 = n333 | n4732 ;
  assign n4734 = n4699 | n4703 ;
  assign n4735 = n4693 | n4696 ;
  assign n4736 = n4687 | n4690 ;
  assign n4737 = n2840 & ~n3835 ;
  assign n4738 = n2830 & ~n3981 ;
  assign n4739 = n4737 | n4738 ;
  assign n4740 = n903 & ~n4739 ;
  assign n4741 = ~n903 & n4739 ;
  assign n4742 = n4740 | n4741 ;
  assign n4743 = n4736 & n4742 ;
  assign n4744 = n4736 | n4742 ;
  assign n4745 = ~n4743 & n4744 ;
  assign n4746 = n4681 & ~n4684 ;
  assign n4747 = n221 & ~n2567 ;
  assign n4748 = n2702 & ~n3329 ;
  assign n4749 = ~n2549 & n2697 ;
  assign n4750 = n2553 & n2695 ;
  assign n4751 = n2557 & n2793 ;
  assign n4752 = n4750 | n4751 ;
  assign n4753 = n4749 | n4752 ;
  assign n4754 = n4748 | n4753 ;
  assign n4755 = n221 & ~n4754 ;
  assign n4756 = ~n221 & n4754 ;
  assign n4757 = n4755 | n4756 ;
  assign n4758 = ~n4747 & n4757 ;
  assign n4759 = n4747 & ~n4757 ;
  assign n4760 = n4758 | n4759 ;
  assign n4761 = n4746 | n4760 ;
  assign n4762 = n4746 & n4760 ;
  assign n4763 = n4761 & ~n4762 ;
  assign n4764 = n2720 & ~n3701 ;
  assign n4765 = n2732 & ~n3694 ;
  assign n4766 = n2661 & n2730 ;
  assign n4767 = n2547 & n2728 ;
  assign n4768 = n4766 | n4767 ;
  assign n4769 = n4765 | n4768 ;
  assign n4770 = n4764 | n4769 ;
  assign n4771 = n372 & ~n4770 ;
  assign n4772 = ~n372 & n4770 ;
  assign n4773 = n4771 | n4772 ;
  assign n4774 = n4763 & n4773 ;
  assign n4775 = n4763 | n4773 ;
  assign n4776 = ~n4774 & n4775 ;
  assign n4777 = n4745 & n4776 ;
  assign n4778 = n4745 | n4776 ;
  assign n4779 = ~n4777 & n4778 ;
  assign n4780 = n4735 & n4779 ;
  assign n4781 = n4735 | n4779 ;
  assign n4782 = ~n4780 & n4781 ;
  assign n4783 = n4734 & n4782 ;
  assign n4784 = n4734 | n4782 ;
  assign n4785 = ~n4783 & n4784 ;
  assign n4786 = n4733 & n4785 ;
  assign n4787 = n4732 | n4785 ;
  assign n4788 = n333 | n4787 ;
  assign n4789 = ~n4786 & n4788 ;
  assign n4790 = n4720 | n4789 ;
  assign n4791 = n4720 & n4788 ;
  assign n4792 = ~n4786 & n4791 ;
  assign n4793 = n4790 & ~n4792 ;
  assign n4794 = n4713 | n4793 ;
  assign n4795 = n4713 & n4793 ;
  assign n4796 = n4794 & ~n4795 ;
  assign n4797 = n4714 | n4715 ;
  assign n4798 = n3811 & n4797 ;
  assign n4799 = ~n4796 & n4798 ;
  assign n4800 = n4796 & ~n4798 ;
  assign n4801 = n4799 | n4800 ;
  assign n4802 = n4786 | n4792 ;
  assign n4803 = n181 | n188 ;
  assign n4804 = n437 | n2027 ;
  assign n4805 = n856 | n2534 ;
  assign n4806 = n4804 | n4805 ;
  assign n4807 = n247 | n450 ;
  assign n4808 = n3623 | n3629 ;
  assign n4809 = n470 | n4808 ;
  assign n4810 = n3549 | n4809 ;
  assign n4811 = n4807 | n4810 ;
  assign n4812 = n334 | n4811 ;
  assign n4813 = n4806 | n4812 ;
  assign n4814 = n984 | n4813 ;
  assign n4815 = n4803 | n4814 ;
  assign n4816 = n316 | n4815 ;
  assign n4817 = n4743 | n4777 ;
  assign n4818 = n4761 & ~n4774 ;
  assign n4819 = n2720 & n3842 ;
  assign n4820 = n2732 & ~n3835 ;
  assign n4821 = n2730 & ~n3694 ;
  assign n4822 = n2661 & n2728 ;
  assign n4823 = n4821 | n4822 ;
  assign n4824 = n4820 | n4823 ;
  assign n4825 = n4819 | n4824 ;
  assign n4826 = n372 | n4825 ;
  assign n4827 = n372 & n4825 ;
  assign n4828 = n4826 & ~n4827 ;
  assign n4829 = ~n4818 & n4828 ;
  assign n4830 = n4818 & ~n4828 ;
  assign n4831 = n4829 | n4830 ;
  assign n4832 = n221 & n2557 ;
  assign n4833 = ~n903 & n4832 ;
  assign n4834 = n903 & ~n4832 ;
  assign n4835 = n4679 & ~n4834 ;
  assign n4836 = ~n4833 & n4835 ;
  assign n4837 = n4679 & ~n4836 ;
  assign n4838 = n4833 | n4836 ;
  assign n4839 = n4834 | n4838 ;
  assign n4840 = ~n4837 & n4839 ;
  assign n4841 = n221 & ~n2561 ;
  assign n4842 = ~n2564 & n4841 ;
  assign n4843 = n4758 | n4842 ;
  assign n4844 = ~n4840 & n4843 ;
  assign n4845 = n4840 & ~n4843 ;
  assign n4846 = n4844 | n4845 ;
  assign n4847 = n2702 & ~n3314 ;
  assign n4848 = n2547 & n2697 ;
  assign n4849 = ~n2549 & n2695 ;
  assign n4850 = n2553 & n2793 ;
  assign n4851 = n4849 | n4850 ;
  assign n4852 = n4848 | n4851 ;
  assign n4853 = n4847 | n4852 ;
  assign n4854 = n221 & ~n4853 ;
  assign n4855 = ~n221 & n4853 ;
  assign n4856 = n4854 | n4855 ;
  assign n4857 = ~n4846 & n4856 ;
  assign n4858 = n4846 & ~n4856 ;
  assign n4859 = n4857 | n4858 ;
  assign n4860 = n4831 | n4859 ;
  assign n4861 = n4831 & n4859 ;
  assign n4862 = n4860 & ~n4861 ;
  assign n4863 = n4817 & n4862 ;
  assign n4864 = n4817 | n4862 ;
  assign n4865 = ~n4863 & n4864 ;
  assign n4866 = n4780 | n4783 ;
  assign n4867 = n4865 & n4866 ;
  assign n4868 = n4865 | n4866 ;
  assign n4869 = ~n4867 & n4868 ;
  assign n4870 = n4816 | n4869 ;
  assign n4871 = n4816 & n4869 ;
  assign n4872 = n4870 & ~n4871 ;
  assign n4873 = n4802 & n4872 ;
  assign n4874 = n4802 | n4872 ;
  assign n4875 = ~n4873 & n4874 ;
  assign n4876 = n4795 | n4875 ;
  assign n4877 = n4795 & n4875 ;
  assign n4878 = n4876 & ~n4877 ;
  assign n4879 = n4796 | n4797 ;
  assign n4880 = n3811 & n4879 ;
  assign n4881 = ~n4878 & n4880 ;
  assign n4882 = n4878 & ~n4880 ;
  assign n4883 = n4881 | n4882 ;
  assign n4884 = n4871 | n4873 ;
  assign n4885 = n197 | n414 ;
  assign n4886 = n2236 | n4885 ;
  assign n4887 = n106 | n2235 ;
  assign n4888 = n193 | n283 ;
  assign n4889 = n121 | n235 ;
  assign n4890 = n4888 | n4889 ;
  assign n4891 = n161 | n510 ;
  assign n4892 = n379 | n390 ;
  assign n4893 = n4891 | n4892 ;
  assign n4894 = n4890 | n4893 ;
  assign n4895 = n231 | n500 ;
  assign n4896 = n244 | n248 ;
  assign n4897 = n4895 | n4896 ;
  assign n4898 = n164 | n380 ;
  assign n4899 = n202 | n302 ;
  assign n4900 = n4898 | n4899 ;
  assign n4901 = n4897 | n4900 ;
  assign n4902 = n4894 | n4901 ;
  assign n4903 = n207 | n397 ;
  assign n4904 = n386 | n4903 ;
  assign n4905 = n162 | n167 ;
  assign n4906 = n204 | n325 ;
  assign n4907 = n4905 | n4906 ;
  assign n4908 = n4904 | n4907 ;
  assign n4909 = n481 | n884 ;
  assign n4910 = n388 | n4909 ;
  assign n4911 = n322 | n396 ;
  assign n4912 = n189 | n192 ;
  assign n4913 = n4911 | n4912 ;
  assign n4914 = n4910 | n4913 ;
  assign n4915 = n4908 | n4914 ;
  assign n4916 = n4902 | n4915 ;
  assign n4917 = n4887 | n4916 ;
  assign n4918 = n4886 | n4917 ;
  assign n4919 = n114 | n277 ;
  assign n4920 = n4918 | n4919 ;
  assign n4921 = n4863 | n4867 ;
  assign n4922 = ~n4829 & n4860 ;
  assign n4923 = n2728 & ~n3694 ;
  assign n4924 = n2730 & ~n3835 ;
  assign n4925 = n2720 & n3983 ;
  assign n4926 = n4924 | n4925 ;
  assign n4927 = n4923 | n4926 ;
  assign n4928 = n372 & n4927 ;
  assign n4929 = n372 | n4927 ;
  assign n4930 = ~n4928 & n4929 ;
  assign n4931 = n4844 | n4857 ;
  assign n4932 = n221 & n2553 ;
  assign n4933 = n4838 & n4932 ;
  assign n4934 = n4838 | n4932 ;
  assign n4935 = ~n4933 & n4934 ;
  assign n4936 = n2667 & n2702 ;
  assign n4937 = n2661 & n2697 ;
  assign n4938 = n2547 & n2695 ;
  assign n4939 = ~n2549 & n2793 ;
  assign n4940 = n4938 | n4939 ;
  assign n4941 = n4937 | n4940 ;
  assign n4942 = n4936 | n4941 ;
  assign n4943 = n221 | n4942 ;
  assign n4944 = n221 & n4942 ;
  assign n4945 = n4943 & ~n4944 ;
  assign n4946 = ~n4935 & n4945 ;
  assign n4947 = n4935 & ~n4945 ;
  assign n4948 = n4946 | n4947 ;
  assign n4949 = n4931 & ~n4948 ;
  assign n4950 = ~n4931 & n4948 ;
  assign n4951 = n4949 | n4950 ;
  assign n4952 = n4930 & ~n4951 ;
  assign n4953 = ~n4930 & n4951 ;
  assign n4954 = n4952 | n4953 ;
  assign n4955 = n4922 | n4954 ;
  assign n4956 = n4922 & n4954 ;
  assign n4957 = n4955 & ~n4956 ;
  assign n4958 = n4921 & n4957 ;
  assign n4959 = n4921 | n4957 ;
  assign n4960 = ~n4958 & n4959 ;
  assign n4961 = n4920 | n4960 ;
  assign n4962 = n4920 & n4960 ;
  assign n4963 = n4961 & ~n4962 ;
  assign n4964 = n4884 & n4963 ;
  assign n4965 = n4884 | n4963 ;
  assign n4966 = ~n4964 & n4965 ;
  assign n4967 = n4877 | n4966 ;
  assign n4968 = n4877 & n4966 ;
  assign n4969 = n4967 & ~n4968 ;
  assign n4970 = n4878 | n4879 ;
  assign n4971 = n3811 & n4970 ;
  assign n4972 = ~n4969 & n4971 ;
  assign n4973 = n4969 & ~n4971 ;
  assign n4974 = n4972 | n4973 ;
  assign n4975 = n4962 | n4964 ;
  assign n4976 = n70 & n124 ;
  assign n4977 = n253 | n318 ;
  assign n4978 = n148 | n4977 ;
  assign n4979 = n197 | n4978 ;
  assign n4980 = n310 | n4979 ;
  assign n4981 = n2275 | n4980 ;
  assign n4982 = n827 | n4981 ;
  assign n4983 = n2157 | n3968 ;
  assign n4984 = n4982 | n4983 ;
  assign n4985 = n4976 | n4984 ;
  assign n4986 = n177 | n389 ;
  assign n4987 = n379 | n4986 ;
  assign n4988 = n294 | n4987 ;
  assign n4989 = n4985 | n4988 ;
  assign n4990 = n260 | n315 ;
  assign n4991 = n252 | n2032 ;
  assign n4992 = n311 | n4991 ;
  assign n4993 = n4990 | n4992 ;
  assign n4994 = n240 | n326 ;
  assign n4995 = n224 | n229 ;
  assign n4996 = n4994 | n4995 ;
  assign n4997 = n4993 | n4996 ;
  assign n4998 = n327 | n446 ;
  assign n4999 = n192 | n4998 ;
  assign n5000 = n4997 | n4999 ;
  assign n5001 = n4989 | n5000 ;
  assign n5002 = n4955 & ~n4958 ;
  assign n5003 = n4949 | n4952 ;
  assign n5004 = n4838 & ~n4932 ;
  assign n5005 = n4946 | n5004 ;
  assign n5006 = n221 & ~n2549 ;
  assign n5007 = n4932 & ~n5006 ;
  assign n5008 = ~n4932 & n5006 ;
  assign n5009 = n5005 & ~n5008 ;
  assign n5010 = ~n5007 & n5009 ;
  assign n5011 = n5005 & ~n5010 ;
  assign n5012 = n5007 | n5010 ;
  assign n5013 = n5008 | n5012 ;
  assign n5014 = ~n5011 & n5013 ;
  assign n5015 = n2702 & ~n3701 ;
  assign n5016 = n2697 & ~n3694 ;
  assign n5017 = n2661 & n2695 ;
  assign n5018 = n2547 & n2793 ;
  assign n5019 = n5017 | n5018 ;
  assign n5020 = n5016 | n5019 ;
  assign n5021 = n5015 | n5020 ;
  assign n5022 = n221 & ~n5021 ;
  assign n5023 = ~n221 & n5021 ;
  assign n5024 = n5022 | n5023 ;
  assign n5025 = n2720 & ~n3981 ;
  assign n5026 = n2728 & ~n3835 ;
  assign n5027 = n5025 | n5026 ;
  assign n5028 = n372 & ~n5027 ;
  assign n5029 = ~n372 & n5027 ;
  assign n5030 = n5028 | n5029 ;
  assign n5031 = n5024 & n5030 ;
  assign n5032 = n5024 | n5030 ;
  assign n5033 = ~n5031 & n5032 ;
  assign n5034 = ~n5014 & n5033 ;
  assign n5035 = n5014 & ~n5033 ;
  assign n5036 = n5034 | n5035 ;
  assign n5037 = n5003 & ~n5036 ;
  assign n5038 = ~n5003 & n5036 ;
  assign n5039 = n5037 | n5038 ;
  assign n5040 = n5002 | n5039 ;
  assign n5041 = n5002 & n5039 ;
  assign n5042 = n5040 & ~n5041 ;
  assign n5043 = n5001 | n5042 ;
  assign n5044 = n5001 & n5042 ;
  assign n5045 = n5043 & ~n5044 ;
  assign n5046 = n4975 & n5045 ;
  assign n5047 = n4975 | n5045 ;
  assign n5048 = ~n5046 & n5047 ;
  assign n5049 = n4968 | n5048 ;
  assign n5050 = n4968 & n5048 ;
  assign n5051 = n5049 & ~n5050 ;
  assign n5052 = n4969 | n4970 ;
  assign n5053 = n3811 & n5052 ;
  assign n5054 = ~n5051 & n5053 ;
  assign n5055 = n5051 & ~n5053 ;
  assign n5056 = n5054 | n5055 ;
  assign n5057 = n5044 | n5046 ;
  assign n5058 = n112 | n430 ;
  assign n5059 = n1357 | n2081 ;
  assign n5060 = n199 | n5059 ;
  assign n5061 = n249 | n267 ;
  assign n5062 = n991 | n2205 ;
  assign n5063 = n160 | n5062 ;
  assign n5064 = n5061 | n5063 ;
  assign n5065 = n5060 | n5064 ;
  assign n5066 = n226 | n2038 ;
  assign n5067 = n3934 | n5066 ;
  assign n5068 = n396 | n510 ;
  assign n5069 = n374 | n5068 ;
  assign n5070 = n5067 | n5069 ;
  assign n5071 = n132 | n317 ;
  assign n5072 = n174 | n5071 ;
  assign n5073 = n240 | n859 ;
  assign n5074 = n230 | n333 ;
  assign n5075 = n5073 | n5074 ;
  assign n5076 = n5072 | n5075 ;
  assign n5077 = n5070 | n5076 ;
  assign n5078 = n5065 | n5077 ;
  assign n5079 = n5058 | n5078 ;
  assign n5080 = n235 | n338 ;
  assign n5081 = n284 | n5080 ;
  assign n5082 = n5079 | n5081 ;
  assign n5083 = n397 | n5082 ;
  assign n5084 = ~n5037 & n5040 ;
  assign n5085 = n5031 | n5034 ;
  assign n5086 = n221 & n2547 ;
  assign n5087 = ~n372 & n5006 ;
  assign n5088 = n372 & ~n5006 ;
  assign n5089 = n5087 | n5088 ;
  assign n5090 = n5086 & ~n5089 ;
  assign n5091 = ~n5086 & n5089 ;
  assign n5092 = n5090 | n5091 ;
  assign n5093 = n2702 & n3842 ;
  assign n5094 = n2697 & ~n3835 ;
  assign n5095 = n2695 & ~n3694 ;
  assign n5096 = n2661 & n2793 ;
  assign n5097 = n5095 | n5096 ;
  assign n5098 = n5094 | n5097 ;
  assign n5099 = n5093 | n5098 ;
  assign n5100 = n221 & ~n5099 ;
  assign n5101 = ~n221 & n5099 ;
  assign n5102 = n5100 | n5101 ;
  assign n5103 = ~n5092 & n5102 ;
  assign n5104 = n5092 & ~n5102 ;
  assign n5105 = n5103 | n5104 ;
  assign n5106 = n5012 & ~n5105 ;
  assign n5107 = ~n5012 & n5105 ;
  assign n5108 = n5106 | n5107 ;
  assign n5109 = n5085 & ~n5108 ;
  assign n5110 = ~n5085 & n5108 ;
  assign n5111 = n5109 | n5110 ;
  assign n5112 = n5084 | n5111 ;
  assign n5113 = ~n5037 & n5111 ;
  assign n5114 = n5040 & n5113 ;
  assign n5115 = n5112 & ~n5114 ;
  assign n5116 = n5083 & n5115 ;
  assign n5117 = n5083 | n5115 ;
  assign n5118 = ~n5116 & n5117 ;
  assign n5119 = n5057 & n5118 ;
  assign n5120 = n5057 | n5118 ;
  assign n5121 = ~n5119 & n5120 ;
  assign n5122 = n5050 | n5121 ;
  assign n5123 = n5050 & n5121 ;
  assign n5124 = n5122 & ~n5123 ;
  assign n5125 = n5051 | n5052 ;
  assign n5126 = n3811 & n5125 ;
  assign n5127 = ~n5124 & n5126 ;
  assign n5128 = n5124 & ~n5126 ;
  assign n5129 = n5127 | n5128 ;
  assign n5130 = n5116 | n5119 ;
  assign n5131 = n283 | n293 ;
  assign n5132 = n114 | n5131 ;
  assign n5133 = n255 | n2088 ;
  assign n5134 = n240 | n2087 ;
  assign n5135 = n853 | n5134 ;
  assign n5136 = n5133 | n5135 ;
  assign n5137 = n155 | n1372 ;
  assign n5138 = n396 | n5137 ;
  assign n5139 = n2084 | n5138 ;
  assign n5140 = n2275 | n2351 ;
  assign n5141 = n325 | n496 ;
  assign n5142 = n167 | n5141 ;
  assign n5143 = n5140 | n5142 ;
  assign n5144 = n5139 | n5143 ;
  assign n5145 = n2368 | n3964 ;
  assign n5146 = n272 | n444 ;
  assign n5147 = n470 | n5146 ;
  assign n5148 = n5145 | n5147 ;
  assign n5149 = n5144 | n5148 ;
  assign n5150 = n2090 | n5149 ;
  assign n5151 = n119 | n2534 ;
  assign n5152 = n5150 | n5151 ;
  assign n5153 = n5136 | n5152 ;
  assign n5154 = n142 | n165 ;
  assign n5155 = n5153 | n5154 ;
  assign n5156 = n5132 | n5155 ;
  assign n5157 = n328 | n5156 ;
  assign n5158 = n2014 & ~n2691 ;
  assign n5159 = ~n2694 & n5158 ;
  assign n5160 = ~n3694 & n5159 ;
  assign n5161 = n2695 & ~n3835 ;
  assign n5162 = n2702 & n3983 ;
  assign n5163 = n5161 | n5162 ;
  assign n5164 = n5160 | n5163 ;
  assign n5165 = n221 | n5164 ;
  assign n5166 = n221 & n5164 ;
  assign n5167 = n5165 & ~n5166 ;
  assign n5168 = n221 & n2661 ;
  assign n5169 = n5087 | n5090 ;
  assign n5170 = ~n5168 & n5169 ;
  assign n5171 = ~n5087 & n5168 ;
  assign n5172 = ~n5090 & n5171 ;
  assign n5173 = n5170 | n5172 ;
  assign n5174 = n5167 & ~n5173 ;
  assign n5175 = ~n5167 & n5173 ;
  assign n5176 = n5174 | n5175 ;
  assign n5177 = n5103 | n5106 ;
  assign n5178 = ~n5176 & n5177 ;
  assign n5179 = n5176 & ~n5177 ;
  assign n5180 = n5178 | n5179 ;
  assign n5181 = ~n5109 & n5112 ;
  assign n5182 = n5180 | n5181 ;
  assign n5183 = n5180 & n5181 ;
  assign n5184 = n5182 & ~n5183 ;
  assign n5185 = n5157 | n5184 ;
  assign n5186 = n5157 & n5184 ;
  assign n5187 = n5185 & ~n5186 ;
  assign n5188 = n5130 & n5187 ;
  assign n5189 = n5130 | n5187 ;
  assign n5190 = ~n5188 & n5189 ;
  assign n5191 = n5123 | n5190 ;
  assign n5192 = n5123 & n5190 ;
  assign n5193 = n5191 & ~n5192 ;
  assign n5194 = n5124 | n5125 ;
  assign n5195 = n3811 & n5194 ;
  assign n5196 = ~n5193 & n5195 ;
  assign n5197 = n5193 & ~n5195 ;
  assign n5198 = n5196 | n5197 ;
  assign n5199 = n5186 | n5188 ;
  assign n5200 = n283 | n332 ;
  assign n5201 = n1015 | n5200 ;
  assign n5202 = n230 | n340 ;
  assign n5203 = n149 | n236 ;
  assign n5204 = n5202 | n5203 ;
  assign n5205 = n5201 | n5204 ;
  assign n5206 = n227 | n315 ;
  assign n5207 = n785 | n5206 ;
  assign n5208 = n165 | n248 ;
  assign n5209 = n461 | n5208 ;
  assign n5210 = n5207 | n5209 ;
  assign n5211 = n5205 | n5210 ;
  assign n5212 = n374 | n3564 ;
  assign n5213 = n2284 | n5212 ;
  assign n5214 = n386 | n811 ;
  assign n5215 = n279 | n445 ;
  assign n5216 = n1046 | n5215 ;
  assign n5217 = n193 | n5216 ;
  assign n5218 = n1044 | n5217 ;
  assign n5219 = n198 | n5218 ;
  assign n5220 = n5214 | n5219 ;
  assign n5221 = n174 | n650 ;
  assign n5222 = n132 | n4980 ;
  assign n5223 = n5221 | n5222 ;
  assign n5224 = n5220 | n5223 ;
  assign n5225 = n5213 | n5224 ;
  assign n5226 = n5211 | n5225 ;
  assign n5227 = n142 | n240 ;
  assign n5228 = n328 | n5227 ;
  assign n5229 = n5226 | n5228 ;
  assign n5230 = n456 | n5229 ;
  assign n5231 = n584 | n5230 ;
  assign n5232 = n5170 | n5174 ;
  assign n5233 = n221 & ~n3697 ;
  assign n5234 = n2793 & ~n3835 ;
  assign n5235 = n2702 & ~n3981 ;
  assign n5236 = n5234 | n5235 ;
  assign n5237 = n221 & ~n5236 ;
  assign n5238 = ~n221 & n5236 ;
  assign n5239 = n5237 | n5238 ;
  assign n5240 = ~n5233 & n5239 ;
  assign n5241 = n5233 & ~n5239 ;
  assign n5242 = n5240 | n5241 ;
  assign n5243 = ~n5232 & n5242 ;
  assign n5244 = n5232 & ~n5242 ;
  assign n5245 = n5243 | n5244 ;
  assign n5246 = ~n5178 & n5182 ;
  assign n5247 = n5245 & n5246 ;
  assign n5248 = n5245 | n5246 ;
  assign n5249 = ~n5247 & n5248 ;
  assign n5250 = n5231 & n5249 ;
  assign n5251 = n5231 | n5249 ;
  assign n5252 = ~n5250 & n5251 ;
  assign n5253 = n5199 & n5252 ;
  assign n5254 = n5199 | n5252 ;
  assign n5255 = ~n5253 & n5254 ;
  assign n5256 = n5192 | n5255 ;
  assign n5257 = n5192 & n5255 ;
  assign n5258 = n5256 & ~n5257 ;
  assign n5259 = n5193 | n5194 ;
  assign n5260 = n3811 & n5259 ;
  assign n5261 = ~n5258 & n5260 ;
  assign n5262 = n5258 & ~n5260 ;
  assign n5263 = n5261 | n5262 ;
  assign n5264 = n5258 | n5259 ;
  assign n5265 = n3811 & n5264 ;
  assign n5266 = n5250 | n5253 ;
  assign n5267 = n294 | n396 ;
  assign n5268 = n432 | n2144 ;
  assign n5269 = n204 | n246 ;
  assign n5270 = n5268 | n5269 ;
  assign n5271 = n5267 | n5270 ;
  assign n5272 = n2213 | n3570 ;
  assign n5273 = n3646 | n5072 ;
  assign n5274 = n5272 | n5273 ;
  assign n5275 = n5271 | n5274 ;
  assign n5276 = n5061 | n5275 ;
  assign n5277 = n221 & ~n3694 ;
  assign n5278 = ~n2661 & n5277 ;
  assign n5279 = n5240 | n5278 ;
  assign n5280 = ~n5244 & n5248 ;
  assign n5281 = n2661 & ~n3835 ;
  assign n5282 = ~n2661 & n3835 ;
  assign n5283 = n5281 | n5282 ;
  assign n5284 = n221 & n5283 ;
  assign n5285 = ~n5280 & n5284 ;
  assign n5286 = n5244 | n5284 ;
  assign n5287 = n5248 & ~n5286 ;
  assign n5288 = n5285 | n5287 ;
  assign n5289 = ~n5279 & n5288 ;
  assign n5290 = n5279 & ~n5287 ;
  assign n5291 = ~n5285 & n5290 ;
  assign n5292 = n5289 | n5291 ;
  assign n5293 = n5276 | n5292 ;
  assign n5294 = n5276 & n5292 ;
  assign n5295 = n5293 & ~n5294 ;
  assign n5296 = n5266 & n5295 ;
  assign n5297 = n5266 | n5295 ;
  assign n5298 = ~n5296 & n5297 ;
  assign n5299 = n5257 & n5298 ;
  assign n5300 = n5257 | n5298 ;
  assign n5301 = ~n5299 & n5300 ;
  assign n5302 = n5265 & ~n5301 ;
  assign n5303 = ~n5265 & n5301 ;
  assign n5304 = n5302 | n5303 ;
  assign n5305 = n5294 | n5296 ;
  assign n5306 = n146 | n2038 ;
  assign n5307 = n809 | n5306 ;
  assign n5308 = n229 | n2491 ;
  assign n5309 = n164 | n331 ;
  assign n5310 = n5308 | n5309 ;
  assign n5311 = n252 | n272 ;
  assign n5312 = n118 | n248 ;
  assign n5313 = n5311 | n5312 ;
  assign n5314 = n5310 | n5313 ;
  assign n5315 = n5307 | n5314 ;
  assign n5316 = n521 | n2027 ;
  assign n5317 = n205 | n859 ;
  assign n5318 = n197 | n5317 ;
  assign n5319 = n5316 | n5318 ;
  assign n5320 = n5315 | n5319 ;
  assign n5321 = n463 | n5320 ;
  assign n5322 = n389 | n5321 ;
  assign n5323 = n5305 & n5322 ;
  assign n5324 = n5294 | n5322 ;
  assign n5325 = n5296 | n5324 ;
  assign n5326 = ~n5323 & n5325 ;
  assign n5327 = ~n5299 & n5326 ;
  assign n5328 = n5299 & ~n5326 ;
  assign n5329 = n5327 | n5328 ;
  assign n5330 = n5264 | n5301 ;
  assign n5331 = n3811 & n5330 ;
  assign n5332 = ~n5329 & n5331 ;
  assign n5333 = n5329 & ~n5331 ;
  assign n5334 = n5332 | n5333 ;
  assign n5335 = n5329 | n5330 ;
  assign n5336 = n3811 & n5335 ;
  assign n5337 = n5299 & n5326 ;
  assign n5338 = n197 | n327 ;
  assign n5339 = n500 | n5338 ;
  assign n5340 = n1060 | n2074 ;
  assign n5341 = n421 | n476 ;
  assign n5342 = n1038 | n5341 ;
  assign n5343 = n5340 | n5342 ;
  assign n5344 = n176 | n5343 ;
  assign n5345 = n165 | n3607 ;
  assign n5346 = n5344 | n5345 ;
  assign n5347 = n867 | n5346 ;
  assign n5348 = n5339 | n5347 ;
  assign n5349 = n5323 | n5348 ;
  assign n5350 = n5337 & n5349 ;
  assign n5351 = n5337 | n5349 ;
  assign n5352 = n5322 & n5348 ;
  assign n5353 = n5305 & n5352 ;
  assign n5354 = n5351 & ~n5353 ;
  assign n5355 = ~n5350 & n5354 ;
  assign n5356 = n5336 & ~n5355 ;
  assign n5357 = ~n5336 & n5355 ;
  assign n5358 = n5356 | n5357 ;
  assign n5359 = n313 | n325 ;
  assign n5360 = n390 | n4313 ;
  assign n5361 = n5218 | n5360 ;
  assign n5362 = n5359 | n5361 ;
  assign n5363 = n795 | n2457 ;
  assign n5364 = n145 | n3615 ;
  assign n5365 = n204 | n5364 ;
  assign n5366 = n5363 | n5365 ;
  assign n5367 = n5362 | n5366 ;
  assign n5368 = n160 | n5367 ;
  assign n5369 = n5353 | n5368 ;
  assign n5370 = n5353 & n5368 ;
  assign n5371 = n5369 & ~n5370 ;
  assign n5372 = n5350 | n5371 ;
  assign n5373 = n5350 & n5371 ;
  assign n5374 = n5372 & ~n5373 ;
  assign n5375 = n5335 | n5355 ;
  assign n5376 = n3811 & n5375 ;
  assign n5377 = ~n5374 & n5376 ;
  assign n5378 = n5374 & ~n5376 ;
  assign n5379 = n5377 | n5378 ;
  assign n5380 = n5374 | n5375 ;
  assign n5381 = n3811 & n5380 ;
  assign n5382 = n121 | n4634 ;
  assign n5383 = n154 | n3577 ;
  assign n5384 = n176 | n5383 ;
  assign n5385 = n5382 | n5384 ;
  assign n5386 = n150 | n181 ;
  assign n5387 = n174 | n288 ;
  assign n5388 = n374 | n5387 ;
  assign n5389 = n224 | n243 ;
  assign n5390 = n165 | n271 ;
  assign n5391 = n5389 | n5390 ;
  assign n5392 = n5388 | n5391 ;
  assign n5393 = n183 | n2028 ;
  assign n5394 = n874 | n5393 ;
  assign n5395 = n5392 | n5394 ;
  assign n5396 = n868 | n872 ;
  assign n5397 = n324 | n787 ;
  assign n5398 = n287 | n5397 ;
  assign n5399 = n862 | n5398 ;
  assign n5400 = n5396 | n5399 ;
  assign n5401 = n5395 | n5400 ;
  assign n5402 = n5386 | n5401 ;
  assign n5403 = n5385 | n5402 ;
  assign n5404 = n386 | n5403 ;
  assign n5405 = n5370 & n5404 ;
  assign n5406 = n5370 | n5404 ;
  assign n5407 = ~n5405 & n5406 ;
  assign n5408 = n5373 | n5407 ;
  assign n5409 = n5348 & n5406 ;
  assign n5410 = n5371 & n5409 ;
  assign n5411 = n5337 & n5410 ;
  assign n5412 = n5408 & ~n5411 ;
  assign n5413 = n5381 & ~n5412 ;
  assign n5414 = ~n5381 & n5412 ;
  assign n5415 = n5413 | n5414 ;
  assign n5416 = n5380 | n5412 ;
  assign n5417 = n3811 & n5416 ;
  assign n5418 = n168 | n445 ;
  assign n5419 = n226 | n5418 ;
  assign n5420 = n164 | n1030 ;
  assign n5421 = n315 | n5420 ;
  assign n5422 = n313 | n5421 ;
  assign n5423 = n5419 | n5422 ;
  assign n5424 = n320 | n651 ;
  assign n5425 = n291 | n849 ;
  assign n5426 = n160 | n5425 ;
  assign n5427 = n259 | n5426 ;
  assign n5428 = n5424 | n5427 ;
  assign n5429 = n132 | n227 ;
  assign n5430 = n131 | n150 ;
  assign n5431 = n235 | n310 ;
  assign n5432 = n163 | n5431 ;
  assign n5433 = n213 | n5432 ;
  assign n5434 = n5430 | n5433 ;
  assign n5435 = n145 | n230 ;
  assign n5436 = n142 | n430 ;
  assign n5437 = n134 | n261 ;
  assign n5438 = n5436 | n5437 ;
  assign n5439 = n5435 | n5438 ;
  assign n5440 = n5434 | n5439 ;
  assign n5441 = n5429 | n5440 ;
  assign n5442 = n5428 | n5441 ;
  assign n5443 = n260 | n314 ;
  assign n5444 = n139 | n155 ;
  assign n5445 = n174 | n5444 ;
  assign n5446 = n5443 | n5445 ;
  assign n5447 = n309 | n5446 ;
  assign n5448 = n5442 | n5447 ;
  assign n5449 = n5423 | n5448 ;
  assign n5450 = n402 | n5449 ;
  assign n5451 = n2170 | n5450 ;
  assign n5452 = n5405 | n5451 ;
  assign n5453 = n5405 & n5451 ;
  assign n5454 = n5452 & ~n5453 ;
  assign n5455 = n5411 & n5454 ;
  assign n5456 = n5411 | n5454 ;
  assign n5457 = ~n5455 & n5456 ;
  assign n5458 = n5417 & n5457 ;
  assign n5459 = n5417 | n5457 ;
  assign n5460 = ~n5458 & n5459 ;
  assign n5461 = n5416 | n5457 ;
  assign n5462 = n3811 & n5461 ;
  assign n5463 = n5411 | n5453 ;
  assign n5464 = n5452 & n5463 ;
  assign n5465 = n145 | n342 ;
  assign n5466 = n135 | n303 ;
  assign n5467 = n5418 | n5466 ;
  assign n5468 = n5465 | n5467 ;
  assign n5469 = n154 | n186 ;
  assign n5470 = n173 | n212 ;
  assign n5471 = n137 | n246 ;
  assign n5472 = n5470 | n5471 ;
  assign n5473 = n150 | n5472 ;
  assign n5474 = n337 | n5436 ;
  assign n5475 = n5420 | n5474 ;
  assign n5476 = n5473 | n5475 ;
  assign n5477 = n131 | n300 ;
  assign n5478 = n160 | n402 ;
  assign n5479 = n255 | n5478 ;
  assign n5480 = n163 | n5479 ;
  assign n5481 = n5477 | n5480 ;
  assign n5482 = n5476 | n5481 ;
  assign n5483 = n5469 | n5482 ;
  assign n5484 = n5468 | n5483 ;
  assign n5485 = n5445 | n5484 ;
  assign n5486 = n5464 & n5485 ;
  assign n5487 = n5464 | n5485 ;
  assign n5488 = ~n5486 & n5487 ;
  assign n5489 = n5462 & n5488 ;
  assign n5490 = n5462 | n5488 ;
  assign n5491 = ~n5489 & n5490 ;
  assign n5492 = ~n5462 & n5486 ;
  assign n5493 = pi21 | n62 ;
  assign n5494 = pi22 | n5493 ;
  assign n5495 = ~n5492 & n5494 ;
  assign n5496 = n4620 | n5485 ;
  assign n5497 = n4619 | n5496 ;
  assign n5498 = n4714 | n5497 ;
  assign n5499 = n4796 | n5498 ;
  assign n5500 = n4878 | n5499 ;
  assign n5501 = n4969 | n5500 ;
  assign n5502 = n5051 | n5501 ;
  assign n5503 = n5124 | n5502 ;
  assign n5504 = n5193 | n5503 ;
  assign n5505 = n5258 | n5504 ;
  assign n5506 = n5301 | n5505 ;
  assign n5507 = n5329 | n5506 ;
  assign n5508 = n5374 | n5507 ;
  assign n5509 = n5457 | n5508 ;
  assign n5510 = n5355 | n5412 ;
  assign n5511 = n5464 | n5510 ;
  assign n5512 = n5509 | n5511 ;
  assign n5513 = n3811 & n5512 ;
  assign n5514 = ~n5486 & n5513 ;
  assign n5515 = n5495 & ~n5514 ;
  assign n5516 = n5494 & ~n5512 ;
  assign n5517 = n3811 & ~n5516 ;
  assign po0 = n3808 ;
  assign po1 = n3957 ;
  assign po2 = n4077 ;
  assign po3 = n4190 ;
  assign po4 = n4305 ;
  assign po5 = n4412 ;
  assign po6 = n4516 ;
  assign po7 = n4624 ;
  assign po8 = n4719 ;
  assign po9 = n4801 ;
  assign po10 = n4883 ;
  assign po11 = n4974 ;
  assign po12 = n5056 ;
  assign po13 = n5129 ;
  assign po14 = n5198 ;
  assign po15 = n5263 ;
  assign po16 = n5304 ;
  assign po17 = n5334 ;
  assign po18 = n5358 ;
  assign po19 = n5379 ;
  assign po20 = n5415 ;
  assign po21 = n5460 ;
  assign po22 = n5491 ;
  assign po23 = ~n5515 ;
  assign po24 = n5517 ;
endmodule
