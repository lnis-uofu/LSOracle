/****************************************************************************
 *                                                                          *
 *  VERILOG VERSION of ORIGINAL NETLIST for c2670                           *
 *                                                                          *  
 *                                                                          *
 *  Generated by: Hakan Yalcin (hyalcin@cadence.com)                        *
 *                                                                          *
 *                Sep 16, 1998                                              *
 *                                                                          *
****************************************************************************/

module c2670g (
        L81, L92, L91, L90, L89, L88, L87, 
        L86, L85, L93, L43, L54, L53, L52, L51, 
        L50, L49, L48, L47, L55, L56, L66, L65, 
        L64, L63, L62, L61, L60, L67, L68, L79, 
        L78, L77, L76, L75, L74, L73, L72, L80, 
        L131, L141, L140, L139, L138, L137, L136, L135, 
        L142, L95, L105, L104, L103, L102, L101, L100, 
        L99, L106, L119, L129, L128, L127, L126, L125, 
        L124, L123, L130, L107, L117, L116, L115, L114, 
        L113, L112, L111, L118, L1971, L1966, L1961, L1956, 
        L1348, L1341, L2090, L2084, L2078, L2072, L2067, L1996, 
        L1991, L1986, L1981, L1976, L2096, L2100, L2678, L2474, 
        L2427, L2430, L2451, L2454, L2443, L2446, L2435, L2438, 
        L24, L6, L23, L22, L21, L5, L20, L4, 
        L19, L28, L35, L34, L27, L33, L26, L32, 
        L25, L651, L543, L2105, L2104, L1384, L40, L16, 
        L29, L11, L8, L37, L14, L44, L132, L82, 
        L96, L69, L120, L57, L108, L2106, L567, L559, 
        L860, L868, L452, L2066, L1083, L94, L7, L661, 
        L1, L2, L3, L15, L36, L483, L169, L174, 
        L177, L178, L179, L180, L181, L182, L183, L184, 
        L185, L186, L189, L190, L191, L192, L193, L194, 
        L195, L196, L197, L198, L199, L200, L201, L202, 
        L203, L204, L205, L206, L207, L208, L209, L210, 
        L211, L212, L213, L214, L215, L239, L240, L241, 
        L242, L243, L244, L245, L246, L247, L248, L249, 
        L250, L251, L252, L253, L254, L255, L256, L257, 
        L262, L263, L264, L265, L266, L267, L268, L269, 
        L270, L271, L272, L273, L274, L275, L276, L277, 
        L278, L279,
        L329, L231, L311, L150, L308, L225, L395, 
        L397, L227, L229, L401, L319, L325, L261, L220, 
        L221, L219, L218, L235, L236, L237, L238, L335, 
        L350, L391, L409, L337, L384, L411, L367, L369, 
        L173, L295, L331, L145, L148, L282, L323, L284, 
        L321, L297, L280, L153, L290, L305, L288, L303, 
        L286, L301, L299, L166, L168, L171, L162, L160, 
        L164, L156, L223, L217, L234, L259, L176, L188, 
        L158, L169o, L174o, L177o, L178o, L179o, L180o, L181o,
        L182o, L183o, L184o, L185o, L186o, L189o, L190o, L191o,
        L192o, L193o, L194o, L195o, L196o, L197o, L198o, L199o, 
        L200o, L201o, L202o, L203o, L204o, L205o, L206o, L207o, 
        L208o, L209o, L210o, L211o, L212o, L213o, L214o, L215o, 
        L239o, L240o, L241o, L242o, L243o, L244o, L245o, L246o, 
        L247o, L248o, L249o, L250o, L251o, L252o, L253o, L254o, 
        L255o, L256o, L257o, L262o, L263o, L264o, L265o, L266o, 
        L267o, L268o, L269o, L270o, L271o, L272o, L273o, L274o, 
        L275o, L276o, L277o, L278o, L279o);

 
   input
        L81, L92, L91, L90, L89, L88, L87, 
        L86, L85, L93, L43, L54, L53, L52, L51, 
        L50, L49, L48, L47, L55, L56, L66, L65, 
        L64, L63, L62, L61, L60, L67, L68, L79, 
        L78, L77, L76, L75, L74, L73, L72, L80, 
        L131, L141, L140, L139, L138, L137, L136, L135, 
        L142, L95, L105, L104, L103, L102, L101, L100, 
        L99, L106, L119, L129, L128, L127, L126, L125, 
        L124, L123, L130, L107, L117, L116, L115, L114, 
        L113, L112, L111, L118, L1971, L1966, L1961, L1956, 
        L1348, L1341, L2090, L2084, L2078, L2072, L2067, L1996, 
        L1991, L1986, L1981, L1976, L2096, L2100, L2678, L2474, 
        L2427, L2430, L2451, L2454, L2443, L2446, L2435, L2438, 
        L24, L6, L23, L22, L21, L5, L20, L4, 
        L19, L28, L35, L34, L27, L33, L26, L32, 
        L25, L651, L543, L2105, L2104, L1384, L40, L16, 
        L29, L11, L8, L37, L14, L44, L132, L82, 
        L96, L69, L120, L57, L108, L2106, L567, L559, 
        L860, L868, L452, L2066, L1083, L94, L7, L661, 
        L1, L2, L3, L15, L36, L483, L169, L174, 
        L177, L178, L179, L180, L181, L182, L183, L184, 
        L185, L186, L189, L190, L191, L192, L193, L194, 
        L195, L196, L197, L198, L199, L200, L201, L202, 
        L203, L204, L205, L206, L207, L208, L209, L210, 
        L211, L212, L213, L214, L215, L239, L240, L241, 
        L242, L243, L244, L245, L246, L247, L248, L249, 
        L250, L251, L252, L253, L254, L255, L256, L257, 
        L262, L263, L264, L265, L266, L267, L268, L269, 
        L270, L271, L272, L273, L274, L275, L276, L277, 
        L278, L279;
 
   output
        L329, L231, L311, L150, L308, L225, L395, 
        L397, L227, L229, L401, L319, L325, L261, L220, 
        L221, L219, L218, L235, L236, L237, L238, L335, 
        L350, L391, L409, L337, L384, L411, L367, L369, 
        L173, L295, L331, L145, L148, L282, L323, L284, 
        L321, L297, L280, L153, L290, L305, L288, L303, 
        L286, L301, L299, L166, L168, L171, L162, L160, 
        L164, L156, L223, L217, L234, L259, L176, L188, 
        L158, L169o, L174o, L177o, L178o, L179o, L180o, L181o, 
        L182o, L183o, L184o, L185o, L186o, L189o, L190o, L191o, 
        L192o, L193o, L194o, L195o, L196o, L197o, L198o, L199o, 
        L200o, L201o, L202o, L203o, L204o, L205o, L206o, L207o, 
        L208o, L209o, L210o, L211o, L212o, L213o, L214o, L215o, 
        L239o, L240o, L241o, L242o, L243o, L244o, L245o, L246o, 
        L247o, L248o, L249o, L250o, L251o, L252o, L253o, L254o, 
        L255o, L256o, L257o, L262o, L263o, L264o, L265o, L266o, 
        L267o, L268o, L269o, L270o, L271o, L272o, L273o, L274o, 
        L275o, L276o, L277o, L278o, L279o;


   assign L169o = L169; 
   assign L174o = L174; 
   assign L177o = L177; 
   assign L178o = L178; 
   assign L179o = L179; 
   assign L180o = L180; 
   assign L181o = L181; 
   assign L182o = L182; 
   assign L183o = L183; 
   assign L184o = L184; 
   assign L185o = L185; 
   assign L186o = L186; 
   assign L189o = L189; 
   assign L190o = L190; 
   assign L191o = L191; 
   assign L192o = L192; 
   assign L193o = L193; 
   assign L194o = L194; 
   assign L195o = L195; 
   assign L196o = L196; 
   assign L197o = L197; 
   assign L198o = L198; 
   assign L199o = L199; 
   assign L200o = L200; 
   assign L201o = L201; 
   assign L202o = L202; 
   assign L203o = L203; 
   assign L204o = L204; 
   assign L205o = L205; 
   assign L206o = L206; 
   assign L207o = L207; 
   assign L208o = L208; 
   assign L209o = L209; 
   assign L210o = L210; 
   assign L211o = L211; 
   assign L212o = L212; 
   assign L213o = L213; 
   assign L214o = L214; 
   assign L215o = L215; 
   assign L239o = L239; 
   assign L240o = L240; 
   assign L241o = L241; 
   assign L242o = L242; 
   assign L243o = L243; 
   assign L244o = L244; 
   assign L245o = L245; 
   assign L246o = L246; 
   assign L247o = L247; 
   assign L248o = L248; 
   assign L249o = L249; 
   assign L250o = L250; 
   assign L251o = L251; 
   assign L252o = L252; 
   assign L253o = L253; 
   assign L254o = L254; 
   assign L255o = L255; 
   assign L256o = L256; 
   assign L257o = L257; 
   assign L262o = L262; 
   assign L263o = L263; 
   assign L264o = L264; 
   assign L265o = L265; 
   assign L266o = L266; 
   assign L267o = L267; 
   assign L268o = L268; 
   assign L269o = L269; 
   assign L270o = L270; 
   assign L271o = L271; 
   assign L272o = L272; 
   assign L273o = L273; 
   assign L274o = L274; 
   assign L275o = L275; 
   assign L276o = L276; 
   assign L277o = L277; 
   assign L278o = L278; 
   assign L279o = L279; 


   buffer U77 ( L452, L350 ); 
   buffer U78 ( L452, L335 ); 
   buffer U79 ( L452, L409 ); 
   and2 U80 ( L1, L3, L546 ); 
   inv U81 ( L559, L560 ); 
   buffer U82 ( L1083, L369 ); 
   buffer U83 ( L1083, L367 ); 
   inv U84 ( L1384, L1385 ); 
   buffer U85 ( L2066, L411 ); 
   buffer U86 ( L2066, L337 ); 
   buffer U87 ( L2066, L384 ); 
   and4 U88 ( L2090, L2084, L2078, L2072, L157 ); 
   inv U89 ( L546, L547 ); 
   inv U90 ( L44, L218 ); 
   inv U91 ( L132, L219 ); 
   inv U92 ( L82, L220 ); 
   inv U93 ( L96, L221 ); 
   inv U94 ( L69, L235 ); 
   inv U95 ( L120, L236 ); 
   inv U96 ( L57, L237 ); 
   inv U97 ( L108, L238 ); 
   and3 U98 ( L2, L15, L661, L258 ); 
   buffer U99 ( L661, L480 ); 
   buffer U100 ( L37, L486 ); 
   buffer U101 ( L452, L654 ); 
   buffer U102 ( L8, L655 ); 
   buffer U103 ( L8, L658 ); 
   buffer U104 ( L543, L772 ); 
   buffer U105 ( L651, L795 ); 
   inv U106 ( L860, L865 ); 
   inv U107 ( L868, L875 ); 
   and2 U108 ( L11, L868, L882 ); 
   and4 U109 ( L132, L82, L96, L44, L1251 ); 
   and4 U110 ( L120, L57, L108, L69, L1254 ); 
   buffer U111 ( L543, L1261 ); 
   buffer U112 ( L651, L1284 ); 
   inv U113 ( L1341, L1344 ); 
   inv U114 ( L1348, L1351 ); 
   buffer U115 ( L2104, L1394 ); 
   buffer U116 ( L2105, L1418 ); 
   inv U117 ( L2427, L2433 ); 
   inv U118 ( L2430, L2434 ); 
   inv U119 ( L2435, L2441 ); 
   inv U120 ( L2438, L2442 ); 
   inv U121 ( L2443, L2449 ); 
   inv U122 ( L2446, L2450 ); 
   inv U123 ( L2474, L2478 ); 
   buffer U124 ( L2104, L1631 ); 
   buffer U125 ( L2105, L1655 ); 
   buffer U126 ( L16, L1710 ); 
   buffer U127 ( L16, L1721 ); 
   inv U128 ( L2678, L2682 ); 
   and2 U129 ( L7, L661, L1955 ); 
   inv U130 ( L1956, L1959 ); 
   inv U131 ( L1961, L1964 ); 
   inv U132 ( L1966, L1969 ); 
   inv U133 ( L1971, L1974 ); 
   inv U134 ( L1976, L1979 ); 
   inv U135 ( L1981, L1984 ); 
   inv U136 ( L1986, L1989 ); 
   inv U137 ( L1991, L1994 ); 
   inv U138 ( L1996, L1999 ); 
   buffer U139 ( L29, L2001 ); 
   buffer U140 ( L29, L2012 ); 
   inv U141 ( L2067, L2070 ); 
   inv U142 ( L2072, L2076 ); 
   inv U143 ( L2078, L2082 ); 
   inv U144 ( L2084, L2088 ); 
   inv U145 ( L2090, L2094 ); 
   inv U146 ( L2096, L2099 ); 
   inv U147 ( L2100, L2103 ); 
   inv U148 ( L2451, L2457 ); 
   inv U149 ( L2454, L2458 ); 
   buffer U150 ( L1348, L2461 ); 
   buffer U151 ( L1341, L2464 ); 
   buffer U152 ( L1956, L2471 ); 
   buffer U153 ( L1966, L2479 ); 
   buffer U154 ( L1961, L2482 ); 
   buffer U155 ( L1976, L2487 ); 
   buffer U156 ( L1971, L2490 ); 
   buffer U157 ( L1986, L2495 ); 
   buffer U158 ( L1981, L2498 ); 
   buffer U159 ( L1996, L2505 ); 
   buffer U160 ( L1991, L2508 ); 
   buffer U161 ( L2067, L2675 ); 
   buffer U162 ( L2078, L2683 ); 
   buffer U163 ( L2072, L2686 ); 
   buffer U164 ( L2090, L2691 ); 
   buffer U165 ( L2084, L2694 ); 
   buffer U166 ( L2100, L2699 ); 
   buffer U167 ( L2096, L2702 ); 
   inv U168 ( L157, L158 ); 
   inv U169 ( L258, L259 ); 
   inv U170 ( L486, L487 ); 
   buffer U171 ( L654, L391 ); 
   nand2 U172 ( L2430, L2433, L1475 ); 
   nand2 U173 ( L2427, L2434, L1476 ); 
   nand2 U174 ( L2438, L2441, L1484 ); 
   nand2 U175 ( L2435, L2442, L1485 ); 
   nand2 U176 ( L2446, L2449, L1493 ); 
   nand2 U177 ( L2443, L2450, L1494 ); 
   nand2 U178 ( L2454, L2457, L2459 ); 
   nand2 U179 ( L2451, L2458, L2460 ); 
   and2 U180 ( L94, L654, L173 ); 
   and2 U181 ( L2106, L1955, L216 ); 
   inv U182 ( L1955, L223 ); 
   nand2 U183 ( L567, L1955, L234 ); 
   inv U184 ( L1251, L1253 ); 
   inv U185 ( L1254, L1256 ); 
   and2 U186 ( L1254, L1251, L558 ); 
   buffer U187 ( L655, L748 ); 
   inv U188 ( L772, L784 ); 
   inv U189 ( L795, L807 ); 
   and3 U190 ( L80, L772, L795, L821 ); 
   and3 U191 ( L68, L772, L795, L825 ); 
   and3 U192 ( L79, L772, L795, L829 ); 
   and3 U193 ( L78, L772, L795, L833 ); 
   and3 U194 ( L77, L772, L795, L837 ); 
   and2 U195 ( L11, L875, L881 ); 
   buffer U196 ( L655, L994 ); 
   inv U197 ( L1261, L1273 ); 
   inv U198 ( L1284, L1296 ); 
   and3 U199 ( L76, L1261, L1284, L1310 ); 
   and3 U200 ( L75, L1261, L1284, L1314 ); 
   and3 U201 ( L74, L1261, L1284, L1318 ); 
   and3 U202 ( L73, L1261, L1284, L1322 ); 
   and3 U203 ( L72, L1261, L1284, L1326 ); 
   inv U204 ( L1394, L1406 ); 
   inv U205 ( L1418, L1430 ); 
   and3 U206 ( L114, L1394, L1418, L1444 ); 
   and3 U207 ( L113, L1394, L1418, L1448 ); 
   and3 U208 ( L112, L1394, L1418, L1452 ); 
   and3 U209 ( L111, L1394, L1418, L1456 ); 
   and2 U210 ( L1394, L1418, L1460 ); 
   nand2 U211 ( L1475, L1476, L1477 ); 
   nand2 U212 ( L1484, L1485, L1486 ); 
   nand2 U213 ( L1493, L1494, L1495 ); 
   inv U214 ( L2471, L2477 ); 
   nand2 U215 ( L2471, L2478, L1499 ); 
   inv U216 ( L2479, L2485 ); 
   inv U217 ( L2482, L2486 ); 
   inv U218 ( L2487, L2493 ); 
   inv U219 ( L2490, L2494 ); 
   inv U220 ( L1631, L1643 ); 
   inv U221 ( L1655, L1667 ); 
   and3 U222 ( L118, L1631, L1655, L1681 ); 
   and3 U223 ( L107, L1631, L1655, L1685 ); 
   and3 U224 ( L117, L1631, L1655, L1689 ); 
   and3 U225 ( L116, L1631, L1655, L1693 ); 
   and3 U226 ( L115, L1631, L1655, L1697 ); 
   inv U227 ( L1710, L1716 ); 
   inv U228 ( L1721, L1728 ); 
   inv U229 ( L2675, L2681 ); 
   nand2 U230 ( L2675, L2682, L1776 ); 
   inv U231 ( L2683, L2689 ); 
   inv U232 ( L2686, L2690 ); 
   inv U233 ( L2691, L2697 ); 
   inv U234 ( L2694, L2698 ); 
   buffer U235 ( L658, L1831 ); 
   buffer U236 ( L658, L1893 ); 
   inv U237 ( L2001, L2007 ); 
   inv U238 ( L2012, L2018 ); 
   inv U239 ( L2461, L2467 ); 
   inv U240 ( L2464, L2468 ); 
   inv U241 ( L2495, L2501 ); 
   inv U242 ( L2498, L2502 ); 
   inv U243 ( L2505, L2511 ); 
   inv U244 ( L2508, L2512 ); 
   nand2 U245 ( L2459, L2460, L2518 ); 
   buffer U246 ( L1344, L2551 ); 
   buffer U247 ( L1351, L2559 ); 
   buffer U248 ( L1959, L2567 ); 
   buffer U249 ( L1964, L2575 ); 
   buffer U250 ( L1969, L2583 ); 
   buffer U251 ( L1974, L2591 ); 
   buffer U252 ( L1979, L2599 ); 
   buffer U253 ( L1984, L2607 ); 
   buffer U254 ( L1989, L2615 ); 
   buffer U255 ( L1994, L2623 ); 
   inv U256 ( L2699, L2705 ); 
   inv U257 ( L2702, L2706 ); 
   buffer U258 ( L1999, L2735 ); 
   buffer U259 ( L2070, L2743 ); 
   buffer U260 ( L2076, L2751 ); 
   buffer U261 ( L2082, L2759 ); 
   buffer U262 ( L2088, L2767 ); 
   buffer U263 ( L2094, L2775 ); 
   inv U264 ( L216, L217 ); 
   and2 U265 ( L2106, L1253, L550 ); 
   and2 U266 ( L567, L1256, L552 ); 
   buffer U267 ( L558, L325 ); 
   or2 U268 ( L881, L882, L894 ); 
   nand2 U269 ( L2474, L2477, L1498 ); 
   nand2 U270 ( L2482, L2485, L1507 ); 
   nand2 U271 ( L2479, L2486, L1508 ); 
   nand2 U272 ( L2490, L2493, L1516 ); 
   nand2 U273 ( L2487, L2494, L1517 ); 
   nand2 U274 ( L2678, L2681, L1775 ); 
   nand2 U275 ( L2686, L2689, L1784 ); 
   nand2 U276 ( L2683, L2690, L1785 ); 
   nand2 U277 ( L2694, L2697, L1793 ); 
   nand2 U278 ( L2691, L2698, L1794 ); 
   nand2 U279 ( L2464, L2467, L2469 ); 
   nand2 U280 ( L2461, L2468, L2470 ); 
   nand2 U281 ( L2498, L2501, L2503 ); 
   nand2 U282 ( L2495, L2502, L2504 ); 
   nand2 U283 ( L2508, L2511, L2513 ); 
   nand2 U284 ( L2505, L2512, L2514 ); 
   nand2 U285 ( L2702, L2705, L2707 ); 
   nand2 U286 ( L2699, L2706, L2708 ); 
   inv U287 ( L558, L261 ); 
   inv U288 ( L550, L551 ); 
   inv U289 ( L552, L553 ); 
   and3 U290 ( L93, L784, L807, L818 ); 
   and3 U291 ( L55, L772, L807, L819 ); 
   and3 U292 ( L67, L784, L795, L820 ); 
   and3 U293 ( L81, L784, L807, L822 ); 
   and3 U294 ( L43, L772, L807, L823 ); 
   and3 U295 ( L56, L784, L795, L824 ); 
   and3 U296 ( L92, L784, L807, L826 ); 
   and3 U297 ( L54, L772, L807, L827 ); 
   and3 U298 ( L66, L784, L795, L828 ); 
   and3 U299 ( L91, L784, L807, L830 ); 
   and3 U300 ( L53, L772, L807, L831 ); 
   and3 U301 ( L65, L784, L795, L832 ); 
   and3 U302 ( L90, L784, L807, L834 ); 
   and3 U303 ( L52, L772, L807, L835 ); 
   and3 U304 ( L64, L784, L795, L836 ); 
   and3 U305 ( L89, L1273, L1296, L1307 ); 
   and3 U306 ( L51, L1261, L1296, L1308 ); 
   and3 U307 ( L63, L1273, L1284, L1309 ); 
   and3 U308 ( L88, L1273, L1296, L1311 ); 
   and3 U309 ( L50, L1261, L1296, L1312 ); 
   and3 U310 ( L62, L1273, L1284, L1313 ); 
   and3 U311 ( L87, L1273, L1296, L1315 ); 
   and3 U312 ( L49, L1261, L1296, L1316 ); 
   and2 U313 ( L1273, L1284, L1317 ); 
   and3 U314 ( L86, L1273, L1296, L1319 ); 
   and3 U315 ( L48, L1261, L1296, L1320 ); 
   and3 U316 ( L61, L1273, L1284, L1321 ); 
   and3 U317 ( L85, L1273, L1296, L1323 ); 
   and3 U318 ( L47, L1261, L1296, L1324 ); 
   and3 U319 ( L60, L1273, L1284, L1325 ); 
   and3 U320 ( L138, L1406, L1430, L1441 ); 
   and3 U321 ( L102, L1394, L1430, L1442 ); 
   and3 U322 ( L126, L1406, L1418, L1443 ); 
   and3 U323 ( L137, L1406, L1430, L1445 ); 
   and3 U324 ( L101, L1394, L1430, L1446 ); 
   and3 U325 ( L125, L1406, L1418, L1447 ); 
   and3 U326 ( L136, L1406, L1430, L1449 ); 
   and3 U327 ( L100, L1394, L1430, L1450 ); 
   and3 U328 ( L124, L1406, L1418, L1451 ); 
   and3 U329 ( L135, L1406, L1430, L1453 ); 
   and3 U330 ( L99, L1394, L1430, L1454 ); 
   and3 U331 ( L123, L1406, L1418, L1455 ); 
   and2 U332 ( L1406, L1430, L1457 ); 
   and2 U333 ( L1394, L1430, L1458 ); 
   and2 U334 ( L1406, L1418, L1459 ); 
   inv U335 ( L1477, L1481 ); 
   inv U336 ( L1486, L1490 ); 
   nand2 U337 ( L1498, L1499, L1500 ); 
   nand2 U338 ( L1507, L1508, L1509 ); 
   nand2 U339 ( L1516, L1517, L1518 ); 
   buffer U340 ( L1495, L1521 ); 
   buffer U341 ( L1495, L1525 ); 
   inv U342 ( L2551, L2557 ); 
   inv U343 ( L2559, L2565 ); 
   inv U344 ( L2567, L2573 ); 
   inv U345 ( L2575, L2581 ); 
   inv U346 ( L2583, L2589 ); 
   inv U347 ( L2591, L2597 ); 
   inv U348 ( L2599, L2605 ); 
   inv U349 ( L2607, L2613 ); 
   inv U350 ( L2615, L2621 ); 
   inv U351 ( L2623, L2629 ); 
   and3 U352 ( L142, L1643, L1667, L1678 ); 
   and3 U353 ( L106, L1631, L1667, L1679 ); 
   and3 U354 ( L130, L1643, L1655, L1680 ); 
   and3 U355 ( L131, L1643, L1667, L1682 ); 
   and3 U356 ( L95, L1631, L1667, L1683 ); 
   and3 U357 ( L119, L1643, L1655, L1684 ); 
   and3 U358 ( L141, L1643, L1667, L1686 ); 
   and3 U359 ( L105, L1631, L1667, L1687 ); 
   and3 U360 ( L129, L1643, L1655, L1688 ); 
   and3 U361 ( L140, L1643, L1667, L1690 ); 
   and3 U362 ( L104, L1631, L1667, L1691 ); 
   and3 U363 ( L128, L1643, L1655, L1692 ); 
   and3 U364 ( L139, L1643, L1667, L1694 ); 
   and3 U365 ( L103, L1631, L1667, L1695 ); 
   and3 U366 ( L127, L1643, L1655, L1696 ); 
   and2 U367 ( L19, L1716, L1734 ); 
   and2 U368 ( L4, L1716, L1736 ); 
   and2 U369 ( L20, L1716, L1738 ); 
   and2 U370 ( L5, L1716, L1740 ); 
   and2 U371 ( L21, L1728, L1742 ); 
   and2 U372 ( L22, L1728, L1744 ); 
   and2 U373 ( L23, L1728, L1746 ); 
   and2 U374 ( L6, L1728, L1748 ); 
   and2 U375 ( L24, L1728, L1750 ); 
   nand2 U376 ( L1775, L1776, L1777 ); 
   nand2 U377 ( L1784, L1785, L1786 ); 
   nand2 U378 ( L1793, L1794, L1795 ); 
   and2 U379 ( L25, L2007, L2023 ); 
   and2 U380 ( L32, L2007, L2025 ); 
   and2 U381 ( L26, L2007, L2027 ); 
   and2 U382 ( L33, L2007, L2029 ); 
   and2 U383 ( L27, L2018, L2031 ); 
   and2 U384 ( L34, L2018, L2033 ); 
   and2 U385 ( L35, L2018, L2035 ); 
   and2 U386 ( L28, L2018, L2037 ); 
   inv U387 ( L2735, L2741 ); 
   inv U388 ( L2743, L2749 ); 
   inv U389 ( L2751, L2757 ); 
   inv U390 ( L2759, L2765 ); 
   inv U391 ( L2767, L2773 ); 
   inv U392 ( L2775, L2781 ); 
   nand2 U393 ( L2469, L2470, L2515 ); 
   inv U394 ( L2518, L2522 ); 
   nand2 U395 ( L2513, L2514, L2525 ); 
   nand2 U396 ( L2503, L2504, L2528 ); 
   nand2 U397 ( L2707, L2708, L2730 ); 
   and2 U398 ( L551, L553, L554 ); 
   or4 U399 ( L818, L819, L820, L821, L838 ); 
   or4 U400 ( L822, L823, L824, L825, L841 ); 
   or4 U401 ( L826, L827, L828, L829, L846 ); 
   or4 U402 ( L830, L831, L832, L833, L854 ); 
   or4 U403 ( L834, L835, L836, L837, L857 ); 
   or4 U404 ( L1307, L1308, L1309, L1310, L1327 ); 
   or4 U405 ( L1311, L1312, L1313, L1314, L1329 ); 
   or4 U406 ( L1315, L1316, L1317, L1318, L1331 ); 
   or4 U407 ( L1319, L1320, L1321, L1322, L1333 ); 
   or4 U408 ( L1323, L1324, L1325, L1326, L1335 ); 
   or4 U409 ( L1441, L1442, L1443, L1444, L1461 ); 
   or4 U410 ( L1445, L1446, L1447, L1448, L1464 ); 
   or4 U411 ( L1449, L1450, L1451, L1452, L1467 ); 
   or4 U412 ( L1453, L1454, L1455, L1456, L1470 ); 
   or4 U413 ( L1457, L1458, L1459, L1460, L1473 ); 
   or4 U414 ( L1682, L1683, L1684, L1685, L1698 ); 
   or4 U415 ( L1686, L1687, L1688, L1689, L1701 ); 
   or4 U416 ( L1690, L1691, L1692, L1693, L1704 ); 
   or4 U417 ( L1694, L1695, L1696, L1697, L1707 ); 
   or4 U418 ( L1678, L1679, L1680, L1681, L2634 ); 
   buffer U419 ( L554, L319 ); 
   inv U420 ( L1500, L1504 ); 
   inv U421 ( L1509, L1513 ); 
   inv U422 ( L1521, L1524 ); 
   inv U423 ( L1525, L1528 ); 
   buffer U424 ( L1518, L1529 ); 
   buffer U425 ( L1518, L1533 ); 
   and3 U426 ( L1486, L1477, L1521, L1538 ); 
   and3 U427 ( L1490, L1481, L1525, L1541 ); 
   inv U428 ( L1777, L1781 ); 
   inv U429 ( L1786, L1790 ); 
   buffer U430 ( L1795, L1806 ); 
   buffer U431 ( L1795, L1810 ); 
   inv U432 ( L2730, L2734 ); 
   inv U433 ( L2515, L2521 ); 
   nand2 U434 ( L2515, L2522, L2524 ); 
   inv U435 ( L2525, L2531 ); 
   inv U436 ( L2528, L2532 ); 
   and2 U437 ( L838, L860, L144 ); 
   and2 U438 ( L846, L860, L147 ); 
   and2 U439 ( L841, L860, L152 ); 
   inv U440 ( L1464, L160 ); 
   inv U441 ( L1467, L162 ); 
   inv U442 ( L1461, L164 ); 
   inv U443 ( L1329, L166 ); 
   inv U444 ( L1327, L168 ); 
   inv U445 ( L857, L171 ); 
   and4 U446 ( L480, L483, L36, L554, L175 ); 
   and4 U447 ( L480, L483, L554, L547, L187 ); 
   buffer U448 ( L838, L516 ); 
   inv U449 ( L846, L852 ); 
   and2 U450 ( L841, L875, L885 ); 
   and2 U451 ( L846, L875, L887 ); 
   and2 U452 ( L1327, L868, L893 ); 
   inv U453 ( L838, L1028 ); 
   inv U454 ( L841, L1031 ); 
   inv U455 ( L846, L1035 ); 
   buffer U456 ( L854, L1041 ); 
   buffer U457 ( L857, L1049 ); 
   buffer U458 ( L1327, L1057 ); 
   buffer U459 ( L1329, L1060 ); 
   buffer U460 ( L1331, L1066 ); 
   buffer U461 ( L1333, L1072 ); 
   buffer U462 ( L1335, L1078 ); 
   nand2 U463 ( L2099, L1470, L1213 ); 
   nand2 U464 ( L2103, L1473, L1218 ); 
   buffer U465 ( L1704, L1250 ); 
   and2 U466 ( L1461, L1385, L1387 ); 
   inv U467 ( L1464, L1389 ); 
   and3 U468 ( L1481, L1486, L1524, L1537 ); 
   and3 U469 ( L1477, L1490, L1528, L1540 ); 
   and2 U470 ( L841, L1710, L1735 ); 
   and2 U471 ( L846, L1710, L1737 ); 
   and2 U472 ( L854, L1710, L1739 ); 
   and2 U473 ( L857, L1710, L1741 ); 
   and2 U474 ( L1327, L1721, L1743 ); 
   and2 U475 ( L1329, L1721, L1745 ); 
   and2 U476 ( L1331, L1721, L1747 ); 
   and2 U477 ( L1333, L1721, L1749 ); 
   and2 U478 ( L1335, L1721, L1751 ); 
   inv U479 ( L2634, L2638 ); 
   and2 U480 ( L1698, L2001, L2024 ); 
   and2 U481 ( L1701, L2001, L2026 ); 
   and2 U482 ( L1704, L2001, L2028 ); 
   and2 U483 ( L1707, L2001, L2030 ); 
   and2 U484 ( L1461, L2012, L2032 ); 
   and2 U485 ( L1464, L2012, L2034 ); 
   and2 U486 ( L1467, L2012, L2036 ); 
   and2 U487 ( L1470, L2012, L2038 ); 
   buffer U488 ( L841, L2154 ); 
   nand2 U489 ( L2518, L2521, L2523 ); 
   nand2 U490 ( L2528, L2531, L2533 ); 
   nand2 U491 ( L2525, L2532, L2534 ); 
   buffer U492 ( L1698, L2631 ); 
   buffer U493 ( L1704, L2639 ); 
   buffer U494 ( L1701, L2642 ); 
   buffer U495 ( L1461, L2647 ); 
   buffer U496 ( L1707, L2650 ); 
   buffer U497 ( L1467, L2655 ); 
   buffer U498 ( L1464, L2658 ); 
   buffer U499 ( L1473, L2665 ); 
   buffer U500 ( L1470, L2668 ); 
   or2 U501 ( L865, L152, L153 ); 
   inv U502 ( L175, L176 ); 
   inv U503 ( L187, L188 ); 
   buffer U504 ( L1041, L299 ); 
   buffer U505 ( L1049, L301 ); 
   buffer U506 ( L1057, L286 ); 
   buffer U507 ( L1060, L303 ); 
   buffer U508 ( L1066, L288 ); 
   buffer U509 ( L1072, L305 ); 
   buffer U510 ( L1078, L290 ); 
   inv U511 ( L1529, L1532 ); 
   inv U512 ( L1533, L1536 ); 
   nor2 U513 ( L1537, L1538, L1539 ); 
   nor2 U514 ( L1540, L1541, L1542 ); 
   and3 U515 ( L1509, L1500, L1529, L1544 ); 
   and3 U516 ( L1513, L1504, L1533, L1547 ); 
   or2 U517 ( L2037, L2038, L2065 ); 
   inv U518 ( L1806, L1809 ); 
   inv U519 ( L1810, L1813 ); 
   and3 U520 ( L1786, L1777, L1806, L1821 ); 
   and3 U521 ( L1790, L1781, L1810, L1824 ); 
   nand2 U522 ( L2523, L2524, L2538 ); 
   nand2 U523 ( L2533, L2534, L2546 ); 
   or2 U524 ( L1734, L1735, L2554 ); 
   or2 U525 ( L1736, L1737, L2562 ); 
   or2 U526 ( L1738, L1739, L2570 ); 
   or2 U527 ( L1740, L1741, L2578 ); 
   or2 U528 ( L1742, L1743, L2586 ); 
   or2 U529 ( L1744, L1745, L2594 ); 
   or2 U530 ( L1746, L1747, L2602 ); 
   or2 U531 ( L1748, L1749, L2610 ); 
   or2 U532 ( L1750, L1751, L2618 ); 
   or2 U533 ( L2023, L2024, L2626 ); 
   or2 U534 ( L2025, L2026, L2738 ); 
   or2 U535 ( L2027, L2028, L2746 ); 
   or2 U536 ( L2029, L2030, L2754 ); 
   or2 U537 ( L2031, L2032, L2762 ); 
   or2 U538 ( L2033, L2034, L2770 ); 
   or2 U539 ( L2035, L2036, L2778 ); 
   and3 U540 ( L1389, L1387, L40, L456 ); 
   inv U541 ( L1387, L466 ); 
   nand2 U542 ( L560, L852, L562 ); 
   and2 U543 ( L516, L875, L883 ); 
   and2 U544 ( L1049, L868, L889 ); 
   and2 U545 ( L1041, L875, L891 ); 
   inv U546 ( L1041, L1043 ); 
   inv U547 ( L1049, L1051 ); 
   inv U548 ( L1060, L1062 ); 
   inv U549 ( L1066, L1068 ); 
   inv U550 ( L1072, L1074 ); 
   inv U551 ( L1078, L1080 ); 
   and2 U552 ( L2099, L1213, L1225 ); 
   and2 U553 ( L1213, L1470, L1227 ); 
   and2 U554 ( L2103, L1218, L1232 ); 
   and2 U555 ( L1218, L1473, L1234 ); 
   and3 U556 ( L1504, L1509, L1532, L1543 ); 
   and3 U557 ( L1500, L1513, L1536, L1546 ); 
   inv U558 ( L2631, L2637 ); 
   nand2 U559 ( L2631, L2638, L1753 ); 
   inv U560 ( L2639, L2645 ); 
   inv U561 ( L2642, L2646 ); 
   inv U562 ( L2647, L2653 ); 
   inv U563 ( L2650, L2654 ); 
   and3 U564 ( L1781, L1786, L1809, L1820 ); 
   and3 U565 ( L1777, L1790, L1813, L1823 ); 
   buffer U566 ( L1031, L2107 ); 
   buffer U567 ( L1028, L2110 ); 
   buffer U568 ( L1035, L2118 ); 
   inv U569 ( L1057, L2123 ); 
   inv U570 ( L852, L2151 ); 
   inv U571 ( L2154, L2158 ); 
   buffer U572 ( L1031, L2161 ); 
   buffer U573 ( L1028, L2164 ); 
   buffer U574 ( L1035, L2172 ); 
   buffer U575 ( L516, L2235 ); 
   buffer U576 ( L1035, L2262 ); 
   buffer U577 ( L1035, L2350 ); 
   nand2 U578 ( L1542, L1539, L2535 ); 
   inv U579 ( L2655, L2661 ); 
   inv U580 ( L2658, L2662 ); 
   inv U581 ( L2665, L2671 ); 
   inv U582 ( L2668, L2672 ); 
   and3 U583 ( L40, L1389, L466, L468 ); 
   or2 U584 ( L887, L889, L897 ); 
   or2 U585 ( L891, L893, L898 ); 
   or2 U586 ( L1225, L1227, L1228 ); 
   or2 U587 ( L1232, L1234, L1235 ); 
   nor2 U588 ( L1543, L1544, L1545 ); 
   nor2 U589 ( L1546, L1547, L1548 ); 
   inv U590 ( L2538, L2542 ); 
   inv U591 ( L2546, L2550 ); 
   nand2 U592 ( L2554, L2557, L1561 ); 
   inv U593 ( L2554, L2558 ); 
   nand2 U594 ( L2562, L2565, L1565 ); 
   inv U595 ( L2562, L2566 ); 
   nand2 U596 ( L2570, L2573, L1569 ); 
   inv U597 ( L2570, L2574 ); 
   nand2 U598 ( L2578, L2581, L1573 ); 
   inv U599 ( L2578, L2582 ); 
   nand2 U600 ( L2586, L2589, L1577 ); 
   inv U601 ( L2586, L2590 ); 
   nand2 U602 ( L2594, L2597, L1581 ); 
   inv U603 ( L2594, L2598 ); 
   nand2 U604 ( L2602, L2605, L1585 ); 
   inv U605 ( L2602, L2606 ); 
   nand2 U606 ( L2610, L2613, L1589 ); 
   inv U607 ( L2610, L2614 ); 
   nand2 U608 ( L2618, L2621, L1593 ); 
   inv U609 ( L2618, L2622 ); 
   nand2 U610 ( L2626, L2629, L1597 ); 
   inv U611 ( L2626, L2630 ); 
   nand2 U612 ( L2634, L2637, L1752 ); 
   nand2 U613 ( L2642, L2645, L1761 ); 
   nand2 U614 ( L2639, L2646, L1762 ); 
   nand2 U615 ( L2650, L2653, L1770 ); 
   nand2 U616 ( L2647, L2654, L1771 ); 
   nor2 U617 ( L1820, L1821, L1822 ); 
   nor2 U618 ( L1823, L1824, L1825 ); 
   nand2 U619 ( L2738, L2741, L2039 ); 
   inv U620 ( L2738, L2742 ); 
   nand2 U621 ( L2746, L2749, L2043 ); 
   inv U622 ( L2746, L2750 ); 
   nand2 U623 ( L2754, L2757, L2047 ); 
   inv U624 ( L2754, L2758 ); 
   nand2 U625 ( L2762, L2765, L2051 ); 
   inv U626 ( L2762, L2766 ); 
   nand2 U627 ( L2770, L2773, L2055 ); 
   inv U628 ( L2770, L2774 ); 
   nand2 U629 ( L2778, L2781, L2059 ); 
   inv U630 ( L2778, L2782 ); 
   nand2 U631 ( L2658, L2661, L2663 ); 
   nand2 U632 ( L2655, L2662, L2664 ); 
   nand2 U633 ( L2668, L2671, L2673 ); 
   nand2 U634 ( L2665, L2672, L2674 ); 
   and2 U635 ( L562, L865, L146 ); 
   inv U636 ( L456, L462 ); 
   inv U637 ( L2107, L2113 ); 
   inv U638 ( L2110, L2114 ); 
   inv U639 ( L2118, L2122 ); 
   inv U640 ( L2123, L2129 ); 
   buffer U641 ( L562, L592 ); 
   inv U642 ( L2161, L2167 ); 
   inv U643 ( L2164, L2168 ); 
   inv U644 ( L2172, L2176 ); 
   inv U645 ( L2235, L2241 ); 
   inv U646 ( L2262, L2266 ); 
   inv U647 ( L456, L743 ); 
   buffer U648 ( L456, L749 ); 
   and2 U649 ( L562, L868, L886 ); 
   buffer U650 ( L897, L284 ); 
   buffer U651 ( L897, L321 ); 
   buffer U652 ( L898, L297 ); 
   buffer U653 ( L898, L280 ); 
   buffer U654 ( L456, L995 ); 
   inv U655 ( L456, L1006 ); 
   nand2 U656 ( L2535, L2542, L1550 ); 
   inv U657 ( L2350, L2354 ); 
   inv U658 ( L2535, L2541 ); 
   nand2 U659 ( L2551, L2558, L1562 ); 
   nand2 U660 ( L2559, L2566, L1566 ); 
   nand2 U661 ( L2567, L2574, L1570 ); 
   nand2 U662 ( L2575, L2582, L1574 ); 
   nand2 U663 ( L2583, L2590, L1578 ); 
   nand2 U664 ( L2591, L2598, L1582 ); 
   nand2 U665 ( L2599, L2606, L1586 ); 
   nand2 U666 ( L2607, L2614, L1590 ); 
   nand2 U667 ( L2615, L2622, L1594 ); 
   nand2 U668 ( L2623, L2630, L1598 ); 
   nand2 U669 ( L1752, L1753, L1754 ); 
   nand2 U670 ( L1761, L1762, L1763 ); 
   nand2 U671 ( L1770, L1771, L1772 ); 
   nand2 U672 ( L2735, L2742, L2040 ); 
   nand2 U673 ( L2743, L2750, L2044 ); 
   nand2 U674 ( L2751, L2758, L2048 ); 
   nand2 U675 ( L2759, L2766, L2052 ); 
   nand2 U676 ( L2767, L2774, L2056 ); 
   nand2 U677 ( L2775, L2782, L2060 ); 
   buffer U678 ( L1043, L2115 ); 
   buffer U679 ( L1051, L2126 ); 
   buffer U680 ( L1068, L2131 ); 
   buffer U681 ( L1062, L2134 ); 
   buffer U682 ( L1080, L2141 ); 
   buffer U683 ( L1074, L2144 ); 
   inv U684 ( L2151, L2157 ); 
   nand2 U685 ( L2151, L2158, L2160 ); 
   buffer U686 ( L1043, L2169 ); 
   buffer U687 ( L1068, L2177 ); 
   buffer U688 ( L1062, L2180 ); 
   buffer U689 ( L1080, L2187 ); 
   buffer U690 ( L1074, L2190 ); 
   inv U691 ( L562, L2207 ); 
   buffer U692 ( L1043, L2254 ); 
   buffer U693 ( L1051, L2334 ); 
   buffer U694 ( L1043, L2342 ); 
   buffer U695 ( L1051, L2422 ); 
   nand2 U696 ( L1548, L1545, L2543 ); 
   nand2 U697 ( L2673, L2674, L2709 ); 
   nand2 U698 ( L2663, L2664, L2712 ); 
   nand2 U699 ( L1825, L1822, L2727 ); 
   or2 U700 ( L146, L147, L148 ); 
   nand2 U701 ( L2110, L2113, L569 ); 
   nand2 U702 ( L2107, L2114, L570 ); 
   nand2 U703 ( L2164, L2167, L599 ); 
   nand2 U704 ( L2161, L2168, L600 ); 
   or2 U705 ( L885, L886, L896 ); 
   nand2 U706 ( L2538, L2541, L1549 ); 
   inv U707 ( L1228, L1243 ); 
   inv U708 ( L1235, L1245 ); 
   buffer U709 ( L468, L1257 ); 
   buffer U710 ( L468, L1258 ); 
   nand2 U711 ( L1561, L1562, L1563 ); 
   nand2 U712 ( L1565, L1566, L1567 ); 
   nand2 U713 ( L1569, L1570, L1571 ); 
   nand2 U714 ( L1573, L1574, L1575 ); 
   nand2 U715 ( L1577, L1578, L1579 ); 
   nand2 U716 ( L1581, L1582, L1583 ); 
   nand2 U717 ( L1585, L1586, L1587 ); 
   nand2 U718 ( L1589, L1590, L1591 ); 
   nand2 U719 ( L1593, L1594, L1595 ); 
   nand2 U720 ( L1597, L1598, L1599 ); 
   nand2 U721 ( L2039, L2040, L2041 ); 
   nand2 U722 ( L2043, L2044, L2045 ); 
   nand2 U723 ( L2047, L2048, L2049 ); 
   nand2 U724 ( L2051, L2052, L2053 ); 
   nand2 U725 ( L2055, L2056, L2057 ); 
   nand2 U726 ( L2059, L2060, L2061 ); 
   nand2 U727 ( L2154, L2157, L2159 ); 
   buffer U728 ( L462, L475 ); 
   and2 U729 ( L1078, L743, L490 ); 
   and2 U730 ( L1698, L743, L496 ); 
   and2 U731 ( L1701, L743, L502 ); 
   and2 U732 ( L1250, L743, L508 ); 
   and2 U733 ( L1057, L749, L765 ); 
   and2 U734 ( L1060, L749, L769 ); 
   nand2 U735 ( L569, L570, L571 ); 
   inv U736 ( L2115, L2121 ); 
   nand2 U737 ( L2115, L2122, L579 ); 
   nand2 U738 ( L2126, L2129, L587 ); 
   inv U739 ( L2126, L2130 ); 
   inv U740 ( L592, L596 ); 
   nand2 U741 ( L599, L600, L601 ); 
   inv U742 ( L2169, L2175 ); 
   nand2 U743 ( L2169, L2176, L609 ); 
   inv U744 ( L2254, L2258 ); 
   and2 U745 ( L1057, L995, L1014 ); 
   and2 U746 ( L1060, L995, L1018 ); 
   and2 U747 ( L1078, L1006, L717 ); 
   and2 U748 ( L1698, L1006, L723 ); 
   and2 U749 ( L1701, L1006, L729 ); 
   and2 U750 ( L1250, L1006, L735 ); 
   inv U751 ( L749, L753 ); 
   buffer U752 ( L896, L282 ); 
   buffer U753 ( L896, L323 ); 
   inv U754 ( L2334, L2338 ); 
   inv U755 ( L995, L999 ); 
   nand2 U756 ( L1549, L1550, L1091 ); 
   inv U757 ( L2342, L2346 ); 
   inv U758 ( L2422, L2426 ); 
   buffer U759 ( L462, L1337 ); 
   inv U760 ( L2543, L2549 ); 
   nand2 U761 ( L2543, L2550, L1552 ); 
   inv U762 ( L1599, L1600 ); 
   inv U763 ( L1595, L1596 ); 
   inv U764 ( L1591, L1592 ); 
   inv U765 ( L1587, L1588 ); 
   inv U766 ( L1583, L1584 ); 
   inv U767 ( L1579, L1580 ); 
   inv U768 ( L1575, L1576 ); 
   inv U769 ( L1571, L1572 ); 
   inv U770 ( L1567, L1568 ); 
   inv U771 ( L1563, L1564 ); 
   inv U772 ( L2061, L2062 ); 
   inv U773 ( L2057, L2058 ); 
   inv U774 ( L2053, L2054 ); 
   inv U775 ( L2049, L2050 ); 
   inv U776 ( L2045, L2046 ); 
   inv U777 ( L2041, L2042 ); 
   inv U778 ( L1754, L1758 ); 
   inv U779 ( L1763, L1767 ); 
   buffer U780 ( L1772, L1798 ); 
   buffer U781 ( L1772, L1802 ); 
   inv U782 ( L2727, L2733 ); 
   nand2 U783 ( L2727, L2734, L1829 ); 
   inv U784 ( L2131, L2137 ); 
   inv U785 ( L2134, L2138 ); 
   inv U786 ( L2141, L2147 ); 
   inv U787 ( L2144, L2148 ); 
   inv U788 ( L2177, L2183 ); 
   inv U789 ( L2180, L2184 ); 
   inv U790 ( L2187, L2193 ); 
   inv U791 ( L2190, L2194 ); 
   nand2 U792 ( L2159, L2160, L2210 ); 
   inv U793 ( L2207, L2213 ); 
   inv U794 ( L2709, L2715 ); 
   inv U795 ( L2712, L2716 ); 
   and2 U796 ( L1235, L1245, L1094 ); 
   and2 U797 ( L1228, L1243, L1096 ); 
   nand2 U798 ( L2118, L2121, L578 ); 
   nand2 U799 ( L2123, L2130, L588 ); 
   nand2 U800 ( L2172, L2175, L608 ); 
   buffer U801 ( L1257, L742 ); 
   buffer U802 ( L1257, L1005 ); 
   inv U803 ( L1091, L1092 ); 
   nand2 U804 ( L2546, L2549, L1551 ); 
   and5 U805 ( L1600, L1596, L1592, L1588, L1584, L1554 ); 
   and5 U806 ( L1580, L1576, L1572, L1568, L1564, L1555 ); 
   and2 U807 ( L2065, L2062, L1557 ); 
   and5 U808 ( L2058, L2054, L2050, L2046, L2042, L1558 ); 
   nand2 U809 ( L2730, L2733, L1828 ); 
   buffer U810 ( L1258, L1845 ); 
   buffer U811 ( L1258, L1907 ); 
   nand2 U812 ( L2134, L2137, L2139 ); 
   nand2 U813 ( L2131, L2138, L2140 ); 
   nand2 U814 ( L2144, L2147, L2149 ); 
   nand2 U815 ( L2141, L2148, L2150 ); 
   nand2 U816 ( L2180, L2183, L2185 ); 
   nand2 U817 ( L2177, L2184, L2186 ); 
   nand2 U818 ( L2190, L2193, L2195 ); 
   nand2 U819 ( L2187, L2194, L2196 ); 
   nand2 U820 ( L2712, L2715, L2717 ); 
   nand2 U821 ( L2709, L2716, L2718 ); 
   or2 U822 ( L1094, L1245, L154 ); 
   or2 U823 ( L1096, L1243, L155 ); 
   and2 U824 ( L1057, L753, L763 ); 
   and2 U825 ( L1060, L753, L767 ); 
   and2 U826 ( L1066, L753, L531 ); 
   and2 U827 ( L1072, L753, L537 ); 
   inv U828 ( L571, L575 ); 
   nand2 U829 ( L578, L579, L580 ); 
   nand2 U830 ( L587, L588, L589 ); 
   inv U831 ( L601, L605 ); 
   nand2 U832 ( L608, L609, L610 ); 
   and2 U833 ( L1057, L999, L1012 ); 
   and2 U834 ( L1060, L999, L1016 ); 
   and2 U835 ( L1066, L999, L705 ); 
   and2 U836 ( L1072, L999, L711 ); 
   and2 U837 ( L1092, L14, L1093 ); 
   buffer U838 ( L475, L1355 ); 
   nand2 U839 ( L1551, L1552, L1553 ); 
   and2 U840 ( L1554, L1555, L1556 ); 
   and2 U841 ( L1557, L1558, L1559 ); 
   buffer U842 ( L1337, L1601 ); 
   inv U843 ( L1798, L1801 ); 
   inv U844 ( L1802, L1805 ); 
   and3 U845 ( L1763, L1754, L1798, L1815 ); 
   and3 U846 ( L1767, L1758, L1802, L1818 ); 
   nand2 U847 ( L1828, L1829, L1830 ); 
   buffer U848 ( L475, L1836 ); 
   buffer U849 ( L475, L1850 ); 
   buffer U850 ( L1337, L1898 ); 
   buffer U851 ( L1337, L1912 ); 
   nand2 U852 ( L2149, L2150, L2197 ); 
   nand2 U853 ( L2139, L2140, L2200 ); 
   inv U854 ( L2210, L2214 ); 
   nand2 U855 ( L2210, L2213, L2215 ); 
   nand2 U856 ( L2195, L2196, L2217 ); 
   nand2 U857 ( L2185, L2186, L2220 ); 
   nand2 U858 ( L2717, L2718, L2722 ); 
   nand2 U859 ( L154, L155, L156 ); 
   and2 U860 ( L490, L742, L492 ); 
   and2 U861 ( L496, L742, L498 ); 
   and2 U862 ( L502, L742, L504 ); 
   and2 U863 ( L508, L742, L510 ); 
   or2 U864 ( L763, L765, L519 ); 
   or2 U865 ( L767, L769, L525 ); 
   and2 U866 ( L531, L748, L533 ); 
   and2 U867 ( L537, L748, L539 ); 
   or2 U868 ( L1012, L1014, L693 ); 
   or2 U869 ( L1016, L1018, L699 ); 
   and2 U870 ( L705, L994, L707 ); 
   and2 U871 ( L711, L994, L713 ); 
   and2 U872 ( L717, L1005, L719 ); 
   and2 U873 ( L723, L1005, L725 ); 
   and2 U874 ( L729, L1005, L731 ); 
   and2 U875 ( L735, L1005, L737 ); 
   buffer U876 ( L1093, L401 ); 
   and3 U877 ( L1556, L1559, L894, L1560 ); 
   and3 U878 ( L1758, L1763, L1801, L1814 ); 
   and3 U879 ( L1754, L1767, L1805, L1817 ); 
   nand2 U880 ( L2207, L2214, L2216 ); 
   inv U881 ( L1830, L227 ); 
   inv U882 ( L1553, L229 ); 
   inv U883 ( L492, L493 ); 
   inv U884 ( L498, L499 ); 
   inv U885 ( L504, L505 ); 
   inv U886 ( L510, L511 ); 
   and2 U887 ( L519, L748, L521 ); 
   and2 U888 ( L525, L748, L527 ); 
   inv U889 ( L533, L534 ); 
   inv U890 ( L539, L540 ); 
   inv U891 ( L580, L584 ); 
   buffer U892 ( L589, L613 ); 
   buffer U893 ( L589, L617 ); 
   buffer U894 ( L610, L621 ); 
   buffer U895 ( L610, L625 ); 
   and2 U896 ( L1344, L1355, L676 ); 
   and2 U897 ( L693, L994, L695 ); 
   and2 U898 ( L699, L994, L701 ); 
   inv U899 ( L707, L708 ); 
   inv U900 ( L713, L714 ); 
   inv U901 ( L719, L720 ); 
   inv U902 ( L725, L726 ); 
   inv U903 ( L731, L732 ); 
   inv U904 ( L737, L738 ); 
   inv U905 ( L1093, L1087 ); 
   and2 U906 ( L1344, L1601, L1108 ); 
   inv U907 ( L1355, L1361 ); 
   and2 U908 ( L1351, L1355, L1369 ); 
   and2 U909 ( L1959, L1355, L1373 ); 
   and2 U910 ( L1964, L1355, L1377 ); 
   buffer U911 ( L1560, L311 ); 
   inv U912 ( L1601, L1607 ); 
   and2 U913 ( L1351, L1601, L1615 ); 
   and2 U914 ( L1959, L1601, L1619 ); 
   and2 U915 ( L1964, L1601, L1623 ); 
   nor2 U916 ( L1814, L1815, L1816 ); 
   nor2 U917 ( L1817, L1818, L1819 ); 
   inv U918 ( L2722, L2726 ); 
   inv U919 ( L1836, L1842 ); 
   and2 U920 ( L1969, L1836, L1858 ); 
   and2 U921 ( L1974, L1836, L1863 ); 
   and2 U922 ( L1979, L1836, L1866 ); 
   and2 U923 ( L1984, L1836, L1868 ); 
   and2 U924 ( L1989, L1850, L1870 ); 
   and2 U925 ( L1994, L1850, L1872 ); 
   and2 U926 ( L1999, L1850, L1874 ); 
   and2 U927 ( L2070, L1850, L1876 ); 
   inv U928 ( L1898, L1904 ); 
   and2 U929 ( L1969, L1898, L1920 ); 
   and2 U930 ( L1974, L1898, L1925 ); 
   and2 U931 ( L1979, L1898, L1928 ); 
   and2 U932 ( L1984, L1898, L1930 ); 
   and2 U933 ( L1989, L1912, L1932 ); 
   and2 U934 ( L1994, L1912, L1934 ); 
   and2 U935 ( L1999, L1912, L1936 ); 
   and2 U936 ( L2070, L1912, L1938 ); 
   inv U937 ( L2197, L2203 ); 
   inv U938 ( L2200, L2204 ); 
   inv U939 ( L2217, L2223 ); 
   inv U940 ( L2220, L2224 ); 
   nand2 U941 ( L2215, L2216, L2238 ); 
   inv U942 ( L1560, L150 ); 
   inv U943 ( L521, L522 ); 
   inv U944 ( L527, L528 ); 
   inv U945 ( L695, L696 ); 
   inv U946 ( L701, L702 ); 
   and2 U947 ( L1866, L1831, L1881 ); 
   and2 U948 ( L1868, L1831, L1883 ); 
   and2 U949 ( L1870, L1845, L1885 ); 
   and2 U950 ( L1872, L1845, L1887 ); 
   and2 U951 ( L1874, L1845, L1889 ); 
   and2 U952 ( L1876, L1845, L1891 ); 
   and2 U953 ( L1928, L1893, L1943 ); 
   and2 U954 ( L1930, L1893, L1945 ); 
   and2 U955 ( L1932, L1907, L1947 ); 
   and2 U956 ( L1934, L1907, L1949 ); 
   and2 U957 ( L1936, L1907, L1951 ); 
   and2 U958 ( L1938, L1907, L1953 ); 
   nand2 U959 ( L2200, L2203, L2205 ); 
   nand2 U960 ( L2197, L2204, L2206 ); 
   nand2 U961 ( L2220, L2223, L2225 ); 
   nand2 U962 ( L2217, L2224, L2226 ); 
   nand2 U963 ( L1819, L1816, L2719 ); 
   inv U964 ( L613, L616 ); 
   inv U965 ( L617, L620 ); 
   inv U966 ( L621, L624 ); 
   inv U967 ( L625, L628 ); 
   and3 U968 ( L580, L571, L613, L630 ); 
   and3 U969 ( L584, L575, L617, L633 ); 
   and3 U970 ( L601, L592, L621, L636 ); 
   and3 U971 ( L605, L596, L625, L639 ); 
   nand2 U972 ( L2238, L2241, L645 ); 
   inv U973 ( L2238, L2242 ); 
   and2 U974 ( L1999, L1361, L675 ); 
   and2 U975 ( L1999, L1607, L1107 ); 
   and2 U976 ( L2070, L1361, L1368 ); 
   and2 U977 ( L2076, L1361, L1371 ); 
   and2 U978 ( L2082, L1361, L1375 ); 
   and2 U979 ( L2070, L1607, L1614 ); 
   and2 U980 ( L2076, L1607, L1617 ); 
   and2 U981 ( L2082, L1607, L1621 ); 
   and2 U982 ( L2088, L1842, L1856 ); 
   and2 U983 ( L2094, L1842, L1861 ); 
   and2 U984 ( L2088, L1904, L1918 ); 
   and2 U985 ( L2094, L1904, L1923 ); 
   nand2 U986 ( L2205, L2206, L2230 ); 
   nand2 U987 ( L2225, L2226, L2246 ); 
   buffer U988 ( L511, L2270 ); 
   buffer U989 ( L505, L2278 ); 
   buffer U990 ( L499, L2286 ); 
   buffer U991 ( L493, L2294 ); 
   buffer U992 ( L540, L2302 ); 
   buffer U993 ( L534, L2310 ); 
   buffer U994 ( L738, L2358 ); 
   buffer U995 ( L732, L2366 ); 
   buffer U996 ( L726, L2374 ); 
   buffer U997 ( L720, L2382 ); 
   buffer U998 ( L714, L2390 ); 
   buffer U999 ( L708, L2398 ); 
   and3 U1000 ( L575, L580, L616, L629 ); 
   and3 U1001 ( L571, L584, L620, L632 ); 
   and3 U1002 ( L596, L601, L624, L635 ); 
   and3 U1003 ( L592, L605, L628, L638 ); 
   nand2 U1004 ( L2235, L2242, L646 ); 
   or2 U1005 ( L675, L676, L677 ); 
   nand2 U1006 ( L2719, L2726, L1827 ); 
   and2 U1007 ( L1891, L511, L907 ); 
   and2 U1008 ( L1889, L505, L915 ); 
   and2 U1009 ( L1887, L499, L922 ); 
   and2 U1010 ( L493, L1885, L924 ); 
   and2 U1011 ( L1883, L540, L937 ); 
   and2 U1012 ( L1881, L534, L946 ); 
   or2 U1013 ( L1107, L1108, L1109 ); 
   and2 U1014 ( L1953, L738, L1125 ); 
   and2 U1015 ( L1951, L732, L1133 ); 
   and2 U1016 ( L1949, L726, L1140 ); 
   and2 U1017 ( L720, L1947, L1142 ); 
   and2 U1018 ( L1945, L714, L1155 ); 
   and2 U1019 ( L1943, L708, L1164 ); 
   or2 U1020 ( L1368, L1369, L1378 ); 
   or2 U1021 ( L1371, L1373, L1380 ); 
   or2 U1022 ( L1375, L1377, L1382 ); 
   or2 U1023 ( L1614, L1615, L1624 ); 
   or2 U1024 ( L1617, L1619, L1626 ); 
   or2 U1025 ( L1621, L1623, L1628 ); 
   inv U1026 ( L2719, L2725 ); 
   or2 U1027 ( L1856, L1858, L1859 ); 
   or2 U1028 ( L1861, L1863, L1864 ); 
   or2 U1029 ( L1918, L1920, L1921 ); 
   or2 U1030 ( L1923, L1925, L1926 ); 
   buffer U1031 ( L1891, L2267 ); 
   buffer U1032 ( L1889, L2275 ); 
   buffer U1033 ( L1887, L2283 ); 
   buffer U1034 ( L1885, L2291 ); 
   buffer U1035 ( L1883, L2299 ); 
   buffer U1036 ( L1881, L2307 ); 
   buffer U1037 ( L528, L2318 ); 
   buffer U1038 ( L522, L2326 ); 
   buffer U1039 ( L1953, L2355 ); 
   buffer U1040 ( L1951, L2363 ); 
   buffer U1041 ( L1949, L2371 ); 
   buffer U1042 ( L1947, L2379 ); 
   buffer U1043 ( L1945, L2387 ); 
   buffer U1044 ( L1943, L2395 ); 
   buffer U1045 ( L702, L2406 ); 
   buffer U1046 ( L696, L2414 ); 
   nand2 U1047 ( L645, L646, L647 ); 
   nor2 U1048 ( L629, L630, L631 ); 
   nor2 U1049 ( L632, L633, L634 ); 
   nor2 U1050 ( L635, L636, L637 ); 
   nor2 U1051 ( L638, L639, L640 ); 
   inv U1052 ( L2230, L2234 ); 
   inv U1053 ( L2246, L2250 ); 
   and2 U1054 ( L677, L1031, L679 ); 
   nand2 U1055 ( L2722, L2725, L1826 ); 
   inv U1056 ( L2270, L2274 ); 
   inv U1057 ( L2278, L2282 ); 
   inv U1058 ( L2286, L2290 ); 
   inv U1059 ( L2294, L2298 ); 
   inv U1060 ( L2302, L2306 ); 
   inv U1061 ( L2310, L2314 ); 
   and2 U1062 ( L1109, L1031, L1110 ); 
   inv U1063 ( L2358, L2362 ); 
   inv U1064 ( L2366, L2370 ); 
   inv U1065 ( L2374, L2378 ); 
   inv U1066 ( L2382, L2386 ); 
   inv U1067 ( L2390, L2394 ); 
   inv U1068 ( L2398, L2402 ); 
   and2 U1069 ( L1859, L1831, L1877 ); 
   and2 U1070 ( L1864, L1831, L1879 ); 
   and2 U1071 ( L1921, L1893, L1939 ); 
   and2 U1072 ( L1926, L1893, L1941 ); 
   and2 U1073 ( L647, L865, L143 ); 
   and2 U1074 ( L1380, L1043, L671 ); 
   and2 U1075 ( L1378, L1035, L674 ); 
   nand2 U1076 ( L1826, L1827, L686 ); 
   inv U1077 ( L2267, L2273 ); 
   nand2 U1078 ( L2267, L2274, L900 ); 
   inv U1079 ( L2275, L2281 ); 
   nand2 U1080 ( L2275, L2282, L909 ); 
   inv U1081 ( L2283, L2289 ); 
   nand2 U1082 ( L2283, L2290, L917 ); 
   inv U1083 ( L2291, L2297 ); 
   nand2 U1084 ( L2291, L2298, L926 ); 
   inv U1085 ( L2299, L2305 ); 
   nand2 U1086 ( L2299, L2306, L929 ); 
   inv U1087 ( L2307, L2313 ); 
   nand2 U1088 ( L2307, L2314, L939 ); 
   inv U1089 ( L2318, L2322 ); 
   inv U1090 ( L2326, L2330 ); 
   and2 U1091 ( L1382, L1051, L967 ); 
   and2 U1092 ( L1626, L1043, L1104 ); 
   and2 U1093 ( L1624, L1035, L1106 ); 
   inv U1094 ( L2355, L2361 ); 
   nand2 U1095 ( L2355, L2362, L1118 ); 
   inv U1096 ( L2363, L2369 ); 
   nand2 U1097 ( L2363, L2370, L1127 ); 
   inv U1098 ( L2371, L2377 ); 
   nand2 U1099 ( L2371, L2378, L1135 ); 
   inv U1100 ( L2379, L2385 ); 
   nand2 U1101 ( L2379, L2386, L1144 ); 
   inv U1102 ( L2387, L2393 ); 
   nand2 U1103 ( L2387, L2394, L1147 ); 
   inv U1104 ( L2395, L2401 ); 
   nand2 U1105 ( L2395, L2402, L1157 ); 
   inv U1106 ( L2406, L2410 ); 
   inv U1107 ( L2414, L2418 ); 
   and2 U1108 ( L1628, L1051, L1184 ); 
   nand2 U1109 ( L634, L631, L2227 ); 
   nand2 U1110 ( L640, L637, L2243 ); 
   buffer U1111 ( L1380, L2251 ); 
   buffer U1112 ( L1378, L2259 ); 
   buffer U1113 ( L1382, L2331 ); 
   buffer U1114 ( L1626, L2339 ); 
   buffer U1115 ( L1624, L2347 ); 
   buffer U1116 ( L1628, L2419 ); 
   or2 U1117 ( L143, L144, L145 ); 
   inv U1118 ( L686, L687 ); 
   nand2 U1119 ( L2270, L2273, L899 ); 
   nand2 U1120 ( L2278, L2281, L908 ); 
   nand2 U1121 ( L2286, L2289, L916 ); 
   nand2 U1122 ( L2294, L2297, L925 ); 
   nand2 U1123 ( L2302, L2305, L928 ); 
   nand2 U1124 ( L2310, L2313, L938 ); 
   and2 U1125 ( L1879, L528, L954 ); 
   and2 U1126 ( L1877, L522, L961 ); 
   nand2 U1127 ( L2358, L2361, L1117 ); 
   nand2 U1128 ( L2366, L2369, L1126 ); 
   nand2 U1129 ( L2374, L2377, L1134 ); 
   nand2 U1130 ( L2382, L2385, L1143 ); 
   nand2 U1131 ( L2390, L2393, L1146 ); 
   nand2 U1132 ( L2398, L2401, L1156 ); 
   and2 U1133 ( L1941, L702, L1172 ); 
   and2 U1134 ( L1939, L696, L1179 ); 
   buffer U1135 ( L1879, L2315 ); 
   buffer U1136 ( L1877, L2323 ); 
   buffer U1137 ( L1941, L2403 ); 
   buffer U1138 ( L1939, L2411 ); 
   inv U1139 ( L2227, L2233 ); 
   nand2 U1140 ( L2227, L2234, L642 ); 
   inv U1141 ( L2243, L2249 ); 
   nand2 U1142 ( L2243, L2250, L649 ); 
   inv U1143 ( L2251, L2257 ); 
   nand2 U1144 ( L2251, L2258, L665 ); 
   nand2 U1145 ( L2259, L2266, L684 ); 
   inv U1146 ( L2259, L2265 ); 
   and2 U1147 ( L687, L487, L688 ); 
   nand2 U1148 ( L899, L900, L901 ); 
   nand2 U1149 ( L908, L909, L910 ); 
   nand2 U1150 ( L916, L917, L918 ); 
   nand2 U1151 ( L925, L926, L927 ); 
   nand2 U1152 ( L928, L929, L930 ); 
   nand2 U1153 ( L938, L939, L940 ); 
   inv U1154 ( L2331, L2337 ); 
   nand2 U1155 ( L2331, L2338, L963 ); 
   inv U1156 ( L2339, L2345 ); 
   nand2 U1157 ( L2339, L2346, L1099 ); 
   nand2 U1158 ( L2347, L2354, L1115 ); 
   inv U1159 ( L2347, L2353 ); 
   nand2 U1160 ( L1117, L1118, L1119 ); 
   nand2 U1161 ( L1126, L1127, L1128 ); 
   nand2 U1162 ( L1134, L1135, L1136 ); 
   nand2 U1163 ( L1143, L1144, L1145 ); 
   nand2 U1164 ( L1146, L1147, L1148 ); 
   nand2 U1165 ( L1156, L1157, L1158 ); 
   inv U1166 ( L2419, L2425 ); 
   nand2 U1167 ( L2419, L2426, L1181 ); 
   nand2 U1168 ( L2230, L2233, L641 ); 
   nand2 U1169 ( L2246, L2249, L648 ); 
   nand2 U1170 ( L2254, L2257, L664 ); 
   nand2 U1171 ( L2262, L2265, L683 ); 
   buffer U1172 ( L688, L395 ); 
   inv U1173 ( L2315, L2321 ); 
   nand2 U1174 ( L2315, L2322, L948 ); 
   inv U1175 ( L2323, L2329 ); 
   nand2 U1176 ( L2323, L2330, L956 ); 
   nand2 U1177 ( L2334, L2337, L962 ); 
   nand2 U1178 ( L2342, L2345, L1098 ); 
   nand2 U1179 ( L2350, L2353, L1114 ); 
   inv U1180 ( L2403, L2409 ); 
   nand2 U1181 ( L2403, L2410, L1166 ); 
   inv U1182 ( L2411, L2417 ); 
   nand2 U1183 ( L2411, L2418, L1174 ); 
   nand2 U1184 ( L2422, L2425, L1180 ); 
   nand2 U1185 ( L641, L642, L643 ); 
   nand2 U1186 ( L648, L649, L650 ); 
   nand2 U1187 ( L664, L665, L666 ); 
   nand2 U1188 ( L683, L684, L681 ); 
   inv U1189 ( L688, L690 ); 
   nand2 U1190 ( L2318, L2321, L947 ); 
   nand2 U1191 ( L2326, L2329, L955 ); 
   nand2 U1192 ( L962, L963, L964 ); 
   and4 U1193 ( L910, L927, L918, L901, L968 ); 
   and2 U1194 ( L901, L915, L970 ); 
   and3 U1195 ( L910, L901, L922, L971 ); 
   and4 U1196 ( L918, L901, L924, L910, L972 ); 
   and2 U1197 ( L930, L946, L978 ); 
   and3 U1198 ( L940, L930, L954, L979 ); 
   nand2 U1199 ( L1098, L1099, L1100 ); 
   nand2 U1200 ( L1114, L1115, L1112 ); 
   nand2 U1201 ( L2406, L2409, L1165 ); 
   nand2 U1202 ( L2414, L2417, L1173 ); 
   nand2 U1203 ( L1180, L1181, L1182 ); 
   and4 U1204 ( L1128, L1145, L1136, L1119, L1185 ); 
   and2 U1205 ( L1119, L1133, L1187 ); 
   and3 U1206 ( L1128, L1119, L1140, L1188 ); 
   and4 U1207 ( L1136, L1119, L1142, L1128, L1189 ); 
   and2 U1208 ( L1148, L1164, L1195 ); 
   and3 U1209 ( L1158, L1148, L1172, L1196 ); 
   inv U1210 ( L643, L644 ); 
   and2 U1211 ( L650, L868, L884 ); 
   nand2 U1212 ( L947, L948, L949 ); 
   nand2 U1213 ( L955, L956, L957 ); 
   inv U1214 ( L968, L969 ); 
   or4 U1215 ( L907, L970, L971, L972, L973 ); 
   nand2 U1216 ( L1165, L1166, L1167 ); 
   nand2 U1217 ( L1173, L1174, L1175 ); 
   inv U1218 ( L1185, L1186 ); 
   or4 U1219 ( L1125, L1187, L1188, L1189, L1190 ); 
   and2 U1220 ( L666, L674, L680 ); 
   and3 U1221 ( L681, L666, L679, L682 ); 
   or2 U1222 ( L883, L884, L895 ); 
   and2 U1223 ( L644, L487, L1025 ); 
   and2 U1224 ( L1100, L1106, L1111 ); 
   and3 U1225 ( L1112, L1100, L1110, L1113 ); 
   or3 U1226 ( L671, L680, L682, L685 ); 
   buffer U1227 ( L895, L295 ); 
   buffer U1228 ( L895, L331 ); 
   inv U1229 ( L973, L976 ); 
   and5 U1230 ( L940, L964, L949, L930, L957, L977 ); 
   and4 U1231 ( L949, L930, L961, L940, L980 ); 
   and5 U1232 ( L957, L949, L930, L967, L940, L981 ); 
   buffer U1233 ( L1025, L397 ); 
   or3 U1234 ( L1104, L1111, L1113, L1116 ); 
   inv U1235 ( L1190, L1193 ); 
   and5 U1236 ( L1158, L1182, L1167, L1148, L1175, L1194 ); 
   and4 U1237 ( L1167, L1148, L1179, L1158, L1197 ); 
   and5 U1238 ( L1175, L1167, L1148, L1184, L1158, L1198 ); 
   or5 U1239 ( L937, L978, L979, L980, L981, L982 ); 
   and2 U1240 ( L977, L685, L983 ); 
   nand2 U1241 ( L976, L969, L988 ); 
   inv U1242 ( L1025, L1027 ); 
   or5 U1243 ( L1155, L1195, L1196, L1197, L1198, L1199 ); 
   and2 U1244 ( L1194, L1116, L1200 ); 
   nand2 U1245 ( L1193, L1186, L1205 ); 
   or2 U1246 ( L982, L983, L984 ); 
   and3 U1247 ( L690, L1027, L1830, L1085 ); 
   or2 U1248 ( L1199, L1200, L1201 ); 
   inv U1249 ( L984, L987 ); 
   and2 U1250 ( L988, L984, L990 ); 
   inv U1251 ( L1201, L1204 ); 
   and2 U1252 ( L1205, L1201, L1207 ); 
   and2 U1253 ( L973, L987, L989 ); 
   and2 U1254 ( L1190, L1204, L1206 ); 
   or2 U1255 ( L989, L990, L991 ); 
   or2 U1256 ( L1206, L1207, L1208 ); 
   buffer U1257 ( L1208, L329 ); 
   nand2 U1258 ( L1208, L991, L1221 ); 
   and2 U1259 ( L1208, L1221, L1238 ); 
   and2 U1260 ( L1221, L991, L1239 ); 
   or2 U1261 ( L1238, L1239, L1240 ); 
   inv U1262 ( L1240, L1247 ); 
   and2 U1263 ( L1240, L1247, L471 ); 
   or2 U1264 ( L471, L1247, L473 ); 
   inv U1265 ( L473, L231 ); 
   and3 U1266 ( L1553, L1087, L473, L1088 ); 
   and3 U1267 ( L1085, L1088, L554, L1089 ); 
   buffer U1268 ( L1089, L308 ); 
   inv U1269 ( L1089, L225 ); 
endmodule

