module top(G1 , G5 , G9 , G13 , G33 , G41 , G17 , G18 , G19 , G20 , G21 , G22 , G23 , G24 , G4 , G8 , G12 , G16 , G36 , G29 , G30 , G31 , G32 , G3 , G7 , G11 , G15 , G35 , G25 , G26 , G27 , G28 , G2 , G6 , G10 , G14 , G34 , G40 , G39 , G38 , G37 , G1324 , G1344 , G1325 , G1326 , G1327 , G1328 , G1329 , G1330 , G1343 , G1331 , G1332 , G1333 , G1334 , G1335 , G1336 , G1337 , G1338 , G1339 , G1340 , G1341 , G1342 , G1345 , G1346 , G1347 , G1348 , G1349 , G1350 , G1351 , G1352 , G1353 , G1354 , G1355 );
  input G1 , G5 , G9 , G13 , G33 , G41 , G17 , G18 , G19 , G20 , G21 , G22 , G23 , G24 , G4 , G8 , G12 , G16 , G36 , G29 , G30 , G31 , G32 , G3 , G7 , G11 , G15 , G35 , G25 , G26 , G27 , G28 , G2 , G6 , G10 , G14 , G34 , G40 , G39 , G38 , G37 ;
  output G1324 , G1344 , G1325 , G1326 , G1327 , G1328 , G1329 , G1330 , G1343 , G1331 , G1332 , G1333 , G1334 , G1335 , G1336 , G1337 , G1338 , G1339 , G1340 , G1341 , G1342 , G1345 , G1346 , G1347 , G1348 , G1349 , G1350 , G1351 , G1352 , G1353 , G1354 , G1355 ;
  wire n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543;
  assign n42 = G1 & G5 ;
  assign n43 = G1 & ~n42 ;
  assign n44 = G5 & ~n42 ;
  assign n45 = ~n43 & ~n44 ;
  assign n46 = G9 & G13 ;
  assign n47 = G9 & ~n46 ;
  assign n48 = G13 & ~n46 ;
  assign n49 = ~n47 & ~n48 ;
  assign n50 = ~n45 & ~n49 ;
  assign n51 = ~n45 & ~n50 ;
  assign n52 = ~n49 & ~n50 ;
  assign n53 = ~n51 & ~n52 ;
  assign n54 = G33 & G41 ;
  assign n55 = G17 & G18 ;
  assign n56 = G17 & ~n55 ;
  assign n57 = G18 & ~n55 ;
  assign n58 = ~n56 & ~n57 ;
  assign n59 = G19 & G20 ;
  assign n60 = G19 & ~n59 ;
  assign n61 = G20 & ~n59 ;
  assign n62 = ~n60 & ~n61 ;
  assign n63 = ~n58 & ~n62 ;
  assign n64 = ~n58 & ~n63 ;
  assign n65 = ~n62 & ~n63 ;
  assign n66 = ~n64 & ~n65 ;
  assign n67 = G21 & G22 ;
  assign n68 = G21 & ~n67 ;
  assign n69 = G22 & ~n67 ;
  assign n70 = ~n68 & ~n69 ;
  assign n71 = G23 & G24 ;
  assign n72 = G23 & ~n71 ;
  assign n73 = G24 & ~n71 ;
  assign n74 = ~n72 & ~n73 ;
  assign n75 = ~n70 & ~n74 ;
  assign n76 = ~n70 & ~n75 ;
  assign n77 = ~n74 & ~n75 ;
  assign n78 = ~n76 & ~n77 ;
  assign n79 = ~n66 & ~n78 ;
  assign n80 = ~n66 & ~n79 ;
  assign n81 = ~n78 & ~n79 ;
  assign n82 = ~n80 & ~n81 ;
  assign n83 = n54 & ~n82 ;
  assign n84 = n54 & ~n83 ;
  assign n85 = ~n82 & ~n83 ;
  assign n86 = ~n84 & ~n85 ;
  assign n87 = ~n53 & ~n86 ;
  assign n88 = ~n53 & ~n87 ;
  assign n89 = ~n86 & ~n87 ;
  assign n90 = ~n88 & ~n89 ;
  assign n91 = G4 & G8 ;
  assign n92 = G4 & ~n91 ;
  assign n93 = G8 & ~n91 ;
  assign n94 = ~n92 & ~n93 ;
  assign n95 = G12 & G16 ;
  assign n96 = G12 & ~n95 ;
  assign n97 = G16 & ~n95 ;
  assign n98 = ~n96 & ~n97 ;
  assign n99 = ~n94 & ~n98 ;
  assign n100 = ~n94 & ~n99 ;
  assign n101 = ~n98 & ~n99 ;
  assign n102 = ~n100 & ~n101 ;
  assign n103 = G41 & G36 ;
  assign n104 = G29 & G30 ;
  assign n105 = G29 & ~n104 ;
  assign n106 = G30 & ~n104 ;
  assign n107 = ~n105 & ~n106 ;
  assign n108 = G31 & G32 ;
  assign n109 = G31 & ~n108 ;
  assign n110 = G32 & ~n108 ;
  assign n111 = ~n109 & ~n110 ;
  assign n112 = ~n107 & ~n111 ;
  assign n113 = ~n107 & ~n112 ;
  assign n114 = ~n111 & ~n112 ;
  assign n115 = ~n113 & ~n114 ;
  assign n116 = ~n78 & ~n115 ;
  assign n117 = ~n78 & ~n116 ;
  assign n118 = ~n115 & ~n116 ;
  assign n119 = ~n117 & ~n118 ;
  assign n120 = n103 & ~n119 ;
  assign n121 = n103 & ~n120 ;
  assign n122 = ~n119 & ~n120 ;
  assign n123 = ~n121 & ~n122 ;
  assign n124 = ~n102 & ~n123 ;
  assign n125 = ~n102 & ~n124 ;
  assign n126 = ~n123 & ~n124 ;
  assign n127 = ~n125 & ~n126 ;
  assign n128 = G3 & G7 ;
  assign n129 = G3 & ~n128 ;
  assign n130 = G7 & ~n128 ;
  assign n131 = ~n129 & ~n130 ;
  assign n132 = G11 & G15 ;
  assign n133 = G11 & ~n132 ;
  assign n134 = G15 & ~n132 ;
  assign n135 = ~n133 & ~n134 ;
  assign n136 = ~n131 & ~n135 ;
  assign n137 = ~n131 & ~n136 ;
  assign n138 = ~n135 & ~n136 ;
  assign n139 = ~n137 & ~n138 ;
  assign n140 = G41 & G35 ;
  assign n141 = G25 & G26 ;
  assign n142 = G25 & ~n141 ;
  assign n143 = G26 & ~n141 ;
  assign n144 = ~n142 & ~n143 ;
  assign n145 = G27 & G28 ;
  assign n146 = G27 & ~n145 ;
  assign n147 = G28 & ~n145 ;
  assign n148 = ~n146 & ~n147 ;
  assign n149 = ~n144 & ~n148 ;
  assign n150 = ~n144 & ~n149 ;
  assign n151 = ~n148 & ~n149 ;
  assign n152 = ~n150 & ~n151 ;
  assign n153 = ~n66 & ~n152 ;
  assign n154 = ~n66 & ~n153 ;
  assign n155 = ~n152 & ~n153 ;
  assign n156 = ~n154 & ~n155 ;
  assign n157 = n140 & ~n156 ;
  assign n158 = n140 & ~n157 ;
  assign n159 = ~n156 & ~n157 ;
  assign n160 = ~n158 & ~n159 ;
  assign n161 = ~n139 & ~n160 ;
  assign n162 = ~n139 & ~n161 ;
  assign n163 = ~n160 & ~n161 ;
  assign n164 = ~n162 & ~n163 ;
  assign n165 = n127 & n164 ;
  assign n166 = G2 & G6 ;
  assign n167 = G2 & ~n166 ;
  assign n168 = G6 & ~n166 ;
  assign n169 = ~n167 & ~n168 ;
  assign n170 = G10 & G14 ;
  assign n171 = G10 & ~n170 ;
  assign n172 = G14 & ~n170 ;
  assign n173 = ~n171 & ~n172 ;
  assign n174 = ~n169 & ~n173 ;
  assign n175 = ~n169 & ~n174 ;
  assign n176 = ~n173 & ~n174 ;
  assign n177 = ~n175 & ~n176 ;
  assign n178 = G41 & G34 ;
  assign n179 = ~n115 & ~n152 ;
  assign n180 = ~n152 & ~n179 ;
  assign n181 = ~n115 & ~n179 ;
  assign n182 = ~n180 & ~n181 ;
  assign n183 = n178 & ~n182 ;
  assign n184 = n178 & ~n183 ;
  assign n185 = ~n182 & ~n183 ;
  assign n186 = ~n184 & ~n185 ;
  assign n187 = ~n177 & ~n186 ;
  assign n188 = ~n177 & ~n187 ;
  assign n189 = ~n186 & ~n187 ;
  assign n190 = ~n188 & ~n189 ;
  assign n191 = ~n90 & n190 ;
  assign n192 = n165 & n191 ;
  assign n193 = n90 & ~n190 ;
  assign n194 = n165 & n193 ;
  assign n195 = ~n192 & ~n194 ;
  assign n196 = n127 & ~n164 ;
  assign n197 = n90 & n190 ;
  assign n198 = n196 & n197 ;
  assign n199 = ~n127 & n164 ;
  assign n200 = n197 & n199 ;
  assign n201 = ~n198 & ~n200 ;
  assign n202 = n195 & n201 ;
  assign n203 = G20 & G24 ;
  assign n204 = G20 & ~n203 ;
  assign n205 = G24 & ~n203 ;
  assign n206 = ~n204 & ~n205 ;
  assign n207 = G32 & G28 ;
  assign n208 = G28 & ~n207 ;
  assign n209 = G32 & ~n207 ;
  assign n210 = ~n208 & ~n209 ;
  assign n211 = ~n206 & ~n210 ;
  assign n212 = ~n206 & ~n211 ;
  assign n213 = ~n210 & ~n211 ;
  assign n214 = ~n212 & ~n213 ;
  assign n215 = G41 & G40 ;
  assign n216 = G5 & G6 ;
  assign n217 = G5 & ~n216 ;
  assign n218 = G6 & ~n216 ;
  assign n219 = ~n217 & ~n218 ;
  assign n220 = G8 & G7 ;
  assign n221 = G7 & ~n220 ;
  assign n222 = G8 & ~n220 ;
  assign n223 = ~n221 & ~n222 ;
  assign n224 = ~n219 & ~n223 ;
  assign n225 = ~n219 & ~n224 ;
  assign n226 = ~n223 & ~n224 ;
  assign n227 = ~n225 & ~n226 ;
  assign n228 = G13 & G14 ;
  assign n229 = G13 & ~n228 ;
  assign n230 = G14 & ~n228 ;
  assign n231 = ~n229 & ~n230 ;
  assign n232 = G16 & G15 ;
  assign n233 = G15 & ~n232 ;
  assign n234 = G16 & ~n232 ;
  assign n235 = ~n233 & ~n234 ;
  assign n236 = ~n231 & ~n235 ;
  assign n237 = ~n231 & ~n236 ;
  assign n238 = ~n235 & ~n236 ;
  assign n239 = ~n237 & ~n238 ;
  assign n240 = ~n227 & ~n239 ;
  assign n241 = ~n227 & ~n240 ;
  assign n242 = ~n239 & ~n240 ;
  assign n243 = ~n241 & ~n242 ;
  assign n244 = n215 & ~n243 ;
  assign n245 = n215 & ~n244 ;
  assign n246 = ~n243 & ~n244 ;
  assign n247 = ~n245 & ~n246 ;
  assign n248 = ~n214 & ~n247 ;
  assign n249 = ~n214 & ~n248 ;
  assign n250 = ~n247 & ~n248 ;
  assign n251 = ~n249 & ~n250 ;
  assign n252 = ~n202 & n251 ;
  assign n253 = G19 & G23 ;
  assign n254 = G19 & ~n253 ;
  assign n255 = G23 & ~n253 ;
  assign n256 = ~n254 & ~n255 ;
  assign n257 = G31 & G27 ;
  assign n258 = G27 & ~n257 ;
  assign n259 = G31 & ~n257 ;
  assign n260 = ~n258 & ~n259 ;
  assign n261 = ~n256 & ~n260 ;
  assign n262 = ~n256 & ~n261 ;
  assign n263 = ~n260 & ~n261 ;
  assign n264 = ~n262 & ~n263 ;
  assign n265 = G41 & G39 ;
  assign n266 = G1 & G2 ;
  assign n267 = G1 & ~n266 ;
  assign n268 = G2 & ~n266 ;
  assign n269 = ~n267 & ~n268 ;
  assign n270 = G4 & G3 ;
  assign n271 = G3 & ~n270 ;
  assign n272 = G4 & ~n270 ;
  assign n273 = ~n271 & ~n272 ;
  assign n274 = ~n269 & ~n273 ;
  assign n275 = ~n269 & ~n274 ;
  assign n276 = ~n273 & ~n274 ;
  assign n277 = ~n275 & ~n276 ;
  assign n278 = G9 & G10 ;
  assign n279 = G9 & ~n278 ;
  assign n280 = G10 & ~n278 ;
  assign n281 = ~n279 & ~n280 ;
  assign n282 = G12 & G11 ;
  assign n283 = G11 & ~n282 ;
  assign n284 = G12 & ~n282 ;
  assign n285 = ~n283 & ~n284 ;
  assign n286 = ~n281 & ~n285 ;
  assign n287 = ~n281 & ~n286 ;
  assign n288 = ~n285 & ~n286 ;
  assign n289 = ~n287 & ~n288 ;
  assign n290 = ~n277 & ~n289 ;
  assign n291 = ~n277 & ~n290 ;
  assign n292 = ~n289 & ~n290 ;
  assign n293 = ~n291 & ~n292 ;
  assign n294 = n265 & ~n293 ;
  assign n295 = n265 & ~n294 ;
  assign n296 = ~n293 & ~n294 ;
  assign n297 = ~n295 & ~n296 ;
  assign n298 = ~n264 & ~n297 ;
  assign n299 = ~n264 & ~n298 ;
  assign n300 = ~n297 & ~n298 ;
  assign n301 = ~n299 & ~n300 ;
  assign n302 = G18 & G22 ;
  assign n303 = G18 & ~n302 ;
  assign n304 = G22 & ~n302 ;
  assign n305 = ~n303 & ~n304 ;
  assign n306 = G30 & G26 ;
  assign n307 = G26 & ~n306 ;
  assign n308 = G30 & ~n306 ;
  assign n309 = ~n307 & ~n308 ;
  assign n310 = ~n305 & ~n309 ;
  assign n311 = ~n305 & ~n310 ;
  assign n312 = ~n309 & ~n310 ;
  assign n313 = ~n311 & ~n312 ;
  assign n314 = G41 & G38 ;
  assign n315 = ~n239 & ~n289 ;
  assign n316 = ~n289 & ~n315 ;
  assign n317 = ~n239 & ~n315 ;
  assign n318 = ~n316 & ~n317 ;
  assign n319 = n314 & ~n318 ;
  assign n320 = n314 & ~n319 ;
  assign n321 = ~n318 & ~n319 ;
  assign n322 = ~n320 & ~n321 ;
  assign n323 = ~n313 & ~n322 ;
  assign n324 = ~n313 & ~n323 ;
  assign n325 = ~n322 & ~n323 ;
  assign n326 = ~n324 & ~n325 ;
  assign n327 = G17 & G21 ;
  assign n328 = G17 & ~n327 ;
  assign n329 = G21 & ~n327 ;
  assign n330 = ~n328 & ~n329 ;
  assign n331 = G29 & G25 ;
  assign n332 = G25 & ~n331 ;
  assign n333 = G29 & ~n331 ;
  assign n334 = ~n332 & ~n333 ;
  assign n335 = ~n330 & ~n334 ;
  assign n336 = ~n330 & ~n335 ;
  assign n337 = ~n334 & ~n335 ;
  assign n338 = ~n336 & ~n337 ;
  assign n339 = G41 & G37 ;
  assign n340 = ~n227 & ~n277 ;
  assign n341 = ~n277 & ~n340 ;
  assign n342 = ~n227 & ~n340 ;
  assign n343 = ~n341 & ~n342 ;
  assign n344 = n339 & ~n343 ;
  assign n345 = n339 & ~n344 ;
  assign n346 = ~n343 & ~n344 ;
  assign n347 = ~n345 & ~n346 ;
  assign n348 = ~n338 & ~n347 ;
  assign n349 = ~n338 & ~n348 ;
  assign n350 = ~n347 & ~n348 ;
  assign n351 = ~n349 & ~n350 ;
  assign n352 = n326 & ~n351 ;
  assign n353 = ~n301 & n352 ;
  assign n354 = n252 & n353 ;
  assign n355 = ~n90 & n354 ;
  assign n356 = G1 & n355 ;
  assign n357 = G1 & ~n356 ;
  assign n358 = n355 & ~n356 ;
  assign n359 = ~n357 & ~n358 ;
  assign n360 = n251 & n301 ;
  assign n361 = n352 & n360 ;
  assign n362 = ~n326 & n351 ;
  assign n363 = n360 & n362 ;
  assign n364 = ~n361 & ~n363 ;
  assign n365 = n251 & ~n301 ;
  assign n366 = n326 & n351 ;
  assign n367 = n365 & n366 ;
  assign n368 = ~n251 & n301 ;
  assign n369 = n366 & n368 ;
  assign n370 = ~n367 & ~n369 ;
  assign n371 = n364 & n370 ;
  assign n372 = ~n127 & ~n371 ;
  assign n373 = n164 & n191 ;
  assign n374 = n372 & n373 ;
  assign n375 = ~n351 & n374 ;
  assign n376 = G21 & n375 ;
  assign n377 = G21 & ~n376 ;
  assign n378 = n375 & ~n376 ;
  assign n379 = ~n377 & ~n378 ;
  assign n380 = ~n190 & n354 ;
  assign n381 = G2 & n380 ;
  assign n382 = G2 & ~n381 ;
  assign n383 = n380 & ~n381 ;
  assign n384 = ~n382 & ~n383 ;
  assign n385 = ~n164 & n354 ;
  assign n386 = G3 & n385 ;
  assign n387 = G3 & ~n386 ;
  assign n388 = n385 & ~n386 ;
  assign n389 = ~n387 & ~n388 ;
  assign n390 = ~n127 & n354 ;
  assign n391 = G4 & n390 ;
  assign n392 = G4 & ~n391 ;
  assign n393 = n390 & ~n391 ;
  assign n394 = ~n392 & ~n393 ;
  assign n395 = ~n202 & ~n251 ;
  assign n396 = n301 & n352 ;
  assign n397 = n395 & n396 ;
  assign n398 = ~n90 & n397 ;
  assign n399 = G5 & n398 ;
  assign n400 = G5 & ~n399 ;
  assign n401 = n398 & ~n399 ;
  assign n402 = ~n400 & ~n401 ;
  assign n403 = ~n190 & n397 ;
  assign n404 = G6 & n403 ;
  assign n405 = G6 & ~n404 ;
  assign n406 = n403 & ~n404 ;
  assign n407 = ~n405 & ~n406 ;
  assign n408 = ~n164 & n397 ;
  assign n409 = G7 & n408 ;
  assign n410 = G7 & ~n409 ;
  assign n411 = n408 & ~n409 ;
  assign n412 = ~n410 & ~n411 ;
  assign n413 = n127 & ~n371 ;
  assign n414 = ~n164 & n191 ;
  assign n415 = n413 & n414 ;
  assign n416 = ~n251 & n415 ;
  assign n417 = G20 & n416 ;
  assign n418 = G20 & ~n417 ;
  assign n419 = n416 & ~n417 ;
  assign n420 = ~n418 & ~n419 ;
  assign n421 = ~n127 & n397 ;
  assign n422 = G8 & n421 ;
  assign n423 = G8 & ~n422 ;
  assign n424 = n421 & ~n422 ;
  assign n425 = ~n423 & ~n424 ;
  assign n426 = ~n301 & n362 ;
  assign n427 = n252 & n426 ;
  assign n428 = ~n90 & n427 ;
  assign n429 = G9 & n428 ;
  assign n430 = G9 & ~n429 ;
  assign n431 = n428 & ~n429 ;
  assign n432 = ~n430 & ~n431 ;
  assign n433 = ~n190 & n427 ;
  assign n434 = G10 & n433 ;
  assign n435 = G10 & ~n434 ;
  assign n436 = n433 & ~n434 ;
  assign n437 = ~n435 & ~n436 ;
  assign n438 = ~n164 & n427 ;
  assign n439 = G11 & n438 ;
  assign n440 = G11 & ~n439 ;
  assign n441 = n438 & ~n439 ;
  assign n442 = ~n440 & ~n441 ;
  assign n443 = ~n127 & n427 ;
  assign n444 = G12 & n443 ;
  assign n445 = G12 & ~n444 ;
  assign n446 = n443 & ~n444 ;
  assign n447 = ~n445 & ~n446 ;
  assign n448 = n301 & n362 ;
  assign n449 = n395 & n448 ;
  assign n450 = ~n90 & n449 ;
  assign n451 = G13 & n450 ;
  assign n452 = G13 & ~n451 ;
  assign n453 = n450 & ~n451 ;
  assign n454 = ~n452 & ~n453 ;
  assign n455 = ~n190 & n449 ;
  assign n456 = G14 & n455 ;
  assign n457 = G14 & ~n456 ;
  assign n458 = n455 & ~n456 ;
  assign n459 = ~n457 & ~n458 ;
  assign n460 = ~n164 & n449 ;
  assign n461 = G15 & n460 ;
  assign n462 = G15 & ~n461 ;
  assign n463 = n460 & ~n461 ;
  assign n464 = ~n462 & ~n463 ;
  assign n465 = ~n127 & n449 ;
  assign n466 = G16 & n465 ;
  assign n467 = G16 & ~n466 ;
  assign n468 = n465 & ~n466 ;
  assign n469 = ~n467 & ~n468 ;
  assign n470 = ~n351 & n415 ;
  assign n471 = G17 & n470 ;
  assign n472 = G17 & ~n471 ;
  assign n473 = n470 & ~n471 ;
  assign n474 = ~n472 & ~n473 ;
  assign n475 = ~n326 & n415 ;
  assign n476 = G18 & n475 ;
  assign n477 = G18 & ~n476 ;
  assign n478 = n475 & ~n476 ;
  assign n479 = ~n477 & ~n478 ;
  assign n480 = ~n301 & n415 ;
  assign n481 = G19 & n480 ;
  assign n482 = G19 & ~n481 ;
  assign n483 = n480 & ~n481 ;
  assign n484 = ~n482 & ~n483 ;
  assign n485 = ~n326 & n374 ;
  assign n486 = G22 & n485 ;
  assign n487 = G22 & ~n486 ;
  assign n488 = n485 & ~n486 ;
  assign n489 = ~n487 & ~n488 ;
  assign n490 = ~n301 & n374 ;
  assign n491 = G23 & n490 ;
  assign n492 = G23 & ~n491 ;
  assign n493 = n490 & ~n491 ;
  assign n494 = ~n492 & ~n493 ;
  assign n495 = ~n251 & n374 ;
  assign n496 = G24 & n495 ;
  assign n497 = G24 & ~n496 ;
  assign n498 = n495 & ~n496 ;
  assign n499 = ~n497 & ~n498 ;
  assign n500 = ~n164 & n193 ;
  assign n501 = n413 & n500 ;
  assign n502 = ~n351 & n501 ;
  assign n503 = G25 & n502 ;
  assign n504 = G25 & ~n503 ;
  assign n505 = n502 & ~n503 ;
  assign n506 = ~n504 & ~n505 ;
  assign n507 = ~n326 & n501 ;
  assign n508 = G26 & n507 ;
  assign n509 = G26 & ~n508 ;
  assign n510 = n507 & ~n508 ;
  assign n511 = ~n509 & ~n510 ;
  assign n512 = ~n301 & n501 ;
  assign n513 = G27 & n512 ;
  assign n514 = G27 & ~n513 ;
  assign n515 = n512 & ~n513 ;
  assign n516 = ~n514 & ~n515 ;
  assign n517 = ~n251 & n501 ;
  assign n518 = G28 & n517 ;
  assign n519 = G28 & ~n518 ;
  assign n520 = n517 & ~n518 ;
  assign n521 = ~n519 & ~n520 ;
  assign n522 = n164 & n193 ;
  assign n523 = n372 & n522 ;
  assign n524 = ~n351 & n523 ;
  assign n525 = G29 & n524 ;
  assign n526 = G29 & ~n525 ;
  assign n527 = n524 & ~n525 ;
  assign n528 = ~n526 & ~n527 ;
  assign n529 = ~n326 & n523 ;
  assign n530 = G30 & n529 ;
  assign n531 = G30 & ~n530 ;
  assign n532 = n529 & ~n530 ;
  assign n533 = ~n531 & ~n532 ;
  assign n534 = ~n301 & n523 ;
  assign n535 = G31 & n534 ;
  assign n536 = G31 & ~n535 ;
  assign n537 = n534 & ~n535 ;
  assign n538 = ~n536 & ~n537 ;
  assign n539 = ~n251 & n523 ;
  assign n540 = G32 & n539 ;
  assign n541 = G32 & ~n540 ;
  assign n542 = n539 & ~n540 ;
  assign n543 = ~n541 & ~n542 ;
  assign G1324 = n359 ;
  assign G1344 = n379 ;
  assign G1325 = n384 ;
  assign G1326 = n389 ;
  assign G1327 = n394 ;
  assign G1328 = n402 ;
  assign G1329 = n407 ;
  assign G1330 = n412 ;
  assign G1343 = n420 ;
  assign G1331 = n425 ;
  assign G1332 = n432 ;
  assign G1333 = n437 ;
  assign G1334 = n442 ;
  assign G1335 = n447 ;
  assign G1336 = n454 ;
  assign G1337 = n459 ;
  assign G1338 = n464 ;
  assign G1339 = n469 ;
  assign G1340 = n474 ;
  assign G1341 = n479 ;
  assign G1342 = n484 ;
  assign G1345 = n489 ;
  assign G1346 = n494 ;
  assign G1347 = n499 ;
  assign G1348 = n506 ;
  assign G1349 = n511 ;
  assign G1350 = n516 ;
  assign G1351 = n521 ;
  assign G1352 = n528 ;
  assign G1353 = n533 ;
  assign G1354 = n538 ;
  assign G1355 = n543 ;
endmodule
