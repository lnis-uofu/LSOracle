module top(pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 , pi8 , pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 , pi16 , pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 , po0 , po1 , po2 , po3 , po4 , po5 , po6 , po7 , po8 , po9 , po10 , po11 , po12 , po13 , po14 , po15 , po16 , po17 , po18 , po19 , po20 , po21 , po22 , po23 , po24 );
  input pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 , pi8 , pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 , pi16 , pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 ;
  output po0 , po1 , po2 , po3 , po4 , po5 , po6 , po7 , po8 , po9 , po10 , po11 , po12 , po13 , po14 , po15 , po16 , po17 , po18 , po19 , po20 , po21 , po22 , po23 , po24 ;
  wire n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743;
  assign n25 = pi2 & pi22 ;
  assign n26 = pi0 & ~pi22 ;
  assign n27 = pi1 | pi2 ;
  assign n28 = ( ~pi22 & n26 ) | ( ~pi22 & n27 ) | ( n26 & n27 );
  assign n29 = pi0 | pi1 ;
  assign n30 = pi2 & n29 ;
  assign n31 = n28 & ~n30 ;
  assign n32 = n25 | n31 ;
  assign n33 = pi10 | pi11 ;
  assign n34 = pi12 | pi13 ;
  assign n35 = n33 | n34 ;
  assign n36 = pi14 | n35 ;
  assign n37 = pi0 | n27 ;
  assign n38 = pi3 | n37 ;
  assign n39 = pi4 | n38 ;
  assign n40 = pi5 | pi6 ;
  assign n41 = n39 | n40 ;
  assign n42 = pi7 | pi8 ;
  assign n43 = pi9 | n42 ;
  assign n44 = n41 | n43 ;
  assign n45 = n36 | n44 ;
  assign n46 = pi15 | n45 ;
  assign n47 = pi16 | pi17 ;
  assign n48 = n46 | n47 ;
  assign n49 = pi18 | pi19 ;
  assign n50 = pi20 | n49 ;
  assign n51 = n48 | n50 ;
  assign n52 = ~pi22 & n51 ;
  assign n53 = pi21 | pi22 ;
  assign n54 = n51 & ~n53 ;
  assign n55 = ~pi21 & pi22 ;
  assign n56 = ( pi21 & n51 ) | ( pi21 & ~n55 ) | ( n51 & ~n55 );
  assign n57 = ( ~n52 & n54 ) | ( ~n52 & n56 ) | ( n54 & n56 );
  assign n58 = ~pi22 & n45 ;
  assign n59 = ~pi15 & n58 ;
  assign n60 = pi15 | n58 ;
  assign n61 = ( ~n58 & n59 ) | ( ~n58 & n60 ) | ( n59 & n60 );
  assign n62 = ( ~pi22 & n48 ) | ( ~pi22 & n49 ) | ( n48 & n49 );
  assign n63 = ( pi20 & pi22 ) | ( pi20 & n49 ) | ( pi22 & n49 );
  assign n64 = ( pi20 & n48 ) | ( pi20 & n63 ) | ( n48 & n63 );
  assign n65 = n62 & ~n64 ;
  assign n66 = ~pi22 & n64 ;
  assign n67 = ( pi20 & n65 ) | ( pi20 & ~n66 ) | ( n65 & ~n66 );
  assign n68 = n61 & ~n67 ;
  assign n69 = ~n57 & n68 ;
  assign n70 = pi16 & ~pi22 ;
  assign n71 = ( ~pi22 & n46 ) | ( ~pi22 & n70 ) | ( n46 & n70 );
  assign n72 = pi17 & ~n71 ;
  assign n73 = ~pi17 & n71 ;
  assign n74 = n72 | n73 ;
  assign n75 = ~pi22 & n46 ;
  assign n76 = pi16 | pi22 ;
  assign n77 = n46 & ~n76 ;
  assign n78 = pi16 | n77 ;
  assign n79 = ( ~n75 & n77 ) | ( ~n75 & n78 ) | ( n77 & n78 );
  assign n80 = n74 & n79 ;
  assign n81 = pi18 & ~pi22 ;
  assign n82 = ( ~pi22 & n48 ) | ( ~pi22 & n81 ) | ( n48 & n81 );
  assign n83 = pi19 & n81 ;
  assign n84 = pi19 & ~pi22 ;
  assign n85 = ( n48 & n83 ) | ( n48 & n84 ) | ( n83 & n84 );
  assign n86 = pi19 & ~n85 ;
  assign n87 = ( n82 & ~n85 ) | ( n82 & n86 ) | ( ~n85 & n86 );
  assign n88 = ~pi22 & n48 ;
  assign n89 = pi18 | pi22 ;
  assign n90 = n48 & ~n89 ;
  assign n91 = ~pi18 & n89 ;
  assign n92 = ( pi18 & n48 ) | ( pi18 & ~n91 ) | ( n48 & ~n91 );
  assign n93 = ( ~n88 & n90 ) | ( ~n88 & n92 ) | ( n90 & n92 );
  assign n94 = n87 | n93 ;
  assign n95 = n80 & ~n94 ;
  assign n96 = n69 & n95 ;
  assign n97 = n61 | n67 ;
  assign n98 = n57 | n97 ;
  assign n99 = ~n74 & n79 ;
  assign n100 = ~n94 & n99 ;
  assign n101 = ~n98 & n100 ;
  assign n102 = ~n57 & n67 ;
  assign n103 = n61 & n102 ;
  assign n104 = n87 & n93 ;
  assign n105 = n80 & n104 ;
  assign n106 = n103 & n105 ;
  assign n107 = n74 | n79 ;
  assign n108 = n104 & ~n107 ;
  assign n109 = n103 & n108 ;
  assign n110 = ~n87 & n93 ;
  assign n111 = n80 & n110 ;
  assign n112 = n103 & n111 ;
  assign n113 = n74 & ~n79 ;
  assign n114 = n110 & n113 ;
  assign n115 = n103 & n114 ;
  assign n116 = ~n61 & n67 ;
  assign n117 = ~n57 & n116 ;
  assign n118 = n87 & ~n93 ;
  assign n119 = n80 & n118 ;
  assign n120 = n117 & n119 ;
  assign n121 = n115 | n120 ;
  assign n122 = ~n94 & n113 ;
  assign n123 = n69 & n122 ;
  assign n124 = n108 & n117 ;
  assign n125 = n99 & n110 ;
  assign n126 = n117 & n125 ;
  assign n127 = n103 & n119 ;
  assign n128 = n57 & ~n97 ;
  assign n129 = n100 & n128 ;
  assign n130 = n99 & n104 ;
  assign n131 = n117 & n130 ;
  assign n132 = n57 & n68 ;
  assign n133 = n94 | n107 ;
  assign n134 = n132 & ~n133 ;
  assign n135 = n131 | n134 ;
  assign n136 = n129 | n135 ;
  assign n137 = n127 | n136 ;
  assign n138 = n126 | n137 ;
  assign n139 = n124 | n138 ;
  assign n140 = n123 | n139 ;
  assign n141 = n98 | n133 ;
  assign n142 = n100 & n132 ;
  assign n143 = n95 & ~n98 ;
  assign n144 = n142 | n143 ;
  assign n145 = n141 & ~n144 ;
  assign n146 = ~n98 & n105 ;
  assign n147 = n104 & n113 ;
  assign n148 = ~n98 & n147 ;
  assign n149 = ~n107 & n110 ;
  assign n150 = n128 & n149 ;
  assign n151 = n125 & n128 ;
  assign n152 = n150 | n151 ;
  assign n153 = n69 & n147 ;
  assign n154 = n117 & ~n133 ;
  assign n155 = n153 | n154 ;
  assign n156 = n103 & ~n133 ;
  assign n157 = n132 & n149 ;
  assign n158 = n125 & n132 ;
  assign n159 = n157 | n158 ;
  assign n160 = n156 | n159 ;
  assign n161 = n69 & n108 ;
  assign n162 = n69 & n130 ;
  assign n163 = n161 | n162 ;
  assign n164 = n160 | n163 ;
  assign n165 = n155 | n164 ;
  assign n166 = n152 | n165 ;
  assign n167 = n148 | n166 ;
  assign n168 = n146 | n167 ;
  assign n169 = n69 & n105 ;
  assign n170 = ~n98 & n130 ;
  assign n171 = n169 | n170 ;
  assign n172 = n168 | n171 ;
  assign n173 = n145 & ~n172 ;
  assign n174 = n99 & n118 ;
  assign n175 = n57 & n67 ;
  assign n176 = n61 & n175 ;
  assign n177 = n174 & n176 ;
  assign n178 = n113 & n118 ;
  assign n179 = ~n61 & n175 ;
  assign n180 = n178 & n179 ;
  assign n181 = n119 & n179 ;
  assign n182 = n180 | n181 ;
  assign n183 = n176 & n178 ;
  assign n184 = n108 & n132 ;
  assign n185 = n95 & n179 ;
  assign n186 = n184 | n185 ;
  assign n187 = n183 | n186 ;
  assign n188 = n182 | n187 ;
  assign n189 = n128 & n130 ;
  assign n190 = n95 & n176 ;
  assign n191 = n130 & n132 ;
  assign n192 = n190 | n191 ;
  assign n193 = n189 | n192 ;
  assign n194 = n188 | n193 ;
  assign n195 = n132 & n174 ;
  assign n196 = n149 & n176 ;
  assign n197 = ~n107 & n118 ;
  assign n198 = n132 & n197 ;
  assign n199 = n111 & n176 ;
  assign n200 = n128 & n197 ;
  assign n201 = n199 | n200 ;
  assign n202 = n198 | n201 ;
  assign n203 = n128 & n174 ;
  assign n204 = n114 & n176 ;
  assign n205 = n111 & n179 ;
  assign n206 = n149 & n179 ;
  assign n207 = n205 | n206 ;
  assign n208 = n204 | n207 ;
  assign n209 = n203 | n208 ;
  assign n210 = n202 | n209 ;
  assign n211 = n196 | n210 ;
  assign n212 = n195 | n211 ;
  assign n213 = n108 & n128 ;
  assign n214 = n105 & n132 ;
  assign n215 = ~n133 & n179 ;
  assign n216 = n214 | n215 ;
  assign n217 = n213 | n216 ;
  assign n218 = n212 | n217 ;
  assign n219 = n194 | n218 ;
  assign n220 = ~n133 & n176 ;
  assign n221 = n130 & n179 ;
  assign n222 = n100 & n179 ;
  assign n223 = n221 | n222 ;
  assign n224 = n147 & n179 ;
  assign n225 = n130 & n176 ;
  assign n226 = n224 | n225 ;
  assign n227 = n223 | n226 ;
  assign n228 = n220 | n227 ;
  assign n229 = n219 | n228 ;
  assign n230 = n177 | n229 ;
  assign n231 = n173 & ~n230 ;
  assign n232 = ~n140 & n231 ;
  assign n233 = n128 & ~n133 ;
  assign n234 = n114 & n117 ;
  assign n235 = n111 & n117 ;
  assign n236 = n103 & n125 ;
  assign n237 = n235 | n236 ;
  assign n238 = n234 | n237 ;
  assign n239 = n233 | n238 ;
  assign n240 = n69 & n100 ;
  assign n241 = n69 & ~n133 ;
  assign n242 = n240 | n241 ;
  assign n243 = n239 | n242 ;
  assign n244 = n232 & ~n243 ;
  assign n245 = ~n98 & n122 ;
  assign n246 = ~n98 & n149 ;
  assign n247 = n245 | n246 ;
  assign n248 = n244 & ~n247 ;
  assign n249 = ~n121 & n248 ;
  assign n250 = ~n112 & n249 ;
  assign n251 = ~n109 & n250 ;
  assign n252 = ~n106 & n251 ;
  assign n253 = ~n101 & n252 ;
  assign n254 = ~n96 & n253 ;
  assign n255 = ( pi10 & ~pi22 ) | ( pi10 & n44 ) | ( ~pi22 & n44 );
  assign n256 = ( pi10 & ~pi11 ) | ( pi10 & pi22 ) | ( ~pi11 & pi22 );
  assign n257 = ( ~pi11 & n44 ) | ( ~pi11 & n256 ) | ( n44 & n256 );
  assign n258 = n255 & ~n257 ;
  assign n311 = n69 & n174 ;
  assign n312 = ~n98 & n174 ;
  assign n313 = ~n98 & n178 ;
  assign n314 = n120 | n127 ;
  assign n315 = n103 & n147 ;
  assign n316 = n103 & n130 ;
  assign n317 = n109 | n316 ;
  assign n318 = n131 | n317 ;
  assign n319 = n315 | n318 ;
  assign n320 = n314 | n319 ;
  assign n321 = n117 & n147 ;
  assign n322 = n103 & n178 ;
  assign n323 = n95 & n128 ;
  assign n324 = n129 | n323 ;
  assign n325 = n322 | n324 ;
  assign n326 = n106 | n325 ;
  assign n327 = n321 | n326 ;
  assign n328 = n122 & n132 ;
  assign n329 = n142 | n328 ;
  assign n330 = n105 & n117 ;
  assign n331 = n114 & n128 ;
  assign n332 = n330 | n331 ;
  assign n333 = n122 & n128 ;
  assign n334 = n95 & n132 ;
  assign n335 = n333 | n334 ;
  assign n336 = n332 | n335 ;
  assign n337 = n329 | n336 ;
  assign n338 = n327 | n337 ;
  assign n339 = n320 | n338 ;
  assign n340 = n233 | n339 ;
  assign n341 = n134 | n340 ;
  assign n342 = n124 | n341 ;
  assign n343 = n69 & n197 ;
  assign n344 = n69 & n178 ;
  assign n345 = n69 & n119 ;
  assign n346 = ~n98 & n119 ;
  assign n347 = ~n98 & n108 ;
  assign n348 = n346 | n347 ;
  assign n349 = n345 | n348 ;
  assign n350 = n172 | n349 ;
  assign n351 = n344 | n350 ;
  assign n352 = n343 | n351 ;
  assign n353 = n342 | n352 ;
  assign n354 = n313 | n353 ;
  assign n355 = n312 | n354 ;
  assign n356 = n311 | n355 ;
  assign n357 = n170 | n233 ;
  assign n358 = n69 & n114 ;
  assign n286 = n125 & n176 ;
  assign n305 = n122 & n179 ;
  assign n359 = n183 | n305 ;
  assign n360 = n333 | n359 ;
  assign n361 = n129 | n214 ;
  assign n362 = n360 | n361 ;
  assign n363 = n221 | n362 ;
  assign n364 = n286 | n363 ;
  assign n365 = n169 | n364 ;
  assign n366 = n358 | n365 ;
  assign n367 = n190 | n366 ;
  assign n368 = n142 | n367 ;
  assign n264 = n108 & n179 ;
  assign n369 = n150 | n264 ;
  assign n281 = n176 & n197 ;
  assign n370 = n205 | n281 ;
  assign n371 = n162 | n370 ;
  assign n372 = n369 | n371 ;
  assign n373 = n368 | n372 ;
  assign n374 = n357 | n373 ;
  assign n304 = n105 & n179 ;
  assign n268 = n105 & n128 ;
  assign n375 = n215 | n268 ;
  assign n376 = n117 & n174 ;
  assign n377 = n225 | n376 ;
  assign n378 = n375 | n377 ;
  assign n379 = n304 | n378 ;
  assign n267 = n108 & n176 ;
  assign n380 = n267 | n328 ;
  assign n381 = n379 | n380 ;
  assign n382 = n115 | n381 ;
  assign n383 = ~n98 & n114 ;
  assign n283 = n174 & n179 ;
  assign n284 = n114 & n179 ;
  assign n285 = n283 | n284 ;
  assign n384 = n69 & n149 ;
  assign n385 = n148 | n384 ;
  assign n386 = n285 | n385 ;
  assign n387 = n177 | n204 ;
  assign n388 = n386 | n387 ;
  assign n389 = n103 & n197 ;
  assign n390 = n156 | n389 ;
  assign n391 = n234 | n390 ;
  assign n392 = n388 | n391 ;
  assign n393 = n383 | n392 ;
  assign n394 = ~n98 & n125 ;
  assign n262 = n100 & n176 ;
  assign n263 = n147 & n176 ;
  assign n395 = n262 | n263 ;
  assign n396 = n182 | n395 ;
  assign n397 = n117 & n178 ;
  assign n398 = n112 | n397 ;
  assign n399 = n396 | n398 ;
  assign n400 = n69 & n111 ;
  assign n265 = n119 & n176 ;
  assign n259 = n122 & n176 ;
  assign n401 = n196 | n259 ;
  assign n402 = n155 | n401 ;
  assign n403 = n265 | n402 ;
  assign n404 = n331 | n403 ;
  assign n405 = n151 | n404 ;
  assign n406 = n400 | n405 ;
  assign n407 = n399 | n406 ;
  assign n408 = n206 | n407 ;
  assign n409 = n185 | n408 ;
  assign n410 = n224 | n409 ;
  assign n411 = n158 | n410 ;
  assign n412 = n235 | n411 ;
  assign n413 = n394 | n412 ;
  assign n260 = n105 & n176 ;
  assign n414 = ~n98 & n197 ;
  assign n415 = n260 | n414 ;
  assign n416 = n413 | n415 ;
  assign n282 = n125 & n179 ;
  assign n417 = n220 | n282 ;
  assign n418 = n103 & n174 ;
  assign n419 = n199 | n418 ;
  assign n420 = n417 | n419 ;
  assign n421 = n416 | n420 ;
  assign n422 = n161 | n323 ;
  assign n423 = n117 & n197 ;
  assign n293 = n179 & n197 ;
  assign n424 = n222 | n293 ;
  assign n425 = n423 | n424 ;
  assign n426 = n422 | n425 ;
  assign n427 = n421 | n426 ;
  assign n428 = n393 | n427 ;
  assign n429 = n134 | n157 ;
  assign n430 = n69 & n125 ;
  assign n431 = n246 | n430 ;
  assign n432 = n429 | n431 ;
  assign n433 = n428 | n432 ;
  assign n434 = n382 | n433 ;
  assign n435 = n374 | n434 ;
  assign n436 = ~n98 & n111 ;
  assign n437 = n236 | n334 ;
  assign n438 = n436 | n437 ;
  assign n439 = n146 | n438 ;
  assign n440 = n435 | n439 ;
  assign n272 = n128 & n147 ;
  assign n278 = n132 & n178 ;
  assign n441 = n272 | n278 ;
  assign n442 = n414 | n441 ;
  assign n443 = n158 | n442 ;
  assign n444 = n397 | n443 ;
  assign n277 = n119 & n132 ;
  assign n445 = n204 | n277 ;
  assign n446 = n157 | n445 ;
  assign n447 = n293 | n446 ;
  assign n448 = n334 | n447 ;
  assign n449 = n106 | n448 ;
  assign n450 = n347 | n449 ;
  assign n451 = n103 & n149 ;
  assign n452 = n304 | n451 ;
  assign n453 = n423 | n452 ;
  assign n454 = n376 | n453 ;
  assign n455 = n344 | n454 ;
  assign n456 = n213 | n323 ;
  assign n457 = n151 | n456 ;
  assign n458 = n316 | n457 ;
  assign n459 = n117 & n149 ;
  assign n460 = n263 | n400 ;
  assign n461 = n182 | n460 ;
  assign n462 = n126 | n315 ;
  assign n463 = n221 | n321 ;
  assign n464 = n462 | n463 ;
  assign n465 = n461 | n464 ;
  assign n466 = n205 | n285 ;
  assign n467 = n199 | n466 ;
  assign n468 = n177 | n467 ;
  assign n469 = n465 | n468 ;
  assign n271 = n132 & n147 ;
  assign n470 = n271 | n358 ;
  assign n471 = n469 | n470 ;
  assign n472 = n281 | n471 ;
  assign n473 = n459 | n472 ;
  assign n474 = n143 | n184 ;
  assign n475 = n473 | n474 ;
  assign n476 = n330 | n389 ;
  assign n477 = n154 | n476 ;
  assign n478 = n475 | n477 ;
  assign n479 = n458 | n478 ;
  assign n480 = n455 | n479 ;
  assign n481 = n450 | n480 ;
  assign n292 = n119 & n128 ;
  assign n482 = n225 | n369 ;
  assign n483 = n267 | n482 ;
  assign n484 = n292 | n483 ;
  assign n485 = n156 | n484 ;
  assign n486 = n418 | n485 ;
  assign n487 = n346 | n486 ;
  assign n488 = n123 | n383 ;
  assign n489 = n282 | n286 ;
  assign n490 = n488 | n489 ;
  assign n491 = n146 | n490 ;
  assign n492 = n189 | n191 ;
  assign n493 = n345 | n492 ;
  assign n494 = n95 & n103 ;
  assign n495 = n169 | n494 ;
  assign n496 = n96 | n495 ;
  assign n497 = n260 | n265 ;
  assign n498 = n183 | n497 ;
  assign n499 = n496 | n498 ;
  assign n500 = n493 | n499 ;
  assign n501 = n491 | n500 ;
  assign n502 = n487 | n501 ;
  assign n503 = n224 | n502 ;
  assign n504 = n245 | n331 ;
  assign n505 = n503 | n504 ;
  assign n506 = n481 | n505 ;
  assign n507 = n444 | n506 ;
  assign n508 = n436 | n507 ;
  assign n509 = n440 & n508 ;
  assign n510 = n356 & ~n509 ;
  assign n511 = pi14 & pi22 ;
  assign n512 = pi14 & n35 ;
  assign n513 = ( pi14 & n44 ) | ( pi14 & n512 ) | ( n44 & n512 );
  assign n514 = n45 & ~n513 ;
  assign n515 = pi22 & ~n511 ;
  assign n516 = ( n511 & n514 ) | ( n511 & ~n515 ) | ( n514 & ~n515 );
  assign n517 = n440 | n508 ;
  assign n518 = ~n356 & n517 ;
  assign n519 = n440 & ~n508 ;
  assign n520 = ~n440 & n508 ;
  assign n521 = n519 | n520 ;
  assign n522 = n518 | n521 ;
  assign n523 = n516 & ~n522 ;
  assign n524 = n510 | n521 ;
  assign n525 = n516 & ~n524 ;
  assign n526 = ( n510 & ~n523 ) | ( n510 & n525 ) | ( ~n523 & n525 );
  assign n261 = n259 | n260 ;
  assign n266 = n264 | n265 ;
  assign n269 = n267 | n268 ;
  assign n270 = n266 | n269 ;
  assign n273 = n271 | n272 ;
  assign n274 = n270 | n273 ;
  assign n275 = n263 | n274 ;
  assign n276 = n262 | n275 ;
  assign n279 = n128 & n178 ;
  assign n280 = n278 | n279 ;
  assign n287 = n111 & n132 ;
  assign n288 = n286 | n287 ;
  assign n289 = n114 & n132 ;
  assign n290 = n111 & n128 ;
  assign n291 = n289 | n290 ;
  assign n294 = n292 | n293 ;
  assign n295 = n291 | n294 ;
  assign n296 = n288 | n295 ;
  assign n297 = n285 | n296 ;
  assign n298 = n282 | n297 ;
  assign n299 = n281 | n298 ;
  assign n300 = n280 | n299 ;
  assign n301 = n277 | n300 ;
  assign n302 = n177 | n301 ;
  assign n303 = n276 | n302 ;
  assign n306 = n304 | n305 ;
  assign n307 = n303 | n306 ;
  assign n308 = n228 | n307 ;
  assign n309 = n219 | n308 ;
  assign n310 = n261 | n309 ;
  assign n527 = ~n310 & n526 ;
  assign n528 = ( ~pi11 & n526 ) | ( ~pi11 & n527 ) | ( n526 & n527 );
  assign n529 = ~pi22 & n256 ;
  assign n530 = ( n526 & n527 ) | ( n526 & ~n529 ) | ( n527 & ~n529 );
  assign n531 = pi11 | pi22 ;
  assign n532 = ( n526 & n527 ) | ( n526 & n531 ) | ( n527 & n531 );
  assign n533 = ( ~n44 & n530 ) | ( ~n44 & n532 ) | ( n530 & n532 );
  assign n534 = ( n258 & n528 ) | ( n258 & n533 ) | ( n528 & n533 );
  assign n535 = n310 & ~n526 ;
  assign n536 = pi11 & n535 ;
  assign n537 = n529 & n535 ;
  assign n538 = ~n531 & n535 ;
  assign n539 = ( n44 & n537 ) | ( n44 & n538 ) | ( n537 & n538 );
  assign n540 = ( ~n258 & n536 ) | ( ~n258 & n539 ) | ( n536 & n539 );
  assign n541 = n534 | n540 ;
  assign n542 = pi12 & ~pi22 ;
  assign n543 = ( ~pi22 & n33 ) | ( ~pi22 & n542 ) | ( n33 & n542 );
  assign n544 = pi13 & n543 ;
  assign n545 = pi13 & ~pi22 ;
  assign n546 = ( n44 & n544 ) | ( n44 & n545 ) | ( n544 & n545 );
  assign n547 = pi13 & ~n546 ;
  assign n548 = n100 & n103 ;
  assign n549 = n100 & n117 ;
  assign n550 = n451 | n549 ;
  assign n551 = n548 | n550 ;
  assign n552 = n117 & n122 ;
  assign n553 = n95 & n117 ;
  assign n554 = n552 | n553 ;
  assign n555 = n551 | n554 ;
  assign n556 = n103 & n122 ;
  assign n557 = n459 | n494 ;
  assign n558 = n556 | n557 ;
  assign n559 = n555 | n558 ;
  assign n560 = n238 | n398 ;
  assign n561 = n115 | n560 ;
  assign n562 = n389 | n561 ;
  assign n563 = n418 | n423 ;
  assign n564 = n562 | n563 ;
  assign n565 = n376 | n564 ;
  assign n566 = n342 | n565 ;
  assign n567 = n159 | n566 ;
  assign n568 = n152 | n567 ;
  assign n569 = n559 | n568 ;
  assign n570 = n126 | n569 ;
  assign n571 = n356 | n570 ;
  assign n572 = ~n310 & n571 ;
  assign n573 = ~n356 & n570 ;
  assign n574 = n356 & ~n570 ;
  assign n575 = n573 | n574 ;
  assign n576 = ~n572 & n575 ;
  assign n577 = ~n546 & n576 ;
  assign n578 = ( ~pi22 & n44 ) | ( ~pi22 & n543 ) | ( n44 & n543 );
  assign n579 = n576 & n578 ;
  assign n580 = ( n547 & n577 ) | ( n547 & n579 ) | ( n577 & n579 );
  assign n581 = n541 | n580 ;
  assign n582 = n572 | n575 ;
  assign n583 = pi12 & pi22 ;
  assign n584 = pi12 & n33 ;
  assign n585 = ( pi12 & n44 ) | ( pi12 & n584 ) | ( n44 & n584 );
  assign n586 = n578 & ~n585 ;
  assign n587 = n583 | n586 ;
  assign n588 = n356 & n570 ;
  assign n589 = n310 & ~n588 ;
  assign n590 = n575 & ~n589 ;
  assign n591 = n546 & n590 ;
  assign n592 = ~n578 & n590 ;
  assign n593 = ( ~n547 & n591 ) | ( ~n547 & n592 ) | ( n591 & n592 );
  assign n594 = ( ~n582 & n587 ) | ( ~n582 & n593 ) | ( n587 & n593 );
  assign n595 = n575 | n589 ;
  assign n596 = ( n587 & ~n593 ) | ( n587 & n595 ) | ( ~n593 & n595 );
  assign n597 = ~n594 & n596 ;
  assign n598 = ~n581 & n597 ;
  assign n599 = ( ~n546 & n547 ) | ( ~n546 & n578 ) | ( n547 & n578 );
  assign n600 = ~n515 & n576 ;
  assign n601 = n511 & n576 ;
  assign n602 = ( n514 & n600 ) | ( n514 & n601 ) | ( n600 & n601 );
  assign n603 = n515 & n590 ;
  assign n604 = ~n511 & n590 ;
  assign n605 = ( ~n514 & n603 ) | ( ~n514 & n604 ) | ( n603 & n604 );
  assign n606 = n602 | n605 ;
  assign n607 = ( n595 & n599 ) | ( n595 & ~n606 ) | ( n599 & ~n606 );
  assign n608 = ( ~n582 & n599 ) | ( ~n582 & n606 ) | ( n599 & n606 );
  assign n609 = n607 & ~n608 ;
  assign n610 = n534 & n609 ;
  assign n611 = ( n598 & n609 ) | ( n598 & n610 ) | ( n609 & n610 );
  assign n612 = n534 | n609 ;
  assign n613 = n598 | n612 ;
  assign n614 = ~n611 & n613 ;
  assign n615 = ~n310 & n510 ;
  assign n616 = ( ~pi11 & n510 ) | ( ~pi11 & n615 ) | ( n510 & n615 );
  assign n617 = ( n510 & ~n529 ) | ( n510 & n615 ) | ( ~n529 & n615 );
  assign n618 = ( n510 & n531 ) | ( n510 & n615 ) | ( n531 & n615 );
  assign n619 = ( ~n44 & n617 ) | ( ~n44 & n618 ) | ( n617 & n618 );
  assign n620 = ( n258 & n616 ) | ( n258 & n619 ) | ( n616 & n619 );
  assign n621 = n310 & ~n510 ;
  assign n622 = pi11 & n621 ;
  assign n623 = n529 & n621 ;
  assign n624 = ~n531 & n621 ;
  assign n625 = ( n44 & n623 ) | ( n44 & n624 ) | ( n623 & n624 );
  assign n626 = ( ~n258 & n622 ) | ( ~n258 & n625 ) | ( n622 & n625 );
  assign n627 = n620 | n626 ;
  assign n628 = n310 & n583 ;
  assign n629 = ( n310 & n586 ) | ( n310 & n628 ) | ( n586 & n628 );
  assign n630 = ~n627 & n629 ;
  assign n631 = n627 & ~n629 ;
  assign n632 = n630 | n631 ;
  assign n633 = n614 & ~n632 ;
  assign n634 = ~n614 & n632 ;
  assign n635 = n633 | n634 ;
  assign n636 = n541 & n580 ;
  assign n637 = ( n541 & ~n597 ) | ( n541 & n636 ) | ( ~n597 & n636 );
  assign n638 = n598 | n637 ;
  assign n639 = n177 | n264 ;
  assign n640 = n106 | n639 ;
  assign n641 = n124 | n225 ;
  assign n642 = n347 | n641 ;
  assign n643 = n640 | n642 ;
  assign n644 = n360 | n643 ;
  assign n645 = n184 | n418 ;
  assign n646 = n311 | n330 ;
  assign n647 = n645 | n646 ;
  assign n648 = n190 | n647 ;
  assign n649 = n644 | n648 ;
  assign n650 = n189 | n279 ;
  assign n651 = n271 | n650 ;
  assign n652 = n553 | n651 ;
  assign n653 = n148 | n652 ;
  assign n654 = n649 | n653 ;
  assign n655 = n131 | n272 ;
  assign n656 = n96 | n655 ;
  assign n657 = n162 | n656 ;
  assign n658 = n198 | n221 ;
  assign n659 = n328 | n430 ;
  assign n660 = n144 | n659 ;
  assign n661 = n462 | n660 ;
  assign n662 = n101 | n661 ;
  assign n663 = n313 | n662 ;
  assign n664 = n109 | n663 ;
  assign n665 = n556 | n664 ;
  assign n666 = n416 | n665 ;
  assign n667 = n658 | n666 ;
  assign n668 = n195 | n267 ;
  assign n669 = n191 | n203 ;
  assign n670 = n668 | n669 ;
  assign n671 = n667 | n670 ;
  assign n672 = n657 | n671 ;
  assign n673 = n156 | n672 ;
  assign n674 = n654 | n673 ;
  assign n675 = n452 | n552 ;
  assign n676 = n240 | n675 ;
  assign n677 = n345 | n676 ;
  assign n678 = n674 | n677 ;
  assign n679 = n279 | n331 ;
  assign n680 = n370 | n679 ;
  assign n681 = n126 | n213 ;
  assign n682 = n680 | n681 ;
  assign n683 = n358 | n389 ;
  assign n684 = n150 | n430 ;
  assign n685 = n106 | n170 ;
  assign n686 = n384 | n685 ;
  assign n687 = n684 | n686 ;
  assign n688 = n683 | n687 ;
  assign n689 = n682 | n688 ;
  assign n690 = n185 | n200 ;
  assign n691 = n321 | n436 ;
  assign n692 = n690 | n691 ;
  assign n693 = n312 | n692 ;
  assign n694 = n196 | n220 ;
  assign n695 = n115 | n694 ;
  assign n696 = n199 | n287 ;
  assign n697 = n127 | n553 ;
  assign n698 = n696 | n697 ;
  assign n699 = n169 | n346 ;
  assign n700 = n698 | n699 ;
  assign n701 = n129 | n328 ;
  assign n702 = n191 | n701 ;
  assign n703 = n700 | n702 ;
  assign n704 = n695 | n703 ;
  assign n705 = n693 | n704 ;
  assign n706 = n689 | n705 ;
  assign n707 = n215 | n222 ;
  assign n708 = n190 | n707 ;
  assign n709 = n459 | n708 ;
  assign n710 = n131 | n709 ;
  assign n711 = n313 | n710 ;
  assign n712 = n347 | n711 ;
  assign n713 = n241 | n712 ;
  assign n714 = n293 | n548 ;
  assign n715 = n376 | n714 ;
  assign n716 = n234 | n715 ;
  assign n717 = n414 | n716 ;
  assign n718 = n160 | n717 ;
  assign n719 = n153 | n718 ;
  assign n720 = n195 | n277 ;
  assign n721 = n240 | n397 ;
  assign n722 = n720 | n721 ;
  assign n723 = n283 | n722 ;
  assign n724 = n112 | n723 ;
  assign n725 = n719 | n724 ;
  assign n726 = n109 | n556 ;
  assign n727 = n148 | n726 ;
  assign n728 = n725 | n727 ;
  assign n729 = n123 | n728 ;
  assign n730 = n713 | n729 ;
  assign n731 = n706 | n730 ;
  assign n732 = n206 | n272 ;
  assign n733 = n271 | n732 ;
  assign n734 = n96 | n733 ;
  assign n735 = n731 | n734 ;
  assign n736 = n678 & n735 ;
  assign n737 = n508 & ~n736 ;
  assign n738 = ~pi22 & n41 ;
  assign n739 = ( ~pi22 & n42 ) | ( ~pi22 & n738 ) | ( n42 & n738 );
  assign n740 = pi9 & ~n739 ;
  assign n741 = ~pi9 & n739 ;
  assign n742 = n740 | n741 ;
  assign n743 = n310 & n742 ;
  assign n744 = ~n737 & n743 ;
  assign n745 = n737 & ~n743 ;
  assign n746 = n744 | n745 ;
  assign n747 = ~pi22 & n44 ;
  assign n748 = ~pi10 & n747 ;
  assign n749 = pi10 | n748 ;
  assign n750 = ( ~n747 & n748 ) | ( ~n747 & n749 ) | ( n748 & n749 );
  assign n751 = n310 & n750 ;
  assign n752 = ~n746 & n751 ;
  assign n753 = n744 | n752 ;
  assign n754 = ~n510 & n521 ;
  assign n755 = ~n516 & n754 ;
  assign n756 = ( n524 & n599 ) | ( n524 & ~n755 ) | ( n599 & ~n755 );
  assign n757 = ( ~n522 & n599 ) | ( ~n522 & n755 ) | ( n599 & n755 );
  assign n758 = n756 & ~n757 ;
  assign n759 = n576 & n587 ;
  assign n760 = ( n44 & n529 ) | ( n44 & ~n531 ) | ( n529 & ~n531 );
  assign n761 = ( pi11 & ~n258 ) | ( pi11 & n760 ) | ( ~n258 & n760 );
  assign n762 = ~n587 & n590 ;
  assign n763 = ( ~n582 & n761 ) | ( ~n582 & n762 ) | ( n761 & n762 );
  assign n764 = ( n595 & n761 ) | ( n595 & ~n762 ) | ( n761 & ~n762 );
  assign n765 = ~n763 & n764 ;
  assign n766 = ~n759 & n765 ;
  assign n767 = ~n518 & n521 ;
  assign n768 = ~n516 & n766 ;
  assign n769 = ( n766 & ~n767 ) | ( n766 & n768 ) | ( ~n767 & n768 );
  assign n770 = n758 & n769 ;
  assign n771 = n678 | n735 ;
  assign n772 = ~n508 & n771 ;
  assign n773 = n678 & ~n735 ;
  assign n774 = ~n678 & n735 ;
  assign n775 = n773 | n774 ;
  assign n776 = n772 | n775 ;
  assign n777 = n516 & ~n776 ;
  assign n778 = n737 | n775 ;
  assign n779 = n516 & ~n778 ;
  assign n780 = ( n737 & ~n777 ) | ( n737 & n779 ) | ( ~n777 & n779 );
  assign n781 = ~n743 & n780 ;
  assign n782 = n599 & n767 ;
  assign n783 = ~n599 & n754 ;
  assign n784 = ( n524 & n587 ) | ( n524 & ~n783 ) | ( n587 & ~n783 );
  assign n785 = ( ~n522 & n587 ) | ( ~n522 & n783 ) | ( n587 & n783 );
  assign n786 = n784 & ~n785 ;
  assign n787 = ~n782 & n786 ;
  assign n788 = n743 & ~n780 ;
  assign n789 = n781 | n788 ;
  assign n790 = n787 & ~n789 ;
  assign n791 = n781 | n790 ;
  assign n792 = n516 & ~n766 ;
  assign n793 = n767 & n792 ;
  assign n794 = ( n758 & n766 ) | ( n758 & ~n793 ) | ( n766 & ~n793 );
  assign n795 = ~n770 & n794 ;
  assign n796 = n791 & n795 ;
  assign n797 = n770 | n796 ;
  assign n798 = ( ~n638 & n753 ) | ( ~n638 & n797 ) | ( n753 & n797 );
  assign n799 = ~n635 & n798 ;
  assign n800 = n635 & ~n798 ;
  assign n801 = n799 | n800 ;
  assign n802 = n515 | n582 ;
  assign n803 = n511 & ~n582 ;
  assign n804 = ( n514 & ~n802 ) | ( n514 & n803 ) | ( ~n802 & n803 );
  assign n805 = n511 | n589 ;
  assign n806 = ~n590 & n805 ;
  assign n807 = n515 & ~n589 ;
  assign n808 = n590 | n807 ;
  assign n809 = ( n514 & n806 ) | ( n514 & ~n808 ) | ( n806 & ~n808 );
  assign n810 = ~n804 & n809 ;
  assign n811 = n626 | n629 ;
  assign n812 = ( n626 & ~n627 ) | ( n626 & n811 ) | ( ~n627 & n811 );
  assign n813 = n310 & ~n546 ;
  assign n814 = n310 & n543 ;
  assign n815 = ~pi22 & n310 ;
  assign n816 = ( n44 & n814 ) | ( n44 & n815 ) | ( n814 & n815 );
  assign n817 = ( n547 & n813 ) | ( n547 & n816 ) | ( n813 & n816 );
  assign n818 = ( n810 & n812 ) | ( n810 & ~n817 ) | ( n812 & ~n817 );
  assign n819 = ( n810 & n812 ) | ( n810 & ~n818 ) | ( n812 & ~n818 );
  assign n820 = ( n817 & n818 ) | ( n817 & ~n819 ) | ( n818 & ~n819 );
  assign n821 = ~n609 & n632 ;
  assign n822 = ~n598 & n632 ;
  assign n823 = ( ~n610 & n821 ) | ( ~n610 & n822 ) | ( n821 & n822 );
  assign n824 = n820 & n823 ;
  assign n825 = ~n611 & n820 ;
  assign n826 = ( ~n614 & n824 ) | ( ~n614 & n825 ) | ( n824 & n825 );
  assign n827 = n818 | n826 ;
  assign n828 = n810 | n817 ;
  assign n829 = n812 | n828 ;
  assign n830 = ( n818 & ~n819 ) | ( n818 & n829 ) | ( ~n819 & n829 );
  assign n831 = n823 | n830 ;
  assign n832 = n611 & ~n830 ;
  assign n833 = ( n614 & ~n831 ) | ( n614 & n832 ) | ( ~n831 & n832 );
  assign n834 = ( n801 & n827 ) | ( n801 & ~n833 ) | ( n827 & ~n833 );
  assign n835 = ( n799 & ~n827 ) | ( n799 & n833 ) | ( ~n827 & n833 );
  assign n836 = n753 & n797 ;
  assign n837 = n753 & ~n836 ;
  assign n838 = n797 & ~n836 ;
  assign n839 = n837 | n838 ;
  assign n840 = n638 & ~n839 ;
  assign n841 = ~n638 & n839 ;
  assign n842 = n840 | n841 ;
  assign n843 = n576 & n761 ;
  assign n844 = n590 & ~n761 ;
  assign n845 = ( n595 & n750 ) | ( n595 & ~n844 ) | ( n750 & ~n844 );
  assign n846 = ( ~n582 & n750 ) | ( ~n582 & n844 ) | ( n750 & n844 );
  assign n847 = n845 & ~n846 ;
  assign n848 = ~n843 & n847 ;
  assign n849 = pi7 & ~n738 ;
  assign n850 = ~pi7 & n738 ;
  assign n851 = n849 | n850 ;
  assign n852 = n310 & n851 ;
  assign n853 = n423 | n553 ;
  assign n854 = n224 | n259 ;
  assign n855 = n289 | n854 ;
  assign n856 = n853 | n855 ;
  assign n857 = n268 | n288 ;
  assign n858 = n856 | n857 ;
  assign n859 = n106 | n858 ;
  assign n860 = n292 | n347 ;
  assign n861 = n222 | n279 ;
  assign n862 = n860 | n861 ;
  assign n863 = n241 | n862 ;
  assign n864 = n115 | n124 ;
  assign n865 = n863 | n864 ;
  assign n866 = n859 | n865 ;
  assign n867 = n135 | n463 ;
  assign n868 = n436 | n867 ;
  assign n869 = n123 | n345 ;
  assign n870 = n868 | n869 ;
  assign n871 = n866 | n870 ;
  assign n872 = n181 | n871 ;
  assign n873 = n184 | n304 ;
  assign n874 = n872 | n873 ;
  assign n875 = n112 | n548 ;
  assign n876 = n400 | n875 ;
  assign n877 = n874 | n876 ;
  assign n878 = n183 | n202 ;
  assign n879 = n397 | n878 ;
  assign n880 = n143 | n146 ;
  assign n881 = n879 | n880 ;
  assign n882 = n283 | n290 ;
  assign n883 = n377 | n496 ;
  assign n884 = n882 | n883 ;
  assign n885 = n881 | n884 ;
  assign n886 = n333 | n343 ;
  assign n887 = n330 | n886 ;
  assign n888 = n312 | n887 ;
  assign n889 = n885 | n888 ;
  assign n890 = n190 | n889 ;
  assign n891 = n203 | n890 ;
  assign n892 = n150 | n220 ;
  assign n893 = n213 | n278 ;
  assign n894 = n892 | n893 ;
  assign n895 = n240 | n271 ;
  assign n896 = n161 | n895 ;
  assign n897 = n894 | n896 ;
  assign n898 = n141 & ~n195 ;
  assign n899 = n120 | n260 ;
  assign n900 = n153 | n899 ;
  assign n901 = n196 | n263 ;
  assign n902 = n414 | n901 ;
  assign n903 = n446 | n550 ;
  assign n904 = n902 | n903 ;
  assign n905 = n900 | n904 ;
  assign n906 = n898 & ~n905 ;
  assign n907 = ~n897 & n906 ;
  assign n908 = ~n126 & n907 ;
  assign n909 = ~n891 & n908 ;
  assign n910 = ~n328 & n909 ;
  assign n911 = ~n877 & n910 ;
  assign n912 = n101 | n214 ;
  assign n913 = n245 | n912 ;
  assign n914 = n911 & ~n913 ;
  assign n915 = n213 | n279 ;
  assign n916 = n494 | n915 ;
  assign n917 = n334 | n418 ;
  assign n918 = n127 | n917 ;
  assign n919 = n263 | n918 ;
  assign n920 = n916 | n919 ;
  assign n921 = n235 | n459 ;
  assign n922 = n121 | n292 ;
  assign n923 = n157 | n922 ;
  assign n924 = n346 | n923 ;
  assign n925 = n224 | n264 ;
  assign n926 = n304 | n925 ;
  assign n927 = n316 | n926 ;
  assign n928 = n361 | n927 ;
  assign n929 = n222 | n260 ;
  assign n930 = n206 | n929 ;
  assign n931 = n189 | n281 ;
  assign n932 = n930 | n931 ;
  assign n933 = n888 | n932 ;
  assign n934 = n928 | n933 ;
  assign n935 = n225 | n305 ;
  assign n936 = n204 | n935 ;
  assign n937 = n934 | n936 ;
  assign n938 = n156 | n311 ;
  assign n939 = n655 | n938 ;
  assign n940 = n267 | n293 ;
  assign n941 = n414 | n436 ;
  assign n942 = n940 | n941 ;
  assign n943 = n939 | n942 ;
  assign n944 = n937 | n943 ;
  assign n945 = n924 | n944 ;
  assign n946 = n285 | n945 ;
  assign n947 = n169 | n344 ;
  assign n948 = n200 | n271 ;
  assign n949 = n313 | n948 ;
  assign n950 = n947 | n949 ;
  assign n951 = n221 | n950 ;
  assign n952 = n290 | n951 ;
  assign n953 = n134 | n952 ;
  assign n954 = n553 | n953 ;
  assign n955 = n946 | n954 ;
  assign n956 = n921 | n955 ;
  assign n957 = n406 | n956 ;
  assign n958 = n920 | n957 ;
  assign n959 = n203 | n376 ;
  assign n960 = n146 | n959 ;
  assign n961 = n958 | n960 ;
  assign n962 = ~n914 & n961 ;
  assign n963 = n735 & ~n962 ;
  assign n964 = n852 & ~n963 ;
  assign n965 = pi8 & pi22 ;
  assign n966 = pi7 | n41 ;
  assign n967 = pi8 & n966 ;
  assign n968 = n739 & ~n967 ;
  assign n969 = n965 | n968 ;
  assign n970 = ~n852 & n963 ;
  assign n971 = n964 | n970 ;
  assign n972 = n969 & ~n971 ;
  assign n973 = n310 & n972 ;
  assign n974 = n964 | n973 ;
  assign n975 = n848 & n974 ;
  assign n976 = n848 & ~n975 ;
  assign n977 = n974 & ~n975 ;
  assign n978 = n976 | n977 ;
  assign n979 = n576 & n750 ;
  assign n980 = n590 & ~n750 ;
  assign n981 = ( n595 & n742 ) | ( n595 & ~n980 ) | ( n742 & ~n980 );
  assign n982 = ( ~n582 & n742 ) | ( ~n582 & n980 ) | ( n742 & n980 );
  assign n983 = n981 & ~n982 ;
  assign n984 = ~n979 & n983 ;
  assign n985 = ~n772 & n775 ;
  assign n986 = n516 & n985 ;
  assign n987 = ~n737 & n775 ;
  assign n988 = ~n516 & n987 ;
  assign n989 = ( n599 & n778 ) | ( n599 & ~n988 ) | ( n778 & ~n988 );
  assign n990 = ( n599 & ~n776 ) | ( n599 & n988 ) | ( ~n776 & n988 );
  assign n991 = n989 & ~n990 ;
  assign n992 = ~n986 & n991 ;
  assign n993 = n587 & n767 ;
  assign n994 = ~n587 & n754 ;
  assign n995 = ( n524 & n761 ) | ( n524 & ~n994 ) | ( n761 & ~n994 );
  assign n996 = ( ~n522 & n761 ) | ( ~n522 & n994 ) | ( n761 & n994 );
  assign n997 = n995 & ~n996 ;
  assign n998 = ~n993 & n997 ;
  assign n999 = ( n984 & n992 ) | ( n984 & n998 ) | ( n992 & n998 );
  assign n1000 = n978 & n999 ;
  assign n1001 = n978 & ~n1000 ;
  assign n1002 = n576 & n742 ;
  assign n1003 = n590 & ~n742 ;
  assign n1004 = ( n595 & n969 ) | ( n595 & ~n1003 ) | ( n969 & ~n1003 );
  assign n1005 = ( ~n582 & n969 ) | ( ~n582 & n1003 ) | ( n969 & n1003 );
  assign n1006 = n1004 & ~n1005 ;
  assign n1007 = ~n1002 & n1006 ;
  assign n1008 = n761 & n767 ;
  assign n1009 = n754 & ~n761 ;
  assign n1010 = ( n524 & n750 ) | ( n524 & ~n1009 ) | ( n750 & ~n1009 );
  assign n1011 = ( ~n522 & n750 ) | ( ~n522 & n1009 ) | ( n750 & n1009 );
  assign n1012 = n1010 & ~n1011 ;
  assign n1013 = ~n1008 & n1012 ;
  assign n1014 = n1007 & n1013 ;
  assign n1015 = n225 | n343 ;
  assign n1016 = n335 | n1015 ;
  assign n1017 = n213 | n220 ;
  assign n1018 = n112 | n1017 ;
  assign n1019 = n1016 | n1018 ;
  assign n1020 = n241 | n552 ;
  assign n1021 = n1019 | n1020 ;
  assign n1022 = n153 | n451 ;
  assign n1023 = n280 | n1022 ;
  assign n1024 = n314 | n322 ;
  assign n1025 = n1023 | n1024 ;
  assign n1026 = n246 | n311 ;
  assign n1027 = n198 | n284 ;
  assign n1028 = n1026 | n1027 ;
  assign n1029 = n401 | n1028 ;
  assign n1030 = n146 | n1029 ;
  assign n1031 = n898 & ~n1030 ;
  assign n1032 = ~n490 & n1031 ;
  assign n1033 = ~n1025 & n1032 ;
  assign n1034 = ~n1021 & n1033 ;
  assign n1035 = n369 | n864 ;
  assign n1036 = n659 | n1035 ;
  assign n1037 = n199 | n1036 ;
  assign n1038 = n203 | n1037 ;
  assign n1039 = n157 | n1038 ;
  assign n1040 = n389 | n1039 ;
  assign n1041 = n109 | n1040 ;
  assign n1042 = n345 | n1041 ;
  assign n1043 = n331 | n548 ;
  assign n1044 = n549 | n1043 ;
  assign n1045 = n134 | n272 ;
  assign n1046 = n245 | n1045 ;
  assign n1047 = n267 | n323 ;
  assign n1048 = n376 | n1047 ;
  assign n1049 = n170 | n1048 ;
  assign n1050 = n1046 | n1049 ;
  assign n1051 = n1044 | n1050 ;
  assign n1052 = n932 | n1051 ;
  assign n1053 = n462 | n1052 ;
  assign n1054 = n304 | n1053 ;
  assign n1055 = n106 | n290 ;
  assign n1056 = n1054 | n1055 ;
  assign n1057 = n344 | n1056 ;
  assign n1058 = n1042 | n1057 ;
  assign n1059 = n185 | n1058 ;
  assign n1060 = n1034 & ~n1059 ;
  assign n1061 = ~n271 & n1060 ;
  assign n1062 = ~n556 & n1061 ;
  assign n1063 = ~n131 & n1062 ;
  assign n1064 = ~n436 & n1063 ;
  assign n1065 = n235 | n552 ;
  assign n1066 = n437 | n459 ;
  assign n1067 = n1065 | n1066 ;
  assign n1068 = n206 | n282 ;
  assign n1069 = n321 | n1068 ;
  assign n1070 = n124 | n1069 ;
  assign n1071 = n685 | n1070 ;
  assign n1072 = n318 | n1071 ;
  assign n1073 = n398 | n1072 ;
  assign n1074 = n154 | n1073 ;
  assign n1075 = n285 | n1074 ;
  assign n1076 = n1067 | n1075 ;
  assign n1077 = n375 | n860 ;
  assign n1078 = n220 | n262 ;
  assign n1079 = n331 | n1078 ;
  assign n1080 = n1077 | n1079 ;
  assign n1081 = n203 | n436 ;
  assign n1082 = n240 | n1081 ;
  assign n1083 = n1080 | n1082 ;
  assign n1084 = n345 | n949 ;
  assign n1085 = n492 | n1084 ;
  assign n1086 = n141 & ~n1085 ;
  assign n1087 = ~n159 & n1086 ;
  assign n1088 = ~n1083 & n1087 ;
  assign n1089 = ~n277 & n1088 ;
  assign n1090 = ~n198 & n1089 ;
  assign n1091 = n101 | n241 ;
  assign n1092 = n1090 & ~n1091 ;
  assign n1093 = n384 | n400 ;
  assign n1094 = n1092 & ~n1093 ;
  assign n1095 = ~n1076 & n1094 ;
  assign n1096 = n329 | n1026 ;
  assign n1097 = n668 | n1096 ;
  assign n1098 = n204 | n1097 ;
  assign n1099 = n371 | n902 ;
  assign n1100 = n288 | n1099 ;
  assign n1101 = n1025 | n1100 ;
  assign n1102 = n1098 | n1101 ;
  assign n1103 = n260 | n1102 ;
  assign n1104 = n224 | n304 ;
  assign n1105 = n1103 | n1104 ;
  assign n1106 = n180 | n233 ;
  assign n1107 = n418 | n1106 ;
  assign n1108 = n1105 | n1107 ;
  assign n1109 = n394 | n553 ;
  assign n1110 = n1108 | n1109 ;
  assign n1111 = n1095 & ~n1110 ;
  assign n1112 = n181 | n190 ;
  assign n1113 = n549 | n1112 ;
  assign n1114 = n1111 & ~n1113 ;
  assign n1115 = n1064 | n1114 ;
  assign n1116 = ~n914 & n1115 ;
  assign n1117 = n1064 & ~n1116 ;
  assign n1118 = ~n1064 & n1116 ;
  assign n1119 = pi6 & pi22 ;
  assign n1120 = pi5 | n39 ;
  assign n1121 = pi6 & n1120 ;
  assign n1122 = n738 & ~n1121 ;
  assign n1123 = n1119 | n1122 ;
  assign n1124 = n310 & n1123 ;
  assign n1125 = ~n1117 & n1124 ;
  assign n1126 = ~n1118 & n1125 ;
  assign n1127 = n1117 | n1126 ;
  assign n1128 = n1007 | n1013 ;
  assign n1129 = ~n1014 & n1128 ;
  assign n1130 = n1127 & n1129 ;
  assign n1131 = n1014 | n1130 ;
  assign n1132 = n914 & ~n961 ;
  assign n1133 = n735 | n1132 ;
  assign n1134 = n914 & n961 ;
  assign n1135 = n914 | n961 ;
  assign n1136 = ~n1134 & n1135 ;
  assign n1137 = n1133 & n1136 ;
  assign n1138 = n963 | n1136 ;
  assign n1139 = ( n516 & n1137 ) | ( n516 & ~n1138 ) | ( n1137 & ~n1138 );
  assign n1140 = ( n516 & n963 ) | ( n516 & n1138 ) | ( n963 & n1138 );
  assign n1141 = ~n1139 & n1140 ;
  assign n1142 = ~n852 & n1141 ;
  assign n1143 = n852 & ~n1141 ;
  assign n1144 = n1142 | n1143 ;
  assign n1145 = n599 & n985 ;
  assign n1146 = ~n599 & n987 ;
  assign n1147 = ( n587 & n778 ) | ( n587 & ~n1146 ) | ( n778 & ~n1146 );
  assign n1148 = ( n587 & ~n776 ) | ( n587 & n1146 ) | ( ~n776 & n1146 );
  assign n1149 = n1147 & ~n1148 ;
  assign n1150 = ~n1145 & n1149 ;
  assign n1151 = ~n1144 & n1150 ;
  assign n1152 = n1142 | n1151 ;
  assign n1153 = n1131 & n1152 ;
  assign n1154 = n1131 & ~n1153 ;
  assign n1155 = n1152 & ~n1153 ;
  assign n1156 = n1154 | n1155 ;
  assign n1157 = n310 & ~n973 ;
  assign n1158 = n969 & n1157 ;
  assign n1159 = n971 | n973 ;
  assign n1160 = ~n1158 & n1159 ;
  assign n1161 = n1156 & ~n1160 ;
  assign n1162 = n1153 | n1161 ;
  assign n1163 = ~n787 & n789 ;
  assign n1164 = n790 | n1163 ;
  assign n1165 = n1162 & ~n1164 ;
  assign n1166 = ( n999 & n1162 ) | ( n999 & ~n1164 ) | ( n1162 & ~n1164 );
  assign n1167 = ( ~n978 & n1165 ) | ( ~n978 & n1166 ) | ( n1165 & n1166 );
  assign n1168 = n791 | n795 ;
  assign n1169 = ~n796 & n1168 ;
  assign n1170 = n975 | n1000 ;
  assign n1171 = n746 & ~n751 ;
  assign n1172 = n752 | n1171 ;
  assign n1173 = n1170 & ~n1172 ;
  assign n1174 = ~n1170 & n1172 ;
  assign n1175 = n1173 | n1174 ;
  assign n1176 = n1169 & ~n1175 ;
  assign n1177 = ~n1169 & n1175 ;
  assign n1178 = n1176 | n1177 ;
  assign n1179 = n1167 & ~n1178 ;
  assign n1180 = ~n1162 & n1164 ;
  assign n1181 = n1178 | n1180 ;
  assign n1182 = ( n1001 & n1179 ) | ( n1001 & ~n1181 ) | ( n1179 & ~n1181 );
  assign n1183 = n1156 & ~n1161 ;
  assign n1184 = n1160 | n1161 ;
  assign n1185 = ~n1183 & n1184 ;
  assign n1186 = n984 & ~n1185 ;
  assign n1187 = ( ~n984 & n1185 ) | ( ~n984 & n1186 ) | ( n1185 & n1186 );
  assign n1188 = n1186 | n1187 ;
  assign n1189 = n992 & ~n998 ;
  assign n1190 = ~n992 & n998 ;
  assign n1191 = n1189 | n1190 ;
  assign n1192 = n1144 & ~n1150 ;
  assign n1193 = n1151 | n1192 ;
  assign n1194 = n576 & n969 ;
  assign n1195 = n590 & ~n969 ;
  assign n1196 = ( n595 & n851 ) | ( n595 & ~n1195 ) | ( n851 & ~n1195 );
  assign n1197 = ( ~n582 & n851 ) | ( ~n582 & n1195 ) | ( n851 & n1195 );
  assign n1198 = n1196 & ~n1197 ;
  assign n1199 = ~n1194 & n1198 ;
  assign n1200 = n524 | n742 ;
  assign n1201 = ~n522 & n742 ;
  assign n1202 = n1200 & ~n1201 ;
  assign n1203 = ( n750 & n767 ) | ( n750 & ~n1202 ) | ( n767 & ~n1202 );
  assign n1204 = ( n750 & ~n754 ) | ( n750 & n1202 ) | ( ~n754 & n1202 );
  assign n1205 = ~n1203 & n1204 ;
  assign n1206 = n1133 & ~n1136 ;
  assign n1207 = ~n963 & n1136 ;
  assign n1208 = ~n599 & n1207 ;
  assign n1209 = n599 & n1137 ;
  assign n1210 = n1208 | n1209 ;
  assign n1211 = ( n516 & n1206 ) | ( n516 & n1210 ) | ( n1206 & n1210 );
  assign n1212 = ( n516 & n1138 ) | ( n516 & ~n1210 ) | ( n1138 & ~n1210 );
  assign n1213 = ~n1211 & n1212 ;
  assign n1214 = ( n1199 & n1205 ) | ( n1199 & n1213 ) | ( n1205 & n1213 );
  assign n1215 = ~n1193 & n1214 ;
  assign n1216 = n1127 | n1129 ;
  assign n1217 = ~n1130 & n1216 ;
  assign n1218 = n1193 | n1214 ;
  assign n1219 = ( ~n1214 & n1215 ) | ( ~n1214 & n1218 ) | ( n1215 & n1218 );
  assign n1220 = n1217 & ~n1219 ;
  assign n1221 = n1215 | n1220 ;
  assign n1222 = ( ~n1188 & n1191 ) | ( ~n1188 & n1221 ) | ( n1191 & n1221 );
  assign n1223 = ( n1188 & n1191 ) | ( n1188 & n1221 ) | ( n1191 & n1221 );
  assign n1224 = ( n1188 & n1222 ) | ( n1188 & ~n1223 ) | ( n1222 & ~n1223 );
  assign n1225 = n1118 | n1127 ;
  assign n1226 = n1124 & ~n1126 ;
  assign n1227 = n1225 & ~n1226 ;
  assign n1228 = n587 & n985 ;
  assign n1229 = ~n587 & n987 ;
  assign n1230 = ( n761 & n778 ) | ( n761 & ~n1229 ) | ( n778 & ~n1229 );
  assign n1231 = ( n761 & ~n776 ) | ( n761 & n1229 ) | ( ~n776 & n1229 );
  assign n1232 = n1230 & ~n1231 ;
  assign n1233 = ~n1228 & n1232 ;
  assign n1234 = ~n1227 & n1233 ;
  assign n1235 = ~pi22 & n39 ;
  assign n1236 = pi5 & ~n1235 ;
  assign n1237 = ~pi5 & n1235 ;
  assign n1238 = n1236 | n1237 ;
  assign n1239 = n310 & n1238 ;
  assign n1240 = ~n1064 & n1239 ;
  assign n1241 = n1064 & n1114 ;
  assign n1242 = n914 & ~n1241 ;
  assign n1243 = n1064 & ~n1114 ;
  assign n1244 = ~n1064 & n1114 ;
  assign n1245 = n1243 | n1244 ;
  assign n1246 = n1242 | n1245 ;
  assign n1247 = n516 & ~n1246 ;
  assign n1248 = n1116 | n1245 ;
  assign n1249 = n516 & ~n1248 ;
  assign n1250 = ( n1116 & ~n1247 ) | ( n1116 & n1249 ) | ( ~n1247 & n1249 );
  assign n1251 = ~n1240 & n1250 ;
  assign n1252 = n1064 & ~n1239 ;
  assign n1253 = ~n1240 & n1252 ;
  assign n1254 = ( n1240 & n1251 ) | ( n1240 & ~n1253 ) | ( n1251 & ~n1253 );
  assign n1255 = n1227 & ~n1233 ;
  assign n1256 = n1234 | n1255 ;
  assign n1257 = n1254 & ~n1256 ;
  assign n1258 = n1234 | n1257 ;
  assign n1259 = n599 & n1206 ;
  assign n1260 = n599 | n1138 ;
  assign n1261 = ( n587 & ~n1207 ) | ( n587 & n1260 ) | ( ~n1207 & n1260 );
  assign n1262 = ( n587 & n1137 ) | ( n587 & ~n1260 ) | ( n1137 & ~n1260 );
  assign n1263 = n1261 & ~n1262 ;
  assign n1264 = ~n1259 & n1263 ;
  assign n1265 = n761 & n985 ;
  assign n1266 = ~n761 & n987 ;
  assign n1267 = ( n750 & n778 ) | ( n750 & ~n1266 ) | ( n778 & ~n1266 );
  assign n1268 = ( n750 & ~n776 ) | ( n750 & n1266 ) | ( ~n776 & n1266 );
  assign n1269 = n1267 & ~n1268 ;
  assign n1270 = ~n1265 & n1269 ;
  assign n1271 = n742 & n767 ;
  assign n1272 = ~n742 & n754 ;
  assign n1273 = ( n524 & n969 ) | ( n524 & ~n1272 ) | ( n969 & ~n1272 );
  assign n1274 = ( ~n522 & n969 ) | ( ~n522 & n1272 ) | ( n969 & n1272 );
  assign n1275 = n1273 & ~n1274 ;
  assign n1276 = ~n1271 & n1275 ;
  assign n1277 = ( n1264 & n1270 ) | ( n1264 & n1276 ) | ( n1270 & n1276 );
  assign n1278 = ( n1199 & ~n1205 ) | ( n1199 & n1213 ) | ( ~n1205 & n1213 );
  assign n1279 = ( ~n1199 & n1205 ) | ( ~n1199 & n1278 ) | ( n1205 & n1278 );
  assign n1280 = ( ~n1213 & n1278 ) | ( ~n1213 & n1279 ) | ( n1278 & n1279 );
  assign n1281 = n1277 & n1280 ;
  assign n1282 = n576 & n851 ;
  assign n1283 = n590 & ~n851 ;
  assign n1284 = ( n595 & n1123 ) | ( n595 & ~n1283 ) | ( n1123 & ~n1283 );
  assign n1285 = ( ~n582 & n1123 ) | ( ~n582 & n1283 ) | ( n1123 & n1283 );
  assign n1286 = n1284 & ~n1285 ;
  assign n1287 = ~n1282 & n1286 ;
  assign n1288 = pi4 & pi22 ;
  assign n1289 = pi4 & n38 ;
  assign n1290 = n1235 & ~n1289 ;
  assign n1291 = n1288 | n1290 ;
  assign n1292 = n310 & n1291 ;
  assign n1293 = ~n1064 & n1292 ;
  assign n1294 = n1064 & ~n1292 ;
  assign n1295 = n1293 | n1294 ;
  assign n1296 = ~n1242 & n1245 ;
  assign n1297 = n516 & n1296 ;
  assign n1298 = ~n1116 & n1245 ;
  assign n1299 = ~n516 & n1298 ;
  assign n1300 = ( n599 & n1248 ) | ( n599 & ~n1299 ) | ( n1248 & ~n1299 );
  assign n1301 = ( n599 & ~n1246 ) | ( n599 & n1299 ) | ( ~n1246 & n1299 );
  assign n1302 = n1300 & ~n1301 ;
  assign n1303 = ~n1297 & n1302 ;
  assign n1304 = ~n1295 & n1303 ;
  assign n1305 = n1293 | n1304 ;
  assign n1306 = n1287 & n1305 ;
  assign n1307 = n1287 | n1305 ;
  assign n1308 = ~n1306 & n1307 ;
  assign n1309 = n750 & n985 ;
  assign n1310 = ~n750 & n987 ;
  assign n1311 = ( n742 & n778 ) | ( n742 & ~n1310 ) | ( n778 & ~n1310 );
  assign n1312 = ( n742 & ~n776 ) | ( n742 & n1310 ) | ( ~n776 & n1310 );
  assign n1313 = n1311 & ~n1312 ;
  assign n1314 = ~n1309 & n1313 ;
  assign n1315 = n587 & n1206 ;
  assign n1316 = n587 | n1138 ;
  assign n1317 = ( n761 & ~n1207 ) | ( n761 & n1316 ) | ( ~n1207 & n1316 );
  assign n1318 = ( n761 & n1137 ) | ( n761 & ~n1316 ) | ( n1137 & ~n1316 );
  assign n1319 = n1317 & ~n1318 ;
  assign n1320 = ~n1315 & n1319 ;
  assign n1321 = n767 & n969 ;
  assign n1322 = n754 & ~n969 ;
  assign n1323 = ( n524 & n851 ) | ( n524 & ~n1322 ) | ( n851 & ~n1322 );
  assign n1324 = ( ~n522 & n851 ) | ( ~n522 & n1322 ) | ( n851 & n1322 );
  assign n1325 = n1323 & ~n1324 ;
  assign n1326 = ~n1321 & n1325 ;
  assign n1327 = ( n1314 & n1320 ) | ( n1314 & n1326 ) | ( n1320 & n1326 );
  assign n1328 = n1308 & n1327 ;
  assign n1329 = n1306 | n1328 ;
  assign n1330 = n1277 | n1280 ;
  assign n1331 = ~n1281 & n1330 ;
  assign n1332 = n1329 & n1331 ;
  assign n1333 = n1281 | n1332 ;
  assign n1334 = ~n1217 & n1219 ;
  assign n1335 = n1220 | n1334 ;
  assign n1336 = ( n1258 & n1333 ) | ( n1258 & ~n1335 ) | ( n1333 & ~n1335 );
  assign n1337 = n1224 & ~n1336 ;
  assign n1338 = ~n1224 & n1336 ;
  assign n1339 = n1337 | n1338 ;
  assign n1340 = ( ~n1258 & n1333 ) | ( ~n1258 & n1335 ) | ( n1333 & n1335 );
  assign n1341 = ( n1258 & ~n1335 ) | ( n1258 & n1340 ) | ( ~n1335 & n1340 );
  assign n1342 = ( ~n1333 & n1340 ) | ( ~n1333 & n1341 ) | ( n1340 & n1341 );
  assign n1343 = ~n1254 & n1256 ;
  assign n1344 = n1257 | n1343 ;
  assign n1345 = n1252 | n1254 ;
  assign n1346 = n1250 & n1252 ;
  assign n1347 = ( n1250 & ~n1251 ) | ( n1250 & n1346 ) | ( ~n1251 & n1346 );
  assign n1348 = n595 | n1238 ;
  assign n1349 = ~n582 & n1238 ;
  assign n1350 = n1348 & ~n1349 ;
  assign n1351 = ( ~n590 & n1123 ) | ( ~n590 & n1350 ) | ( n1123 & n1350 );
  assign n1352 = ( n576 & n1123 ) | ( n576 & ~n1350 ) | ( n1123 & ~n1350 );
  assign n1353 = n1351 & ~n1352 ;
  assign n1354 = pi3 & ~n28 ;
  assign n1355 = ~pi3 & n28 ;
  assign n1356 = n1354 | n1355 ;
  assign n1357 = n310 & n1356 ;
  assign n1358 = n188 | n192 ;
  assign n1359 = n141 & ~n334 ;
  assign n1360 = n134 | n156 ;
  assign n1361 = n1359 & ~n1360 ;
  assign n1362 = n154 | n376 ;
  assign n1363 = n397 | n1362 ;
  assign n1364 = n1361 & ~n1363 ;
  assign n1365 = n204 | n279 ;
  assign n1366 = n553 | n1365 ;
  assign n1367 = n395 | n458 ;
  assign n1368 = n1366 | n1367 ;
  assign n1369 = n948 | n1368 ;
  assign n1370 = n357 | n1369 ;
  assign n1371 = n293 | n1370 ;
  assign n1372 = n220 | n1371 ;
  assign n1373 = n189 | n1372 ;
  assign n1374 = n494 | n1373 ;
  assign n1375 = n146 | n1374 ;
  assign n1376 = n161 | n400 ;
  assign n1377 = n385 | n1376 ;
  assign n1378 = n1375 | n1377 ;
  assign n1379 = n1364 & ~n1378 ;
  assign n1380 = ~n1358 & n1379 ;
  assign n1381 = n144 | n286 ;
  assign n1382 = n292 | n1381 ;
  assign n1383 = n328 | n1382 ;
  assign n1384 = n195 | n1383 ;
  assign n1385 = n106 | n1384 ;
  assign n1386 = n330 | n1385 ;
  assign n1387 = n245 | n1386 ;
  assign n1388 = n436 | n1387 ;
  assign n1389 = n1380 & ~n1388 ;
  assign n1390 = ~n264 & n1389 ;
  assign n1391 = ~n282 & n1390 ;
  assign n1392 = ~n451 & n1391 ;
  assign n1393 = ~n236 & n1392 ;
  assign n1394 = ~n101 & n1393 ;
  assign n1395 = ~n246 & n1394 ;
  assign n1396 = ~n430 & n1395 ;
  assign n1397 = n516 & n1396 ;
  assign n1398 = n1064 | n1397 ;
  assign n1399 = n1357 & ~n1398 ;
  assign n1400 = n599 & n1296 ;
  assign n1401 = ~n599 & n1298 ;
  assign n1402 = ( n587 & n1248 ) | ( n587 & ~n1401 ) | ( n1248 & ~n1401 );
  assign n1403 = ( n587 & ~n1246 ) | ( n587 & n1401 ) | ( ~n1246 & n1401 );
  assign n1404 = n1402 & ~n1403 ;
  assign n1405 = ~n1400 & n1404 ;
  assign n1406 = ~n1357 & n1398 ;
  assign n1407 = n1399 | n1406 ;
  assign n1408 = n1405 & ~n1407 ;
  assign n1409 = n1399 | n1408 ;
  assign n1410 = n1353 & n1409 ;
  assign n1411 = n1353 | n1409 ;
  assign n1412 = ~n1410 & n1411 ;
  assign n1413 = n742 & n985 ;
  assign n1414 = ~n742 & n987 ;
  assign n1415 = ( n778 & n969 ) | ( n778 & ~n1414 ) | ( n969 & ~n1414 );
  assign n1416 = ( ~n776 & n969 ) | ( ~n776 & n1414 ) | ( n969 & n1414 );
  assign n1417 = n1415 & ~n1416 ;
  assign n1418 = ~n1413 & n1417 ;
  assign n1419 = n761 & n1206 ;
  assign n1420 = n761 | n1138 ;
  assign n1421 = ( n750 & ~n1207 ) | ( n750 & n1420 ) | ( ~n1207 & n1420 );
  assign n1422 = ( n750 & n1137 ) | ( n750 & ~n1420 ) | ( n1137 & ~n1420 );
  assign n1423 = n1421 & ~n1422 ;
  assign n1424 = ~n1419 & n1423 ;
  assign n1425 = n767 & n851 ;
  assign n1426 = n754 & ~n851 ;
  assign n1427 = ( n524 & n1123 ) | ( n524 & ~n1426 ) | ( n1123 & ~n1426 );
  assign n1428 = ( ~n522 & n1123 ) | ( ~n522 & n1426 ) | ( n1123 & n1426 );
  assign n1429 = n1427 & ~n1428 ;
  assign n1430 = ~n1425 & n1429 ;
  assign n1431 = ( n1418 & n1424 ) | ( n1418 & n1430 ) | ( n1424 & n1430 );
  assign n1432 = n1412 & n1431 ;
  assign n1433 = n1410 | n1432 ;
  assign n1434 = ( n1264 & n1276 ) | ( n1264 & ~n1277 ) | ( n1276 & ~n1277 );
  assign n1435 = ( n1270 & ~n1277 ) | ( n1270 & n1434 ) | ( ~n1277 & n1434 );
  assign n1436 = ( n1347 & n1433 ) | ( n1347 & n1435 ) | ( n1433 & n1435 );
  assign n1437 = n1433 | n1435 ;
  assign n1438 = ( ~n1345 & n1436 ) | ( ~n1345 & n1437 ) | ( n1436 & n1437 );
  assign n1439 = ~n1344 & n1438 ;
  assign n1440 = n1344 & ~n1438 ;
  assign n1441 = n1439 | n1440 ;
  assign n1442 = n1329 | n1331 ;
  assign n1443 = ~n1332 & n1442 ;
  assign n1444 = n1439 | n1443 ;
  assign n1445 = ( n1439 & ~n1441 ) | ( n1439 & n1444 ) | ( ~n1441 & n1444 );
  assign n1446 = n1342 & ~n1445 ;
  assign n1447 = n1339 | n1446 ;
  assign n1448 = ~n1167 & n1178 ;
  assign n1449 = n1178 & n1180 ;
  assign n1450 = ( ~n1001 & n1448 ) | ( ~n1001 & n1449 ) | ( n1448 & n1449 );
  assign n1451 = n1182 | n1450 ;
  assign n1452 = n984 | n1191 ;
  assign n1453 = n984 & n1191 ;
  assign n1454 = n1452 & ~n1453 ;
  assign n1455 = ( ~n1185 & n1221 ) | ( ~n1185 & n1454 ) | ( n1221 & n1454 );
  assign n1456 = n1165 | n1180 ;
  assign n1457 = ( n978 & n999 ) | ( n978 & ~n1456 ) | ( n999 & ~n1456 );
  assign n1458 = ( n978 & n999 ) | ( n978 & ~n1457 ) | ( n999 & ~n1457 );
  assign n1459 = ( n1456 & n1457 ) | ( n1456 & ~n1458 ) | ( n1457 & ~n1458 );
  assign n1460 = n1455 & ~n1459 ;
  assign n1461 = n1455 & n1459 ;
  assign n1462 = ( n1459 & n1460 ) | ( n1459 & ~n1461 ) | ( n1460 & ~n1461 );
  assign n1463 = n1338 | n1460 ;
  assign n1464 = ( n1460 & ~n1462 ) | ( n1460 & n1463 ) | ( ~n1462 & n1463 );
  assign n1465 = ~n1451 & n1464 ;
  assign n1466 = ~n1451 & n1460 ;
  assign n1467 = ( n1451 & n1462 ) | ( n1451 & ~n1466 ) | ( n1462 & ~n1466 );
  assign n1468 = ( n1447 & ~n1465 ) | ( n1447 & n1467 ) | ( ~n1465 & n1467 );
  assign n1469 = ~n1339 & n1445 ;
  assign n1470 = ~n1342 & n1469 ;
  assign n1471 = ( n1465 & ~n1467 ) | ( n1465 & n1470 ) | ( ~n1467 & n1470 );
  assign n1472 = ~n1441 & n1443 ;
  assign n1473 = n1441 & ~n1443 ;
  assign n1474 = n1472 | n1473 ;
  assign n1475 = n1308 | n1327 ;
  assign n1476 = ~n1328 & n1475 ;
  assign n1477 = n1295 & ~n1303 ;
  assign n1478 = n1304 | n1477 ;
  assign n1479 = n589 | n1356 ;
  assign n1480 = n595 & n1479 ;
  assign n1481 = n576 & n1356 ;
  assign n1482 = n589 & ~n1481 ;
  assign n1483 = n1480 & n1482 ;
  assign n1484 = n1064 & ~n1396 ;
  assign n1485 = n1396 | n1484 ;
  assign n1486 = n516 & ~n1485 ;
  assign n1487 = ~n516 & n1484 ;
  assign n1488 = n599 | n1064 ;
  assign n1489 = n1396 & n1488 ;
  assign n1490 = n1487 | n1489 ;
  assign n1491 = n1486 | n1490 ;
  assign n1492 = n1483 & ~n1491 ;
  assign n1493 = n595 | n1291 ;
  assign n1494 = ~n582 & n1291 ;
  assign n1495 = n1493 & ~n1494 ;
  assign n1496 = ( ~n590 & n1238 ) | ( ~n590 & n1495 ) | ( n1238 & n1495 );
  assign n1497 = ( n576 & n1238 ) | ( n576 & ~n1495 ) | ( n1238 & ~n1495 );
  assign n1498 = n1496 & ~n1497 ;
  assign n1499 = n1492 & n1498 ;
  assign n1500 = n1492 | n1498 ;
  assign n1501 = ~n1499 & n1500 ;
  assign n1502 = n750 & n1206 ;
  assign n1503 = n750 | n1138 ;
  assign n1504 = ( n742 & ~n1207 ) | ( n742 & n1503 ) | ( ~n1207 & n1503 );
  assign n1505 = ( n742 & n1137 ) | ( n742 & ~n1503 ) | ( n1137 & ~n1503 );
  assign n1506 = n1504 & ~n1505 ;
  assign n1507 = ~n1502 & n1506 ;
  assign n1508 = n969 & n985 ;
  assign n1509 = ~n969 & n987 ;
  assign n1510 = ( n778 & n851 ) | ( n778 & ~n1509 ) | ( n851 & ~n1509 );
  assign n1511 = ( ~n776 & n851 ) | ( ~n776 & n1509 ) | ( n851 & n1509 );
  assign n1512 = n1510 & ~n1511 ;
  assign n1513 = ~n1508 & n1512 ;
  assign n1514 = n767 & n1123 ;
  assign n1515 = n754 & ~n1123 ;
  assign n1516 = ( n524 & n1238 ) | ( n524 & ~n1515 ) | ( n1238 & ~n1515 );
  assign n1517 = ( ~n522 & n1238 ) | ( ~n522 & n1515 ) | ( n1238 & n1515 );
  assign n1518 = n1516 & ~n1517 ;
  assign n1519 = ~n1514 & n1518 ;
  assign n1520 = ( n1507 & n1513 ) | ( n1507 & n1519 ) | ( n1513 & n1519 );
  assign n1521 = n1499 | n1520 ;
  assign n1522 = ( n1499 & n1501 ) | ( n1499 & n1521 ) | ( n1501 & n1521 );
  assign n1523 = ( n1314 & n1326 ) | ( n1314 & ~n1327 ) | ( n1326 & ~n1327 );
  assign n1524 = ( n1320 & ~n1327 ) | ( n1320 & n1523 ) | ( ~n1327 & n1523 );
  assign n1525 = ( ~n1478 & n1522 ) | ( ~n1478 & n1524 ) | ( n1522 & n1524 );
  assign n1526 = n1476 & n1525 ;
  assign n1527 = n1345 & ~n1347 ;
  assign n1528 = ( n1347 & ~n1433 ) | ( n1347 & n1435 ) | ( ~n1433 & n1435 );
  assign n1529 = n1433 & ~n1435 ;
  assign n1530 = ( n1345 & ~n1528 ) | ( n1345 & n1529 ) | ( ~n1528 & n1529 );
  assign n1531 = ( n1433 & n1527 ) | ( n1433 & ~n1530 ) | ( n1527 & ~n1530 );
  assign n1532 = n1476 | n1525 ;
  assign n1533 = ~n1526 & n1532 ;
  assign n1534 = ~n1530 & n1533 ;
  assign n1535 = ~n1435 & n1533 ;
  assign n1536 = ( n1531 & n1534 ) | ( n1531 & n1535 ) | ( n1534 & n1535 );
  assign n1537 = n1526 | n1536 ;
  assign n1538 = ~n1474 & n1537 ;
  assign n1539 = n1474 & ~n1537 ;
  assign n1540 = n1538 | n1539 ;
  assign n1541 = n1530 & ~n1533 ;
  assign n1542 = n1435 & ~n1533 ;
  assign n1543 = ( ~n1531 & n1541 ) | ( ~n1531 & n1542 ) | ( n1541 & n1542 );
  assign n1544 = n1536 | n1543 ;
  assign n1545 = n1412 | n1431 ;
  assign n1546 = ~n1432 & n1545 ;
  assign n1547 = ~n1483 & n1491 ;
  assign n1548 = n1492 | n1547 ;
  assign n1549 = n595 | n1356 ;
  assign n1550 = ~n582 & n1356 ;
  assign n1551 = n1549 & ~n1550 ;
  assign n1552 = ( ~n590 & n1291 ) | ( ~n590 & n1551 ) | ( n1291 & n1551 );
  assign n1553 = ( n576 & n1291 ) | ( n576 & ~n1551 ) | ( n1291 & ~n1551 );
  assign n1554 = n1552 & ~n1553 ;
  assign n1555 = ~n1405 & n1407 ;
  assign n1556 = n1408 | n1555 ;
  assign n1557 = n1554 & ~n1556 ;
  assign n1558 = n587 & n1296 ;
  assign n1559 = ~n587 & n1298 ;
  assign n1560 = ( n761 & n1248 ) | ( n761 & ~n1559 ) | ( n1248 & ~n1559 );
  assign n1561 = ( n761 & ~n1246 ) | ( n761 & n1559 ) | ( ~n1246 & n1559 );
  assign n1562 = n1560 & ~n1561 ;
  assign n1563 = ~n1558 & n1562 ;
  assign n1564 = ~n1556 & n1563 ;
  assign n1565 = ( ~n1548 & n1557 ) | ( ~n1548 & n1564 ) | ( n1557 & n1564 );
  assign n1566 = ~n1554 & n1556 ;
  assign n1567 = n1556 & ~n1563 ;
  assign n1568 = ( n1548 & n1566 ) | ( n1548 & n1567 ) | ( n1566 & n1567 );
  assign n1569 = n1565 | n1568 ;
  assign n1570 = ( n1418 & n1430 ) | ( n1418 & ~n1431 ) | ( n1430 & ~n1431 );
  assign n1571 = ( n1424 & ~n1431 ) | ( n1424 & n1570 ) | ( ~n1431 & n1570 );
  assign n1572 = n1565 | n1571 ;
  assign n1573 = ( n1565 & ~n1569 ) | ( n1565 & n1572 ) | ( ~n1569 & n1572 );
  assign n1574 = n1546 & n1573 ;
  assign n1575 = n1546 | n1573 ;
  assign n1576 = ~n1574 & n1575 ;
  assign n1577 = ( n1478 & n1522 ) | ( n1478 & ~n1524 ) | ( n1522 & ~n1524 );
  assign n1578 = ( ~n1522 & n1525 ) | ( ~n1522 & n1577 ) | ( n1525 & n1577 );
  assign n1579 = n1576 & ~n1578 ;
  assign n1580 = n1574 | n1579 ;
  assign n1581 = ~n1576 & n1578 ;
  assign n1582 = n1579 | n1581 ;
  assign n1583 = n1501 & n1520 ;
  assign n1584 = n1501 | n1520 ;
  assign n1585 = ~n1583 & n1584 ;
  assign n1586 = n761 & n1296 ;
  assign n1587 = ~n761 & n1298 ;
  assign n1588 = ( n750 & n1248 ) | ( n750 & ~n1587 ) | ( n1248 & ~n1587 );
  assign n1589 = ( n750 & ~n1246 ) | ( n750 & n1587 ) | ( ~n1246 & n1587 );
  assign n1590 = n1588 & ~n1589 ;
  assign n1591 = ~n1586 & n1590 ;
  assign n1592 = n587 | n1064 ;
  assign n1593 = n1396 & n1592 ;
  assign n1594 = ( n599 & n1064 ) | ( n599 & n1396 ) | ( n1064 & n1396 );
  assign n1595 = ( n1488 & n1593 ) | ( n1488 & ~n1594 ) | ( n1593 & ~n1594 );
  assign n1596 = n767 & n1238 ;
  assign n1597 = n754 & ~n1238 ;
  assign n1598 = ( n524 & n1291 ) | ( n524 & ~n1597 ) | ( n1291 & ~n1597 );
  assign n1599 = ( ~n522 & n1291 ) | ( ~n522 & n1597 ) | ( n1291 & n1597 );
  assign n1600 = n1598 & ~n1599 ;
  assign n1601 = ~n1596 & n1600 ;
  assign n1602 = ( n1591 & ~n1595 ) | ( n1591 & n1601 ) | ( ~n1595 & n1601 );
  assign n1603 = n742 & n1206 ;
  assign n1604 = n742 | n1138 ;
  assign n1605 = ( n969 & ~n1207 ) | ( n969 & n1604 ) | ( ~n1207 & n1604 );
  assign n1606 = ( n969 & n1137 ) | ( n969 & ~n1604 ) | ( n1137 & ~n1604 );
  assign n1607 = n1605 & ~n1606 ;
  assign n1608 = ~n1603 & n1607 ;
  assign n1609 = n851 & n985 ;
  assign n1610 = ~n851 & n987 ;
  assign n1611 = ( n778 & n1123 ) | ( n778 & ~n1610 ) | ( n1123 & ~n1610 );
  assign n1612 = ( ~n776 & n1123 ) | ( ~n776 & n1610 ) | ( n1123 & n1610 );
  assign n1613 = n1611 & ~n1612 ;
  assign n1614 = ~n1609 & n1613 ;
  assign n1615 = n761 | n1064 ;
  assign n1616 = n1396 & n1615 ;
  assign n1617 = ( n587 & n1064 ) | ( n587 & n1396 ) | ( n1064 & n1396 );
  assign n1618 = ( n1592 & n1616 ) | ( n1592 & ~n1617 ) | ( n1616 & ~n1617 );
  assign n1619 = n767 & n1356 ;
  assign n1620 = n510 & ~n1619 ;
  assign n1621 = ~n1618 & n1620 ;
  assign n1622 = ( n1608 & n1614 ) | ( n1608 & n1621 ) | ( n1614 & n1621 );
  assign n1623 = ( n1507 & n1519 ) | ( n1507 & ~n1520 ) | ( n1519 & ~n1520 );
  assign n1624 = ( n1513 & ~n1520 ) | ( n1513 & n1623 ) | ( ~n1520 & n1623 );
  assign n1625 = ( n1602 & n1622 ) | ( n1602 & n1624 ) | ( n1622 & n1624 );
  assign n1626 = n1585 & n1625 ;
  assign n1627 = n1585 | n1625 ;
  assign n1628 = ~n1626 & n1627 ;
  assign n1629 = n1568 | n1572 ;
  assign n1630 = n1569 & n1571 ;
  assign n1631 = n1629 & ~n1630 ;
  assign n1632 = ~n1626 & n1631 ;
  assign n1633 = ( n1626 & n1628 ) | ( n1626 & ~n1632 ) | ( n1628 & ~n1632 );
  assign n1634 = ~n1582 & n1633 ;
  assign n1635 = n1628 & ~n1631 ;
  assign n1636 = ~n1628 & n1631 ;
  assign n1637 = n1635 | n1636 ;
  assign n1638 = n742 | n1248 ;
  assign n1639 = n742 & ~n1246 ;
  assign n1640 = n1638 & ~n1639 ;
  assign n1641 = ( n750 & n1296 ) | ( n750 & ~n1640 ) | ( n1296 & ~n1640 );
  assign n1642 = ( n750 & ~n1298 ) | ( n750 & n1640 ) | ( ~n1298 & n1640 );
  assign n1643 = ~n1641 & n1642 ;
  assign n1644 = n778 | n1238 ;
  assign n1645 = ~n776 & n1238 ;
  assign n1646 = n1644 & ~n1645 ;
  assign n1647 = ( ~n987 & n1123 ) | ( ~n987 & n1646 ) | ( n1123 & n1646 );
  assign n1648 = ( n985 & n1123 ) | ( n985 & ~n1646 ) | ( n1123 & ~n1646 );
  assign n1649 = n1647 & ~n1648 ;
  assign n1650 = ~n851 & n1207 ;
  assign n1651 = n851 & n1137 ;
  assign n1652 = n1650 | n1651 ;
  assign n1653 = ( n969 & n1138 ) | ( n969 & ~n1652 ) | ( n1138 & ~n1652 );
  assign n1654 = ( n969 & n1206 ) | ( n969 & n1652 ) | ( n1206 & n1652 );
  assign n1655 = n1653 & ~n1654 ;
  assign n1656 = ( n1643 & n1649 ) | ( n1643 & n1655 ) | ( n1649 & n1655 );
  assign n1657 = ~n1483 & n1656 ;
  assign n1658 = ~n589 & n1481 ;
  assign n1659 = ( n589 & n1480 ) | ( n589 & ~n1658 ) | ( n1480 & ~n1658 );
  assign n1660 = n1657 & n1659 ;
  assign n1661 = n1483 | n1659 ;
  assign n1662 = ( n1483 & n1657 ) | ( n1483 & n1661 ) | ( n1657 & n1661 );
  assign n1663 = n1659 & ~n1662 ;
  assign n1666 = ( n1608 & n1621 ) | ( n1608 & ~n1622 ) | ( n1621 & ~n1622 );
  assign n1667 = ( n1614 & ~n1622 ) | ( n1614 & n1666 ) | ( ~n1622 & n1666 );
  assign n1664 = n1656 & ~n1659 ;
  assign n1665 = ( n1656 & ~n1657 ) | ( n1656 & n1664 ) | ( ~n1657 & n1664 );
  assign n1668 = n1665 & n1667 ;
  assign n1669 = ( n1663 & n1667 ) | ( n1663 & n1668 ) | ( n1667 & n1668 );
  assign n1670 = n1660 | n1669 ;
  assign n1671 = ( ~n1602 & n1622 ) | ( ~n1602 & n1624 ) | ( n1622 & n1624 );
  assign n1672 = ( n1602 & ~n1622 ) | ( n1602 & n1671 ) | ( ~n1622 & n1671 );
  assign n1673 = ( ~n1624 & n1671 ) | ( ~n1624 & n1672 ) | ( n1671 & n1672 );
  assign n1674 = ( ~n1548 & n1554 ) | ( ~n1548 & n1563 ) | ( n1554 & n1563 );
  assign n1675 = ( n1548 & ~n1554 ) | ( n1548 & n1674 ) | ( ~n1554 & n1674 );
  assign n1676 = ( ~n1563 & n1674 ) | ( ~n1563 & n1675 ) | ( n1674 & n1675 );
  assign n1677 = ( n1670 & n1673 ) | ( n1670 & ~n1676 ) | ( n1673 & ~n1676 );
  assign n1678 = ~n1637 & n1677 ;
  assign n1679 = n1637 & ~n1677 ;
  assign n1680 = n1678 | n1679 ;
  assign n1681 = n1670 & n1676 ;
  assign n1682 = n1670 | n1676 ;
  assign n1683 = ~n1681 & n1682 ;
  assign n1684 = n1673 & ~n1683 ;
  assign n1688 = n1618 & ~n1620 ;
  assign n1689 = n1621 | n1688 ;
  assign n1690 = n767 & n1291 ;
  assign n1691 = n754 & ~n1291 ;
  assign n1692 = ( n524 & n1356 ) | ( n524 & ~n1691 ) | ( n1356 & ~n1691 );
  assign n1693 = ( ~n522 & n1356 ) | ( ~n522 & n1691 ) | ( n1356 & n1691 );
  assign n1694 = n1692 & ~n1693 ;
  assign n1695 = ~n1690 & n1694 ;
  assign n1696 = ~n1689 & n1695 ;
  assign n1697 = n969 | n1248 ;
  assign n1698 = n969 & ~n1246 ;
  assign n1699 = n1697 & ~n1698 ;
  assign n1700 = ( n742 & n1296 ) | ( n742 & ~n1699 ) | ( n1296 & ~n1699 );
  assign n1701 = ( n742 & ~n1298 ) | ( n742 & n1699 ) | ( ~n1298 & n1699 );
  assign n1702 = ~n1700 & n1701 ;
  assign n1703 = ~n1123 & n1207 ;
  assign n1704 = n1123 & n1137 ;
  assign n1705 = n1703 | n1704 ;
  assign n1706 = ( n851 & n1138 ) | ( n851 & ~n1705 ) | ( n1138 & ~n1705 );
  assign n1707 = ( n851 & n1206 ) | ( n851 & n1705 ) | ( n1206 & n1705 );
  assign n1708 = n1706 & ~n1707 ;
  assign n1709 = n750 | n1064 ;
  assign n1710 = n1396 & n1709 ;
  assign n1711 = ( n761 & n1064 ) | ( n761 & n1396 ) | ( n1064 & n1396 );
  assign n1712 = ( n1615 & n1710 ) | ( n1615 & ~n1711 ) | ( n1710 & ~n1711 );
  assign n1713 = ( n1702 & n1708 ) | ( n1702 & ~n1712 ) | ( n1708 & ~n1712 );
  assign n1714 = n1695 & ~n1696 ;
  assign n1715 = ( n1689 & n1696 ) | ( n1689 & ~n1714 ) | ( n1696 & ~n1714 );
  assign n1716 = n1713 & ~n1715 ;
  assign n1717 = n1696 | n1716 ;
  assign n1685 = ( n1591 & n1595 ) | ( n1591 & n1601 ) | ( n1595 & n1601 );
  assign n1686 = ( n1595 & n1601 ) | ( n1595 & ~n1685 ) | ( n1601 & ~n1685 );
  assign n1687 = ( n1591 & ~n1685 ) | ( n1591 & n1686 ) | ( ~n1685 & n1686 );
  assign n1718 = ~n1687 & n1717 ;
  assign n1719 = n1717 & ~n1718 ;
  assign n1720 = n1687 | n1718 ;
  assign n1721 = ~n1719 & n1720 ;
  assign n1722 = n1665 | n1667 ;
  assign n1723 = n1663 | n1722 ;
  assign n1724 = ~n1669 & n1723 ;
  assign n1725 = ~n1721 & n1724 ;
  assign n1726 = n1721 & ~n1724 ;
  assign n1727 = n1725 | n1726 ;
  assign n1728 = ( n1702 & n1708 ) | ( n1702 & ~n1713 ) | ( n1708 & ~n1713 );
  assign n1729 = n851 | n1248 ;
  assign n1730 = n851 & ~n1246 ;
  assign n1731 = n1729 & ~n1730 ;
  assign n1732 = ( n969 & n1296 ) | ( n969 & ~n1731 ) | ( n1296 & ~n1731 );
  assign n1733 = ( n969 & ~n1298 ) | ( n969 & n1731 ) | ( ~n1298 & n1731 );
  assign n1734 = ~n1732 & n1733 ;
  assign n1735 = n1207 & ~n1238 ;
  assign n1736 = n1137 & n1238 ;
  assign n1737 = n1735 | n1736 ;
  assign n1738 = ( n1123 & n1138 ) | ( n1123 & ~n1737 ) | ( n1138 & ~n1737 );
  assign n1739 = ( n1123 & n1206 ) | ( n1123 & n1737 ) | ( n1206 & n1737 );
  assign n1740 = n1738 & ~n1739 ;
  assign n1741 = n778 | n1356 ;
  assign n1742 = ~n776 & n1356 ;
  assign n1743 = n1741 & ~n1742 ;
  assign n1744 = ( ~n987 & n1291 ) | ( ~n987 & n1743 ) | ( n1291 & n1743 );
  assign n1745 = ( n985 & n1291 ) | ( n985 & ~n1743 ) | ( n1291 & ~n1743 );
  assign n1746 = n1744 & ~n1745 ;
  assign n1747 = ( n1734 & n1740 ) | ( n1734 & n1746 ) | ( n1740 & n1746 );
  assign n1748 = ~n1713 & n1747 ;
  assign n1749 = ~n1712 & n1747 ;
  assign n1750 = ( n1728 & n1748 ) | ( n1728 & n1749 ) | ( n1748 & n1749 );
  assign n1751 = ( n1712 & n1713 ) | ( n1712 & ~n1728 ) | ( n1713 & ~n1728 );
  assign n1752 = n1750 | n1751 ;
  assign n1753 = n778 | n1291 ;
  assign n1754 = ~n776 & n1291 ;
  assign n1755 = n1753 & ~n1754 ;
  assign n1756 = ( ~n987 & n1238 ) | ( ~n987 & n1755 ) | ( n1238 & n1755 );
  assign n1757 = ( n985 & n1238 ) | ( n985 & ~n1755 ) | ( n1238 & ~n1755 );
  assign n1758 = n1756 & ~n1757 ;
  assign n1759 = n521 & n1356 ;
  assign n1760 = n737 | n1356 ;
  assign n1761 = n778 & n1760 ;
  assign n1762 = n985 & n1356 ;
  assign n1763 = n737 & ~n1762 ;
  assign n1764 = n1761 & n1763 ;
  assign n1765 = n742 | n1064 ;
  assign n1766 = n1396 & n1765 ;
  assign n1767 = ( n750 & n1064 ) | ( n750 & n1396 ) | ( n1064 & n1396 );
  assign n1768 = ( n1709 & n1766 ) | ( n1709 & ~n1767 ) | ( n1766 & ~n1767 );
  assign n1769 = n1764 & ~n1768 ;
  assign n1770 = ( n1758 & n1759 ) | ( n1758 & ~n1769 ) | ( n1759 & ~n1769 );
  assign n1771 = ( ~n1759 & n1769 ) | ( ~n1759 & n1770 ) | ( n1769 & n1770 );
  assign n1772 = ( ~n1758 & n1770 ) | ( ~n1758 & n1771 ) | ( n1770 & n1771 );
  assign n1773 = n1713 & n1747 ;
  assign n1774 = n1712 & n1747 ;
  assign n1775 = ( ~n1728 & n1773 ) | ( ~n1728 & n1774 ) | ( n1773 & n1774 );
  assign n1776 = n1772 & n1775 ;
  assign n1777 = ( ~n1752 & n1772 ) | ( ~n1752 & n1776 ) | ( n1772 & n1776 );
  assign n1778 = n1750 | n1777 ;
  assign n1779 = ( n1643 & n1649 ) | ( n1643 & ~n1655 ) | ( n1649 & ~n1655 );
  assign n1780 = ( n1643 & n1649 ) | ( n1643 & ~n1779 ) | ( n1649 & ~n1779 );
  assign n1781 = ( n1758 & n1759 ) | ( n1758 & n1769 ) | ( n1759 & n1769 );
  assign n1782 = n1779 & n1781 ;
  assign n1783 = n1655 & n1781 ;
  assign n1784 = ( ~n1780 & n1782 ) | ( ~n1780 & n1783 ) | ( n1782 & n1783 );
  assign n1785 = n1779 | n1781 ;
  assign n1786 = n1655 | n1781 ;
  assign n1787 = ( ~n1780 & n1785 ) | ( ~n1780 & n1786 ) | ( n1785 & n1786 );
  assign n1788 = ~n1784 & n1787 ;
  assign n1789 = ~n1713 & n1715 ;
  assign n1790 = n1716 | n1789 ;
  assign n1791 = ~n1788 & n1790 ;
  assign n1792 = n1788 & ~n1790 ;
  assign n1793 = n1791 | n1792 ;
  assign n1794 = ( n1734 & n1740 ) | ( n1734 & ~n1746 ) | ( n1740 & ~n1746 );
  assign n1795 = ( n1734 & n1740 ) | ( n1734 & ~n1794 ) | ( n1740 & ~n1794 );
  assign n1796 = ( n1746 & n1794 ) | ( n1746 & ~n1795 ) | ( n1794 & ~n1795 );
  assign n1797 = n963 & ~n1207 ;
  assign n1798 = ( n1206 & n1356 ) | ( n1206 & ~n1797 ) | ( n1356 & ~n1797 );
  assign n1799 = n1797 & ~n1798 ;
  assign n1800 = n851 | n1064 ;
  assign n1801 = n1396 & n1800 ;
  assign n1802 = n969 | n1064 ;
  assign n1803 = ( n969 & n1064 ) | ( n969 & n1396 ) | ( n1064 & n1396 );
  assign n1804 = ( n1801 & n1802 ) | ( n1801 & ~n1803 ) | ( n1802 & ~n1803 );
  assign n1805 = n1799 & ~n1804 ;
  assign n1806 = ~n1799 & n1804 ;
  assign n1807 = n1805 | n1806 ;
  assign n1808 = n1238 | n1248 ;
  assign n1809 = n1238 & ~n1246 ;
  assign n1810 = n1808 & ~n1809 ;
  assign n1811 = ( n1123 & n1296 ) | ( n1123 & ~n1810 ) | ( n1296 & ~n1810 );
  assign n1812 = ( n1123 & ~n1298 ) | ( n1123 & n1810 ) | ( ~n1298 & n1810 );
  assign n1813 = ~n1811 & n1812 ;
  assign n1814 = n1207 & ~n1356 ;
  assign n1815 = n1137 & n1356 ;
  assign n1816 = n1814 | n1815 ;
  assign n1817 = ( n1138 & n1291 ) | ( n1138 & ~n1816 ) | ( n1291 & ~n1816 );
  assign n1818 = ( n1206 & n1291 ) | ( n1206 & n1816 ) | ( n1291 & n1816 );
  assign n1819 = n1817 & ~n1818 ;
  assign n1820 = ( ~n1807 & n1813 ) | ( ~n1807 & n1819 ) | ( n1813 & n1819 );
  assign n1821 = ( n1813 & n1819 ) | ( n1813 & ~n1820 ) | ( n1819 & ~n1820 );
  assign n1822 = ( n1807 & n1820 ) | ( n1807 & ~n1821 ) | ( n1820 & ~n1821 );
  assign n1823 = n1248 | n1291 ;
  assign n1824 = ~n1246 & n1291 ;
  assign n1825 = n1823 & ~n1824 ;
  assign n1826 = ( n1238 & n1296 ) | ( n1238 & ~n1825 ) | ( n1296 & ~n1825 );
  assign n1827 = ( n1238 & ~n1298 ) | ( n1238 & n1825 ) | ( ~n1298 & n1825 );
  assign n1828 = ~n1826 & n1827 ;
  assign n1829 = n1296 & n1356 ;
  assign n1830 = n1298 & n1356 ;
  assign n1831 = ( n1116 & ~n1829 ) | ( n1116 & n1830 ) | ( ~n1829 & n1830 );
  assign n1832 = n1123 & ~n1396 ;
  assign n1833 = n1238 & n1396 ;
  assign n1834 = ( n1064 & ~n1832 ) | ( n1064 & n1833 ) | ( ~n1832 & n1833 );
  assign n1835 = ~n1484 & n1832 ;
  assign n1836 = n1834 | n1835 ;
  assign n1837 = n1116 & ~n1836 ;
  assign n1838 = n1831 & n1837 ;
  assign n1839 = ~n851 & n1484 ;
  assign n1840 = n1064 | n1123 ;
  assign n1841 = n1396 & n1840 ;
  assign n1842 = n1839 | n1841 ;
  assign n1843 = n851 & ~n1396 ;
  assign n1844 = ~n1484 & n1843 ;
  assign n1845 = n1842 | n1844 ;
  assign n1846 = ( n1828 & n1838 ) | ( n1828 & ~n1845 ) | ( n1838 & ~n1845 );
  assign n1847 = ( n1828 & ~n1838 ) | ( n1828 & n1845 ) | ( ~n1838 & n1845 );
  assign n1848 = ( ~n1828 & n1846 ) | ( ~n1828 & n1847 ) | ( n1846 & n1847 );
  assign n1849 = ~n1116 & n1836 ;
  assign n1850 = ( ~n1831 & n1836 ) | ( ~n1831 & n1849 ) | ( n1836 & n1849 );
  assign n1851 = n1838 | n1850 ;
  assign n1859 = ~n1136 & n1356 ;
  assign n1852 = n1064 | n1291 ;
  assign n1853 = n1396 & n1852 ;
  assign n1854 = ( n1238 & ~n1485 ) | ( n1238 & n1853 ) | ( ~n1485 & n1853 );
  assign n1855 = ( ~n1238 & n1484 ) | ( ~n1238 & n1853 ) | ( n1484 & n1853 );
  assign n1856 = n1854 | n1855 ;
  assign n1857 = ( ~n1064 & n1243 ) | ( ~n1064 & n1356 ) | ( n1243 & n1356 );
  assign n1858 = ( n1114 & n1243 ) | ( n1114 & n1857 ) | ( n1243 & n1857 );
  assign n1860 = n1858 | n1859 ;
  assign n1861 = n1064 | n1356 ;
  assign n1862 = n1291 & ~n1396 ;
  assign n1863 = n1861 | n1862 ;
  assign n1864 = ~n1859 & n1863 ;
  assign n1865 = ( n1856 & ~n1860 ) | ( n1856 & n1864 ) | ( ~n1860 & n1864 );
  assign n1866 = ( n1851 & ~n1859 ) | ( n1851 & n1865 ) | ( ~n1859 & n1865 );
  assign n1867 = n1848 | n1866 ;
  assign n1868 = ~n1246 & n1356 ;
  assign n1869 = ( n1291 & n1296 ) | ( n1291 & n1868 ) | ( n1296 & n1868 );
  assign n1870 = ( ~n1291 & n1298 ) | ( ~n1291 & n1868 ) | ( n1298 & n1868 );
  assign n1871 = n1869 | n1870 ;
  assign n1872 = n1248 | n1356 ;
  assign n1873 = ~n1871 & n1872 ;
  assign n1874 = ( n1856 & ~n1858 ) | ( n1856 & n1863 ) | ( ~n1858 & n1863 );
  assign n1875 = n1872 & ~n1874 ;
  assign n1876 = ~n1871 & n1875 ;
  assign n1877 = ( ~n1851 & n1873 ) | ( ~n1851 & n1876 ) | ( n1873 & n1876 );
  assign n1878 = ( n1848 & n1867 ) | ( n1848 & ~n1877 ) | ( n1867 & ~n1877 );
  assign n1879 = ( n1851 & ~n1873 ) | ( n1851 & n1874 ) | ( ~n1873 & n1874 );
  assign n1880 = n1859 & ~n1879 ;
  assign n1881 = ~n1822 & n1880 ;
  assign n1882 = ( n1822 & n1878 ) | ( n1822 & ~n1881 ) | ( n1878 & ~n1881 );
  assign n1883 = ~n737 & n1762 ;
  assign n1884 = ( n737 & n1761 ) | ( n737 & ~n1883 ) | ( n1761 & ~n1883 );
  assign n1885 = ~n1764 & n1884 ;
  assign n1886 = ( n1805 & ~n1807 ) | ( n1805 & n1885 ) | ( ~n1807 & n1885 );
  assign n1887 = ( n1805 & n1819 ) | ( n1805 & n1885 ) | ( n1819 & n1885 );
  assign n1888 = ( n1813 & n1886 ) | ( n1813 & n1887 ) | ( n1886 & n1887 );
  assign n1889 = ( n1820 & n1885 ) | ( n1820 & ~n1888 ) | ( n1885 & ~n1888 );
  assign n1890 = ( n1805 & ~n1888 ) | ( n1805 & n1889 ) | ( ~n1888 & n1889 );
  assign n1891 = n1882 & ~n1890 ;
  assign n1892 = ~n742 & n1484 ;
  assign n1893 = n1396 & n1802 ;
  assign n1894 = n1892 | n1893 ;
  assign n1895 = n742 & ~n1396 ;
  assign n1896 = ~n1484 & n1895 ;
  assign n1897 = n1894 | n1896 ;
  assign n1898 = n1123 | n1248 ;
  assign n1899 = n1123 & ~n1246 ;
  assign n1900 = n1898 & ~n1899 ;
  assign n1901 = ( n851 & n1296 ) | ( n851 & ~n1900 ) | ( n1296 & ~n1900 );
  assign n1902 = ( n851 & ~n1298 ) | ( n851 & n1900 ) | ( ~n1298 & n1900 );
  assign n1903 = ~n1901 & n1902 ;
  assign n1904 = n1207 & ~n1291 ;
  assign n1905 = n1137 & n1291 ;
  assign n1906 = n1904 | n1905 ;
  assign n1907 = ( n1138 & n1238 ) | ( n1138 & ~n1906 ) | ( n1238 & ~n1906 );
  assign n1908 = ( n1206 & n1238 ) | ( n1206 & n1906 ) | ( n1238 & n1906 );
  assign n1909 = n1907 & ~n1908 ;
  assign n1910 = ( ~n1897 & n1903 ) | ( ~n1897 & n1909 ) | ( n1903 & n1909 );
  assign n1911 = ( n1903 & n1909 ) | ( n1903 & ~n1910 ) | ( n1909 & ~n1910 );
  assign n1912 = ( n1897 & n1910 ) | ( n1897 & ~n1911 ) | ( n1910 & ~n1911 );
  assign n1913 = n1822 & ~n1880 ;
  assign n1914 = n1846 & ~n1848 ;
  assign n1915 = n1846 & n1877 ;
  assign n1916 = ( ~n1867 & n1914 ) | ( ~n1867 & n1915 ) | ( n1914 & n1915 );
  assign n1917 = ( n1846 & ~n1913 ) | ( n1846 & n1916 ) | ( ~n1913 & n1916 );
  assign n1918 = ~n1912 & n1917 ;
  assign n1919 = ( n1891 & n1912 ) | ( n1891 & ~n1918 ) | ( n1912 & ~n1918 );
  assign n1920 = ~n1882 & n1890 ;
  assign n1921 = n1888 | n1917 ;
  assign n1922 = n1888 | n1890 ;
  assign n1923 = ( n1920 & n1921 ) | ( n1920 & n1922 ) | ( n1921 & n1922 );
  assign n1924 = n1919 & ~n1923 ;
  assign n1925 = ~n1764 & n1768 ;
  assign n1926 = n1769 | n1925 ;
  assign n1927 = ~n1909 & n1926 ;
  assign n1928 = n1897 & n1926 ;
  assign n1929 = ( ~n1903 & n1927 ) | ( ~n1903 & n1928 ) | ( n1927 & n1928 );
  assign n1930 = n1926 & ~n1928 ;
  assign n1931 = n1926 & ~n1927 ;
  assign n1932 = ( n1903 & n1930 ) | ( n1903 & n1931 ) | ( n1930 & n1931 );
  assign n1933 = ( n1910 & n1929 ) | ( n1910 & ~n1932 ) | ( n1929 & ~n1932 );
  assign n1934 = ( ~n1796 & n1924 ) | ( ~n1796 & n1933 ) | ( n1924 & n1933 );
  assign n1935 = n1772 | n1775 ;
  assign n1936 = n1752 & ~n1935 ;
  assign n1937 = n1777 | n1936 ;
  assign n1938 = n1888 & n1917 ;
  assign n1939 = n1888 & n1890 ;
  assign n1940 = ( n1920 & n1938 ) | ( n1920 & n1939 ) | ( n1938 & n1939 );
  assign n1941 = ( n1888 & ~n1919 ) | ( n1888 & n1940 ) | ( ~n1919 & n1940 );
  assign n1942 = ( n1794 & n1910 ) | ( n1794 & ~n1926 ) | ( n1910 & ~n1926 );
  assign n1943 = ( n1746 & n1909 ) | ( n1746 & ~n1926 ) | ( n1909 & ~n1926 );
  assign n1944 = ( ~n1746 & n1897 ) | ( ~n1746 & n1926 ) | ( n1897 & n1926 );
  assign n1945 = ( n1903 & n1943 ) | ( n1903 & ~n1944 ) | ( n1943 & ~n1944 );
  assign n1946 = ( ~n1795 & n1942 ) | ( ~n1795 & n1945 ) | ( n1942 & n1945 );
  assign n1947 = ( ~n1937 & n1941 ) | ( ~n1937 & n1946 ) | ( n1941 & n1946 );
  assign n1948 = n1796 & ~n1933 ;
  assign n1949 = ( n1937 & ~n1946 ) | ( n1937 & n1948 ) | ( ~n1946 & n1948 );
  assign n1950 = ( n1934 & ~n1947 ) | ( n1934 & n1949 ) | ( ~n1947 & n1949 );
  assign n1951 = ( ~n1778 & n1793 ) | ( ~n1778 & n1950 ) | ( n1793 & n1950 );
  assign n1952 = n1784 | n1792 ;
  assign n1953 = ~n1951 & n1952 ;
  assign n1954 = n1687 & ~n1953 ;
  assign n1955 = n1717 | n1953 ;
  assign n1956 = ( n1724 & ~n1954 ) | ( n1724 & n1955 ) | ( ~n1954 & n1955 );
  assign n1957 = n1717 | n1952 ;
  assign n1958 = n1951 & ~n1957 ;
  assign n1959 = n1687 & ~n1952 ;
  assign n1960 = n1951 & n1959 ;
  assign n1961 = ( ~n1724 & n1958 ) | ( ~n1724 & n1960 ) | ( n1958 & n1960 );
  assign n1962 = ( n1727 & ~n1956 ) | ( n1727 & n1961 ) | ( ~n1956 & n1961 );
  assign n1963 = ( ~n1673 & n1683 ) | ( ~n1673 & n1962 ) | ( n1683 & n1962 );
  assign n1964 = ~n1687 & n1952 ;
  assign n1965 = n1717 & n1952 ;
  assign n1966 = ( n1724 & n1964 ) | ( n1724 & n1965 ) | ( n1964 & n1965 );
  assign n1967 = n1687 | n1951 ;
  assign n1968 = n1717 & ~n1951 ;
  assign n1969 = ( n1724 & ~n1967 ) | ( n1724 & n1968 ) | ( ~n1967 & n1968 );
  assign n1970 = ( ~n1727 & n1966 ) | ( ~n1727 & n1969 ) | ( n1966 & n1969 );
  assign n1971 = ( n1684 & n1963 ) | ( n1684 & ~n1970 ) | ( n1963 & ~n1970 );
  assign n1972 = ~n1678 & n1971 ;
  assign n1973 = ( ~n1678 & n1680 ) | ( ~n1678 & n1972 ) | ( n1680 & n1972 );
  assign n1974 = n1582 & ~n1633 ;
  assign n1975 = n1634 | n1974 ;
  assign n1976 = ~n1634 & n1975 ;
  assign n1977 = ( ~n1634 & n1973 ) | ( ~n1634 & n1976 ) | ( n1973 & n1976 );
  assign n1978 = ( n1544 & ~n1580 ) | ( n1544 & n1977 ) | ( ~n1580 & n1977 );
  assign n1979 = ~n1538 & n1978 ;
  assign n1980 = ( ~n1538 & n1540 ) | ( ~n1538 & n1979 ) | ( n1540 & n1979 );
  assign n1981 = ( n1468 & ~n1471 ) | ( n1468 & n1980 ) | ( ~n1471 & n1980 );
  assign n1982 = ~n1182 & n1981 ;
  assign n1983 = ~n1173 & n1175 ;
  assign n1984 = ( n1169 & n1173 ) | ( n1169 & ~n1983 ) | ( n1173 & ~n1983 );
  assign n1985 = ( n842 & n1982 ) | ( n842 & ~n1984 ) | ( n1982 & ~n1984 );
  assign n1986 = ~n798 & n1982 ;
  assign n1987 = n798 | n1984 ;
  assign n1988 = ( n842 & n1986 ) | ( n842 & ~n1987 ) | ( n1986 & ~n1987 );
  assign n1989 = ( n635 & n1985 ) | ( n635 & n1988 ) | ( n1985 & n1988 );
  assign n1990 = ( n834 & ~n835 ) | ( n834 & n1989 ) | ( ~n835 & n1989 );
  assign n1991 = n810 & n817 ;
  assign n1992 = n812 & n1991 ;
  assign n1993 = ( n818 & ~n819 ) | ( n818 & n1992 ) | ( ~n819 & n1992 );
  assign n1994 = ( n818 & n823 ) | ( n818 & n1993 ) | ( n823 & n1993 );
  assign n1995 = ( ~n611 & n818 ) | ( ~n611 & n1993 ) | ( n818 & n1993 );
  assign n1996 = ( ~n614 & n1994 ) | ( ~n614 & n1995 ) | ( n1994 & n1995 );
  assign n1997 = n820 & ~n826 ;
  assign n1998 = n826 & n1996 ;
  assign n1999 = ( n611 & n614 ) | ( n611 & ~n823 ) | ( n614 & ~n823 );
  assign n2000 = n1996 & n1999 ;
  assign n2001 = ( ~n1997 & n1998 ) | ( ~n1997 & n2000 ) | ( n1998 & n2000 );
  assign n2002 = ( n801 & n1996 ) | ( n801 & n2001 ) | ( n1996 & n2001 );
  assign n2003 = ( ~n799 & n1996 ) | ( ~n799 & n2001 ) | ( n1996 & n2001 );
  assign n2004 = ( n1989 & n2002 ) | ( n1989 & n2003 ) | ( n2002 & n2003 );
  assign n2005 = n1990 & ~n2004 ;
  assign n2006 = n516 & ~n599 ;
  assign n2007 = ~n516 & n599 ;
  assign n2008 = n2006 | n2007 ;
  assign n2009 = n310 & n2008 ;
  assign n2010 = ( n589 & n2005 ) | ( n589 & n2009 ) | ( n2005 & n2009 );
  assign n2011 = ( n589 & ~n2005 ) | ( n589 & n2009 ) | ( ~n2005 & n2009 );
  assign n2012 = ( n2005 & ~n2010 ) | ( n2005 & n2011 ) | ( ~n2010 & n2011 );
  assign n2013 = n151 | n305 ;
  assign n2014 = n214 | n290 ;
  assign n2015 = n2013 | n2014 ;
  assign n2016 = n346 | n394 ;
  assign n2017 = n2015 | n2016 ;
  assign n2018 = n185 | n293 ;
  assign n2019 = n267 | n2018 ;
  assign n2020 = n198 | n2019 ;
  assign n2021 = n549 | n2020 ;
  assign n2022 = n101 | n200 ;
  assign n2023 = n154 | n1067 ;
  assign n2024 = n183 | n313 ;
  assign n2025 = n146 | n333 ;
  assign n2026 = n2024 | n2025 ;
  assign n2027 = n385 | n2026 ;
  assign n2028 = n2023 | n2027 ;
  assign n2029 = n292 | n444 ;
  assign n2030 = n271 | n2029 ;
  assign n2031 = n315 | n2030 ;
  assign n2032 = n311 | n2031 ;
  assign n2033 = n2028 | n2032 ;
  assign n2034 = n460 | n2033 ;
  assign n2035 = n279 | n2034 ;
  assign n2036 = n332 | n2035 ;
  assign n2037 = n180 | n241 ;
  assign n2038 = n2036 | n2037 ;
  assign n2039 = n2022 | n2038 ;
  assign n2040 = n2021 | n2039 ;
  assign n2041 = n422 | n2040 ;
  assign n2042 = n898 & ~n2041 ;
  assign n2043 = ~n2017 & n2042 ;
  assign n2044 = ~n859 & n2043 ;
  assign n2045 = n282 | n1042 ;
  assign n2046 = n177 | n2045 ;
  assign n2047 = n2044 & ~n2046 ;
  assign n2048 = n2012 | n2047 ;
  assign n2049 = n2012 & n2047 ;
  assign n2050 = n2048 & ~n2049 ;
  assign n2051 = n394 | n423 ;
  assign n2052 = n384 | n684 ;
  assign n2053 = n864 | n2052 ;
  assign n2054 = n882 | n2053 ;
  assign n2055 = n418 | n2054 ;
  assign n2056 = ( n344 & ~n2051 ) | ( n344 & n2055 ) | ( ~n2051 & n2055 );
  assign n2057 = n2051 | n2056 ;
  assign n2058 = n163 | n1044 ;
  assign n2059 = n2057 | n2058 ;
  assign n2060 = n1375 | n2059 ;
  assign n2061 = n185 | n265 ;
  assign n2062 = n292 | n2061 ;
  assign n2063 = n206 | n640 ;
  assign n2064 = n2062 | n2063 ;
  assign n2065 = n313 | n2064 ;
  assign n2066 = n2060 | n2065 ;
  assign n2067 = n366 | n2066 ;
  assign n2068 = n462 | n2067 ;
  assign n2069 = n203 | n2068 ;
  assign n2070 = n899 | n2069 ;
  assign n2071 = n436 | n2070 ;
  assign n2072 = n383 | n2071 ;
  assign n2073 = n311 | n2072 ;
  assign n2074 = n2047 & ~n2073 ;
  assign n2075 = ( n2012 & ~n2073 ) | ( n2012 & n2074 ) | ( ~n2073 & n2074 );
  assign n2076 = ( n635 & ~n798 ) | ( n635 & n1985 ) | ( ~n798 & n1985 );
  assign n2077 = ( n826 & ~n1997 ) | ( n826 & n1999 ) | ( ~n1997 & n1999 );
  assign n2078 = n2076 | n2077 ;
  assign n2079 = n177 | n343 ;
  assign n2080 = n190 | n2079 ;
  assign n2081 = n284 | n647 ;
  assign n2082 = n203 | n2081 ;
  assign n2083 = n142 | n2082 ;
  assign n2084 = n235 | n2083 ;
  assign n2085 = n126 | n2084 ;
  assign n2086 = n245 | n2085 ;
  assign n2087 = n182 | n658 ;
  assign n2088 = n291 | n2087 ;
  assign n2089 = n2086 | n2088 ;
  assign n2090 = n700 | n2089 ;
  assign n2091 = n129 | n151 ;
  assign n2092 = n394 | n552 ;
  assign n2093 = n2091 | n2092 ;
  assign n2094 = n161 | n2093 ;
  assign n2095 = n272 | n2094 ;
  assign n2096 = n685 | n2095 ;
  assign n2097 = n213 | n277 ;
  assign n2098 = n556 | n2097 ;
  assign n2099 = n2096 | n2098 ;
  assign n2100 = n120 | n143 ;
  assign n2101 = n240 | n2100 ;
  assign n2102 = n2099 | n2101 ;
  assign n2103 = n200 | n236 ;
  assign n2104 = n271 | n2103 ;
  assign n2105 = n321 | n488 ;
  assign n2106 = n2104 | n2105 ;
  assign n2107 = n215 | n417 ;
  assign n2108 = n154 | n2107 ;
  assign n2109 = n109 | n2108 ;
  assign n2110 = n160 | n1044 ;
  assign n2111 = n2109 | n2110 ;
  assign n2112 = n2106 | n2111 ;
  assign n2113 = n683 | n927 ;
  assign n2114 = n400 | n2113 ;
  assign n2115 = n2112 | n2114 ;
  assign n2116 = n2102 | n2115 ;
  assign n2117 = n2090 | n2116 ;
  assign n2118 = n2080 | n2117 ;
  assign n2119 = n305 | n2118 ;
  assign n2120 = n281 | n2119 ;
  assign n2121 = n150 | n2120 ;
  assign n2122 = n112 | n2121 ;
  assign n2123 = n146 | n2122 ;
  assign n2124 = n384 | n2123 ;
  assign n2125 = ( n2077 & ~n2078 ) | ( n2077 & n2124 ) | ( ~n2078 & n2124 );
  assign n2126 = ( n2076 & ~n2078 ) | ( n2076 & n2125 ) | ( ~n2078 & n2125 );
  assign n2127 = n920 | n921 ;
  assign n2128 = n463 | n642 ;
  assign n2129 = n855 | n2128 ;
  assign n2130 = n155 | n2129 ;
  assign n2131 = n375 | n2130 ;
  assign n2132 = n722 | n2131 ;
  assign n2133 = n2127 | n2132 ;
  assign n2134 = n393 | n2133 ;
  assign n2135 = n1057 | n2134 ;
  assign n2136 = n142 | n2135 ;
  assign n2137 = n109 | n2136 ;
  assign n2138 = n552 | n2137 ;
  assign n2139 = n346 | n2138 ;
  assign n2140 = n96 | n2139 ;
  assign n2141 = n801 | n1985 ;
  assign n2142 = n801 & n1985 ;
  assign n2143 = n2141 & ~n2142 ;
  assign n2144 = n638 & ~n1984 ;
  assign n2145 = ( ~n638 & n1984 ) | ( ~n638 & n2144 ) | ( n1984 & n2144 );
  assign n2146 = n2144 | n2145 ;
  assign n2147 = n839 & ~n1982 ;
  assign n2148 = ~n839 & n1982 ;
  assign n2149 = ( n839 & ~n1982 ) | ( n839 & n1984 ) | ( ~n1982 & n1984 );
  assign n2150 = ( n638 & n2148 ) | ( n638 & ~n2149 ) | ( n2148 & ~n2149 );
  assign n2151 = ( n2145 & ~n2147 ) | ( n2145 & n2150 ) | ( ~n2147 & n2150 );
  assign n2152 = ( ~n839 & n1982 ) | ( ~n839 & n1984 ) | ( n1982 & n1984 );
  assign n2153 = ( n638 & n2147 ) | ( n638 & ~n2152 ) | ( n2147 & ~n2152 );
  assign n2154 = ( n2145 & ~n2148 ) | ( n2145 & n2153 ) | ( ~n2148 & n2153 );
  assign n2155 = ( ~n2146 & n2151 ) | ( ~n2146 & n2154 ) | ( n2151 & n2154 );
  assign n2156 = n127 | n436 ;
  assign n2157 = n96 | n2156 ;
  assign n2158 = n345 | n384 ;
  assign n2159 = n214 | n2013 ;
  assign n2160 = n321 | n2159 ;
  assign n2161 = n2104 | n2160 ;
  assign n2162 = n153 | n494 ;
  assign n2163 = n659 | n2162 ;
  assign n2164 = n2161 | n2163 ;
  assign n2165 = n375 | n2080 ;
  assign n2166 = n444 | n2165 ;
  assign n2167 = n2164 | n2166 ;
  assign n2168 = n260 | n286 ;
  assign n2169 = n191 | n2168 ;
  assign n2170 = n556 | n2169 ;
  assign n2171 = n2167 | n2170 ;
  assign n2172 = n181 | n2171 ;
  assign n2173 = n2158 | n2172 ;
  assign n2174 = n553 | n2173 ;
  assign n2175 = n1365 | n2174 ;
  assign n2176 = n2157 | n2175 ;
  assign n2177 = n234 | n264 ;
  assign n2178 = n169 | n2177 ;
  assign n2179 = n294 | n2178 ;
  assign n2180 = n318 | n2179 ;
  assign n2181 = n283 | n2180 ;
  assign n2182 = n185 | n2181 ;
  assign n2183 = n224 | n2182 ;
  assign n2184 = n459 | n2183 ;
  assign n2185 = n549 | n2184 ;
  assign n2186 = n146 | n2185 ;
  assign n2187 = n246 | n2186 ;
  assign n2188 = n898 & ~n2086 ;
  assign n2189 = ~n2187 & n2188 ;
  assign n2190 = ~n2176 & n2189 ;
  assign n2191 = n206 | n222 ;
  assign n2192 = n225 | n2191 ;
  assign n2193 = n2190 & ~n2192 ;
  assign n2194 = ~n323 & n2193 ;
  assign n2195 = ~n277 & n2194 ;
  assign n2196 = ~n334 & n2195 ;
  assign n2197 = ~n287 & n2196 ;
  assign n2198 = ~n1460 & n1462 ;
  assign n2199 = ( n1464 & n1470 ) | ( n1464 & ~n2198 ) | ( n1470 & ~n2198 );
  assign n2200 = n1451 & ~n2199 ;
  assign n2201 = ( n1447 & ~n1464 ) | ( n1447 & n2198 ) | ( ~n1464 & n2198 );
  assign n2202 = n1451 & n2201 ;
  assign n2203 = ( n1980 & n2200 ) | ( n1980 & n2202 ) | ( n2200 & n2202 );
  assign n2204 = n1981 & ~n2203 ;
  assign n2205 = n2197 | n2204 ;
  assign n2206 = n2197 & n2204 ;
  assign n2207 = n205 | n265 ;
  assign n2208 = n195 | n2207 ;
  assign n2209 = n156 | n2208 ;
  assign n2210 = n494 | n2209 ;
  assign n2211 = n235 | n2210 ;
  assign n2212 = n397 | n2211 ;
  assign n2213 = n346 | n2212 ;
  assign n2214 = n285 | n1026 ;
  assign n2215 = n357 | n2214 ;
  assign n2216 = n2024 | n2215 ;
  assign n2217 = n897 | n2216 ;
  assign n2218 = n142 | n293 ;
  assign n2219 = n2217 | n2218 ;
  assign n2220 = n127 | n2219 ;
  assign n2221 = n330 | n2220 ;
  assign n2222 = n148 | n877 ;
  assign n2223 = n394 | n2222 ;
  assign n2224 = n158 | n281 ;
  assign n2225 = n315 | n2224 ;
  assign n2226 = n430 | n2225 ;
  assign n2227 = n344 | n2226 ;
  assign n2228 = n2223 | n2227 ;
  assign n2229 = n2221 | n2228 ;
  assign n2230 = n2213 | n2229 ;
  assign n2231 = n305 | n2230 ;
  assign n2232 = n206 | n2231 ;
  assign n2233 = n262 | n2232 ;
  assign n2234 = n190 | n2233 ;
  assign n2235 = n389 | n2234 ;
  assign n2236 = n317 | n2235 ;
  assign n2237 = n312 | n2236 ;
  assign n2238 = n1338 & ~n1462 ;
  assign n2239 = ( n1447 & n1462 ) | ( n1447 & ~n2238 ) | ( n1462 & ~n2238 );
  assign n2240 = ( ~n1462 & n1470 ) | ( ~n1462 & n2238 ) | ( n1470 & n2238 );
  assign n2241 = ( n1980 & n2239 ) | ( n1980 & ~n2240 ) | ( n2239 & ~n2240 );
  assign n2242 = ~n1338 & n1462 ;
  assign n2243 = ~n1470 & n2242 ;
  assign n2244 = n1447 & n2242 ;
  assign n2245 = ( n1980 & n2243 ) | ( n1980 & n2244 ) | ( n2243 & n2244 );
  assign n2246 = n2241 & ~n2245 ;
  assign n2247 = n2237 & ~n2246 ;
  assign n2248 = n243 | n881 ;
  assign n2249 = n181 | n2248 ;
  assign n2250 = n937 | n939 ;
  assign n2251 = n205 | n315 ;
  assign n2252 = n148 | n331 ;
  assign n2253 = n123 | n2252 ;
  assign n2254 = n395 | n2253 ;
  assign n2255 = n2251 | n2254 ;
  assign n2256 = n1023 | n2255 ;
  assign n2257 = n422 | n2256 ;
  assign n2258 = n288 | n2257 ;
  assign n2259 = n2057 | n2258 ;
  assign n2260 = n2250 | n2259 ;
  assign n2261 = n2249 | n2260 ;
  assign n2262 = n158 | n548 ;
  assign n2263 = n2261 | n2262 ;
  assign n2264 = ( n1447 & ~n1470 ) | ( n1447 & n1980 ) | ( ~n1470 & n1980 );
  assign n2265 = n1339 & ~n1445 ;
  assign n2266 = n1339 & n1342 ;
  assign n2267 = ( n1980 & n2265 ) | ( n1980 & n2266 ) | ( n2265 & n2266 );
  assign n2268 = n2264 & ~n2267 ;
  assign n2269 = n2263 & ~n2268 ;
  assign n2270 = ~n2263 & n2268 ;
  assign n2271 = n214 | n316 ;
  assign n2272 = n383 | n2271 ;
  assign n2273 = n96 | n262 ;
  assign n2274 = n2272 | n2273 ;
  assign n2275 = n185 | n870 ;
  assign n2276 = n2274 | n2275 ;
  assign n2277 = n290 | n331 ;
  assign n2278 = n151 | n157 ;
  assign n2279 = n2277 | n2278 ;
  assign n2280 = n376 | n2279 ;
  assign n2281 = n2276 | n2280 ;
  assign n2282 = n268 | n285 ;
  assign n2283 = n189 | n287 ;
  assign n2284 = n2282 | n2283 ;
  assign n2285 = n245 | n322 ;
  assign n2286 = n153 | n2285 ;
  assign n2287 = n2284 | n2286 ;
  assign n2288 = n314 | n2035 ;
  assign n2289 = n683 | n2288 ;
  assign n2290 = n2287 | n2289 ;
  assign n2291 = n2281 | n2290 ;
  assign n2292 = n286 | n304 ;
  assign n2293 = n260 | n2292 ;
  assign n2294 = n277 | n2293 ;
  assign n2295 = n330 | n2294 ;
  assign n2296 = n2291 | n2295 ;
  assign n2297 = n170 | n2296 ;
  assign n2298 = ( n1342 & ~n1445 ) | ( n1342 & n1980 ) | ( ~n1445 & n1980 );
  assign n2299 = ( n1342 & n1980 ) | ( n1342 & ~n2298 ) | ( n1980 & ~n2298 );
  assign n2300 = ( n1445 & n2298 ) | ( n1445 & ~n2299 ) | ( n2298 & ~n2299 );
  assign n2301 = n2297 & ~n2300 ;
  assign n2302 = n152 | n216 ;
  assign n2303 = n389 | n2302 ;
  assign n2304 = n451 | n2303 ;
  assign n2305 = n322 | n2304 ;
  assign n2306 = n146 | n2305 ;
  assign n2307 = n474 | n2306 ;
  assign n2308 = n115 | n287 ;
  assign n2309 = n312 | n2308 ;
  assign n2310 = n498 | n2309 ;
  assign n2311 = n135 | n2310 ;
  assign n2312 = n209 | n2311 ;
  assign n2313 = n334 | n2312 ;
  assign n2314 = n2051 | n2313 ;
  assign n2315 = n311 | n2314 ;
  assign n2316 = n2307 | n2315 ;
  assign n2317 = n123 | n2316 ;
  assign n2318 = n927 | n2317 ;
  assign n2319 = n462 | n2318 ;
  assign n2320 = n281 | n2319 ;
  assign n2321 = n728 | n2320 ;
  assign n2322 = n190 | n272 ;
  assign n2323 = n198 | n2322 ;
  assign n2324 = n494 | n2323 ;
  assign n2325 = n101 | n2324 ;
  assign n2326 = n2321 | n2325 ;
  assign n2327 = n161 | n383 ;
  assign n2328 = n345 | n2327 ;
  assign n2329 = n2326 | n2328 ;
  assign n2330 = n1540 | n1978 ;
  assign n2331 = n1540 & n1978 ;
  assign n2332 = n2330 & ~n2331 ;
  assign n2333 = n2329 & ~n2332 ;
  assign n2334 = n112 | n414 ;
  assign n2335 = n294 | n669 ;
  assign n2336 = n2334 | n2335 ;
  assign n2337 = n2306 | n2336 ;
  assign n2338 = n898 & ~n2337 ;
  assign n2339 = ~n859 & n2338 ;
  assign n2340 = ~n932 & n2339 ;
  assign n2341 = n316 | n345 ;
  assign n2342 = n947 | n2341 ;
  assign n2343 = n247 | n549 ;
  assign n2344 = n124 | n2343 ;
  assign n2345 = n162 | n2344 ;
  assign n2346 = n2342 | n2345 ;
  assign n2347 = n2157 | n2346 ;
  assign n2348 = n385 | n2347 ;
  assign n2349 = n888 | n2348 ;
  assign n2350 = n459 | n2349 ;
  assign n2351 = n243 | n2350 ;
  assign n2352 = n170 | n552 ;
  assign n2353 = n311 | n2352 ;
  assign n2354 = n2351 | n2353 ;
  assign n2355 = n2340 & ~n2354 ;
  assign n2356 = ~n471 & n2355 ;
  assign n2357 = ~n305 & n2356 ;
  assign n2358 = ~n220 & n2357 ;
  assign n2359 = ~n200 & n2358 ;
  assign n2360 = ~n334 & n2359 ;
  assign n2361 = ~n123 & n2360 ;
  assign n2362 = ( ~n1544 & n1580 ) | ( ~n1544 & n1977 ) | ( n1580 & n1977 );
  assign n2363 = ( n1580 & n1977 ) | ( n1580 & ~n2362 ) | ( n1977 & ~n2362 );
  assign n2364 = ( n1544 & n2362 ) | ( n1544 & ~n2363 ) | ( n2362 & ~n2363 );
  assign n2365 = n2361 | n2364 ;
  assign n2366 = n2361 & n2364 ;
  assign n2367 = n361 | n2341 ;
  assign n2368 = n155 | n2367 ;
  assign n2369 = n2057 | n2368 ;
  assign n2370 = n265 | n330 ;
  assign n2371 = n383 | n2370 ;
  assign n2372 = n181 | n1027 ;
  assign n2373 = n2371 | n2372 ;
  assign n2374 = n225 | n268 ;
  assign n2375 = n333 | n2374 ;
  assign n2376 = n236 | n2375 ;
  assign n2377 = n358 | n2376 ;
  assign n2378 = n323 | n2377 ;
  assign n2379 = n2373 | n2378 ;
  assign n2380 = n142 | n459 ;
  assign n2381 = n436 | n2380 ;
  assign n2382 = n400 | n2381 ;
  assign n2383 = n2379 | n2382 ;
  assign n2384 = n2369 | n2383 ;
  assign n2385 = n656 | n2384 ;
  assign n2386 = n162 | n2385 ;
  assign n2387 = n282 | n293 ;
  assign n2388 = n2386 | n2387 ;
  assign n2389 = n177 | n278 ;
  assign n2390 = n195 | n2389 ;
  assign n2391 = n2388 | n2390 ;
  assign n2392 = n235 | n322 ;
  assign n2393 = n312 | n2392 ;
  assign n2394 = n2391 | n2393 ;
  assign n2395 = n1973 | n1975 ;
  assign n2396 = n1973 & n1975 ;
  assign n2397 = n2395 & ~n2396 ;
  assign n2398 = n2394 & ~n2397 ;
  assign n2399 = ~n2394 & n2397 ;
  assign n2400 = n702 | n1049 ;
  assign n2401 = n241 | n2400 ;
  assign n2402 = n385 | n2401 ;
  assign n2403 = n862 | n2402 ;
  assign n2404 = n2315 | n2403 ;
  assign n2405 = n722 | n2115 ;
  assign n2406 = n189 | n2405 ;
  assign n2407 = n2404 | n2406 ;
  assign n2408 = n278 | n552 ;
  assign n2409 = n120 | n2408 ;
  assign n2410 = n246 | n2409 ;
  assign n2411 = n2407 | n2410 ;
  assign n2412 = n1680 | n1971 ;
  assign n2413 = n1680 & ~n1971 ;
  assign n2414 = ( ~n1680 & n2412 ) | ( ~n1680 & n2413 ) | ( n2412 & n2413 );
  assign n2415 = ~n2411 & n2414 ;
  assign n2416 = n2398 | n2415 ;
  assign n2417 = n2399 | n2416 ;
  assign n2418 = ~n2398 & n2417 ;
  assign n2419 = n2365 & ~n2418 ;
  assign n2420 = ~n2366 & n2419 ;
  assign n2421 = n2365 & ~n2420 ;
  assign n2422 = ~n2329 & n2332 ;
  assign n2423 = n2333 | n2422 ;
  assign n2424 = n2421 | n2423 ;
  assign n2425 = ~n2333 & n2424 ;
  assign n2426 = ~n2297 & n2300 ;
  assign n2427 = n2301 | n2426 ;
  assign n2428 = n2425 | n2427 ;
  assign n2429 = ~n2301 & n2428 ;
  assign n2430 = n2269 | n2429 ;
  assign n2431 = n2270 | n2430 ;
  assign n2432 = ~n2269 & n2431 ;
  assign n2433 = n2237 & ~n2247 ;
  assign n2434 = n2246 | n2247 ;
  assign n2435 = ~n2433 & n2434 ;
  assign n2436 = n2432 | n2435 ;
  assign n2437 = ~n2247 & n2436 ;
  assign n2438 = n2205 & ~n2437 ;
  assign n2439 = ~n2206 & n2438 ;
  assign n2440 = n2205 & ~n2439 ;
  assign n2441 = n420 | n455 ;
  assign n2442 = n140 | n2441 ;
  assign n2443 = n265 | n2442 ;
  assign n2444 = n189 | n2443 ;
  assign n2445 = n195 | n2444 ;
  assign n2446 = n240 | n2445 ;
  assign n2447 = n163 | n2309 ;
  assign n2448 = n2178 | n2447 ;
  assign n2449 = n460 | n2448 ;
  assign n2450 = n450 | n2449 ;
  assign n2451 = n357 | n2450 ;
  assign n2452 = n2446 | n2451 ;
  assign n2453 = n2171 | n2452 ;
  assign n2454 = n259 | n2453 ;
  assign n2455 = n198 | n2454 ;
  assign n2456 = n383 | n2455 ;
  assign n2457 = ( n2155 & n2440 ) | ( n2155 & ~n2456 ) | ( n2440 & ~n2456 );
  assign n2458 = n2140 | n2440 ;
  assign n2459 = ~n2140 & n2456 ;
  assign n2460 = ( n2155 & n2458 ) | ( n2155 & ~n2459 ) | ( n2458 & ~n2459 );
  assign n2461 = ( ~n2143 & n2457 ) | ( ~n2143 & n2460 ) | ( n2457 & n2460 );
  assign n2462 = ( ~n2140 & n2143 ) | ( ~n2140 & n2461 ) | ( n2143 & n2461 );
  assign n2463 = ~n2076 & n2077 ;
  assign n2464 = n1982 & ~n2124 ;
  assign n2465 = n1984 | n2124 ;
  assign n2466 = ( n842 & n2464 ) | ( n842 & ~n2465 ) | ( n2464 & ~n2465 );
  assign n2467 = n797 | n2124 ;
  assign n2468 = n753 | n2124 ;
  assign n2469 = ( ~n638 & n2467 ) | ( ~n638 & n2468 ) | ( n2467 & n2468 );
  assign n2470 = ( n635 & n2466 ) | ( n635 & ~n2469 ) | ( n2466 & ~n2469 );
  assign n2471 = ( n2077 & ~n2124 ) | ( n2077 & n2470 ) | ( ~n2124 & n2470 );
  assign n2472 = ( ~n2077 & n2463 ) | ( ~n2077 & n2471 ) | ( n2463 & n2471 );
  assign n2473 = n2126 | n2472 ;
  assign n2474 = ~n2126 & n2473 ;
  assign n2475 = ( ~n2126 & n2462 ) | ( ~n2126 & n2474 ) | ( n2462 & n2474 );
  assign n2476 = n2075 & n2475 ;
  assign n2477 = ( ~n2050 & n2075 ) | ( ~n2050 & n2476 ) | ( n2075 & n2476 );
  assign n2478 = n689 | n693 ;
  assign n2479 = n282 | n556 ;
  assign n2480 = n289 | n2479 ;
  assign n2481 = n262 | n304 ;
  assign n2482 = n157 | n278 ;
  assign n2483 = n2481 | n2482 ;
  assign n2484 = n120 | n2483 ;
  assign n2485 = n328 | n658 ;
  assign n2486 = n394 | n2485 ;
  assign n2487 = n2080 | n2486 ;
  assign n2488 = n2484 | n2487 ;
  assign n2489 = n215 | n272 ;
  assign n2490 = n233 | n2489 ;
  assign n2491 = n2488 | n2490 ;
  assign n2492 = n333 | n2491 ;
  assign n2493 = n127 | n2492 ;
  assign n2494 = n549 | n2493 ;
  assign n2495 = n423 | n2494 ;
  assign n2496 = n552 | n2495 ;
  assign n2497 = n148 | n2496 ;
  assign n2498 = n161 | n2497 ;
  assign n2499 = n717 | n2272 ;
  assign n2500 = n153 | n2499 ;
  assign n2501 = n460 | n2500 ;
  assign n2502 = n2498 | n2501 ;
  assign n2503 = n2480 | n2502 ;
  assign n2504 = n180 | n2503 ;
  assign n2505 = n2478 | n2504 ;
  assign n2506 = n204 | n225 ;
  assign n2507 = n265 | n2506 ;
  assign n2508 = n184 | n2507 ;
  assign n2509 = n134 | n2508 ;
  assign n2510 = n236 | n2509 ;
  assign n2511 = n162 | n2510 ;
  assign n2512 = n2505 | n2511 ;
  assign n2513 = n2477 & ~n2512 ;
  assign n2514 = n254 & n2513 ;
  assign n2515 = n194 | n213 ;
  assign n2516 = n332 | n2515 ;
  assign n2517 = n291 | n1070 ;
  assign n2518 = n2516 | n2517 ;
  assign n2519 = n288 | n2518 ;
  assign n2520 = n274 | n2519 ;
  assign n2521 = n172 | n559 ;
  assign n2522 = n320 | n2521 ;
  assign n2523 = n177 | n196 ;
  assign n2524 = n2522 | n2523 ;
  assign n2525 = n284 | n2524 ;
  assign n2526 = n2520 | n2525 ;
  assign n2527 = n2514 & ~n2526 ;
  assign n2528 = n126 | n331 ;
  assign n2529 = n558 | n2528 ;
  assign n2530 = n555 | n2529 ;
  assign n2531 = n565 | n2530 ;
  assign n2532 = n172 | n212 ;
  assign n2533 = n301 | n2532 ;
  assign n2534 = n2531 | n2533 ;
  assign n2535 = n185 | n190 ;
  assign n2536 = n322 | n2535 ;
  assign n2537 = n2534 | n2536 ;
  assign n2538 = n2527 & ~n2537 ;
  assign n2539 = ~n2527 & n2537 ;
  assign n2540 = n2538 | n2539 ;
  assign n2541 = pi1 & ~n26 ;
  assign n2542 = ~pi1 & n26 ;
  assign n2543 = n2541 | n2542 ;
  assign n2544 = n32 & ~n2543 ;
  assign n2545 = ~n32 & n2543 ;
  assign n2546 = n2544 | n2545 ;
  assign n2547 = pi0 & ~n2546 ;
  assign n2548 = n2540 & n2547 ;
  assign n2549 = n254 | n2513 ;
  assign n2550 = ~n2514 & n2549 ;
  assign n2551 = ~n29 & n2546 ;
  assign n2552 = ~n2550 & n2551 ;
  assign n2553 = n2514 | n2526 ;
  assign n2554 = n2514 & n2526 ;
  assign n2555 = n2553 & ~n2554 ;
  assign n2556 = ~pi0 & n2543 ;
  assign n2557 = n2555 & n2556 ;
  assign n2558 = n2552 | n2557 ;
  assign n2559 = n2548 | n2558 ;
  assign n2560 = n2540 | n2555 ;
  assign n2561 = n2540 & n2555 ;
  assign n2562 = n2560 & ~n2561 ;
  assign n2563 = n2550 & ~n2555 ;
  assign n2564 = ( n2048 & ~n2073 ) | ( n2048 & n2475 ) | ( ~n2073 & n2475 );
  assign n2565 = ~n2048 & n2073 ;
  assign n2566 = ( n2050 & ~n2564 ) | ( n2050 & n2565 ) | ( ~n2564 & n2565 );
  assign n2567 = n2477 | n2566 ;
  assign n2568 = n2050 & ~n2475 ;
  assign n2569 = n2050 | n2475 ;
  assign n2570 = ( ~n2050 & n2568 ) | ( ~n2050 & n2569 ) | ( n2568 & n2569 );
  assign n2571 = n2567 & ~n2570 ;
  assign n2572 = n2462 | n2473 ;
  assign n2573 = n2462 & n2473 ;
  assign n2574 = n2572 & ~n2573 ;
  assign n2575 = ~n2570 & n2574 ;
  assign n2576 = n2570 & ~n2574 ;
  assign n2577 = n2575 | n2576 ;
  assign n2578 = ( ~n2140 & n2143 ) | ( ~n2140 & n2457 ) | ( n2143 & n2457 );
  assign n2579 = ( n2140 & ~n2143 ) | ( n2140 & n2578 ) | ( ~n2143 & n2578 );
  assign n2580 = ( ~n2457 & n2578 ) | ( ~n2457 & n2579 ) | ( n2578 & n2579 );
  assign n2581 = n2574 & n2580 ;
  assign n2582 = ( ~n2155 & n2440 ) | ( ~n2155 & n2456 ) | ( n2440 & n2456 );
  assign n2583 = ( n2440 & n2456 ) | ( n2440 & ~n2582 ) | ( n2456 & ~n2582 );
  assign n2584 = ( n2155 & n2582 ) | ( n2155 & ~n2583 ) | ( n2582 & ~n2583 );
  assign n2585 = n2580 & n2584 ;
  assign n2586 = n2574 | n2580 ;
  assign n2587 = ~n2581 & n2586 ;
  assign n2588 = ~n2206 & n2440 ;
  assign n2589 = n2437 | n2439 ;
  assign n2590 = ~n2588 & n2589 ;
  assign n2591 = ~n2432 & n2436 ;
  assign n2592 = ~n2435 & n2436 ;
  assign n2593 = n2591 | n2592 ;
  assign n2594 = ~n2590 & n2593 ;
  assign n2595 = ~n2429 & n2431 ;
  assign n2596 = ~n2270 & n2432 ;
  assign n2597 = n2595 | n2596 ;
  assign n2598 = n2593 & n2597 ;
  assign n2599 = n2593 | n2597 ;
  assign n2600 = ~n2598 & n2599 ;
  assign n2601 = n2425 & n2427 ;
  assign n2602 = n2428 & ~n2601 ;
  assign n2603 = n2597 & n2602 ;
  assign n2604 = n2421 & n2423 ;
  assign n2605 = n2424 & ~n2604 ;
  assign n2606 = n2602 & n2605 ;
  assign n2607 = n2418 | n2420 ;
  assign n2608 = ~n2366 & n2421 ;
  assign n2609 = n2607 & ~n2608 ;
  assign n2610 = n2605 & ~n2609 ;
  assign n2611 = ~n2605 & n2609 ;
  assign n2612 = ~n2415 & n2417 ;
  assign n2613 = ~n2399 & n2418 ;
  assign n2614 = n2612 | n2613 ;
  assign n2615 = n2411 & ~n2414 ;
  assign n2616 = n2415 | n2615 ;
  assign n2617 = n2609 & ~n2616 ;
  assign n2618 = n2614 & ~n2617 ;
  assign n2619 = ~n2611 & n2618 ;
  assign n2620 = ~n2610 & n2619 ;
  assign n2621 = n2610 | n2620 ;
  assign n2622 = n2602 | n2605 ;
  assign n2623 = n2621 & n2622 ;
  assign n2624 = ~n2606 & n2623 ;
  assign n2625 = n2606 | n2624 ;
  assign n2626 = n2597 | n2602 ;
  assign n2627 = ~n2603 & n2626 ;
  assign n2628 = n2625 & n2627 ;
  assign n2629 = n2603 | n2628 ;
  assign n2630 = n2598 | n2629 ;
  assign n2631 = ( n2598 & n2600 ) | ( n2598 & n2630 ) | ( n2600 & n2630 );
  assign n2632 = n2590 & ~n2593 ;
  assign n2633 = n2594 | n2632 ;
  assign n2634 = ~n2594 & n2633 ;
  assign n2635 = ( n2594 & n2631 ) | ( n2594 & ~n2634 ) | ( n2631 & ~n2634 );
  assign n2636 = n2580 | n2584 ;
  assign n2637 = ~n2585 & n2636 ;
  assign n2638 = n2584 & ~n2590 ;
  assign n2639 = ~n2584 & n2590 ;
  assign n2640 = n2638 | n2639 ;
  assign n2641 = ~n2638 & n2640 ;
  assign n2642 = n2637 & ~n2641 ;
  assign n2643 = n2637 & n2638 ;
  assign n2644 = ( n2635 & n2642 ) | ( n2635 & n2643 ) | ( n2642 & n2643 );
  assign n2645 = ( n2585 & n2587 ) | ( n2585 & n2644 ) | ( n2587 & n2644 );
  assign n2646 = n2581 | n2645 ;
  assign n2647 = n2575 | n2646 ;
  assign n2648 = ( n2575 & ~n2577 ) | ( n2575 & n2647 ) | ( ~n2577 & n2647 );
  assign n2649 = ~n2567 & n2570 ;
  assign n2650 = n2571 | n2649 ;
  assign n2651 = ~n2571 & n2650 ;
  assign n2652 = ( n2571 & n2648 ) | ( n2571 & ~n2651 ) | ( n2648 & ~n2651 );
  assign n2653 = n2477 | n2512 ;
  assign n2654 = n2477 & n2512 ;
  assign n2655 = n2653 & ~n2654 ;
  assign n2656 = ~n2550 & n2655 ;
  assign n2657 = n2550 & ~n2655 ;
  assign n2658 = n2656 | n2657 ;
  assign n2659 = n2567 & n2655 ;
  assign n2660 = n2567 | n2655 ;
  assign n2661 = ~n2659 & n2660 ;
  assign n2662 = n2659 | n2661 ;
  assign n2663 = ~n2658 & n2662 ;
  assign n2664 = ~n2658 & n2659 ;
  assign n2665 = ( n2652 & n2663 ) | ( n2652 & n2664 ) | ( n2663 & n2664 );
  assign n2666 = ( ~n2550 & n2555 ) | ( ~n2550 & n2656 ) | ( n2555 & n2656 );
  assign n2667 = ( ~n2563 & n2665 ) | ( ~n2563 & n2666 ) | ( n2665 & n2666 );
  assign n2668 = n2562 | n2667 ;
  assign n2669 = n2562 & n2666 ;
  assign n2670 = n2562 & ~n2563 ;
  assign n2671 = ( n2665 & n2669 ) | ( n2665 & n2670 ) | ( n2669 & n2670 );
  assign n2672 = n2668 & ~n2671 ;
  assign n2673 = pi0 & n2546 ;
  assign n2674 = n2672 & n2673 ;
  assign n2675 = n2559 | n2674 ;
  assign n2676 = n32 | n2675 ;
  assign n2677 = n32 & n2675 ;
  assign n2678 = n2676 & ~n2677 ;
  assign n2679 = ~n851 & n969 ;
  assign n2680 = n851 & ~n969 ;
  assign n2681 = n2679 | n2680 ;
  assign n2682 = n1123 & ~n1238 ;
  assign n2683 = ~n1123 & n1238 ;
  assign n2684 = n2682 | n2683 ;
  assign n2685 = ~n2681 & n2684 ;
  assign n2686 = n2580 & n2685 ;
  assign n2687 = ~n851 & n1123 ;
  assign n2688 = n851 & ~n1123 ;
  assign n2689 = n2687 | n2688 ;
  assign n2690 = ~n2684 & n2689 ;
  assign n2691 = n2584 & n2690 ;
  assign n2692 = n2684 | n2689 ;
  assign n2693 = n2681 & ~n2692 ;
  assign n2694 = ~n2590 & n2693 ;
  assign n2695 = n2691 | n2694 ;
  assign n2696 = n2686 | n2695 ;
  assign n2697 = n2681 & n2684 ;
  assign n2698 = ~n2637 & n2641 ;
  assign n2699 = n2637 | n2638 ;
  assign n2700 = ( n2635 & ~n2698 ) | ( n2635 & n2699 ) | ( ~n2698 & n2699 );
  assign n2701 = ~n2644 & n2700 ;
  assign n2702 = n2697 & n2701 ;
  assign n2703 = n2696 | n2702 ;
  assign n2704 = n969 | n2703 ;
  assign n2705 = n969 & n2703 ;
  assign n2706 = n2704 & ~n2705 ;
  assign n2707 = ~n742 & n969 ;
  assign n2708 = n742 & ~n969 ;
  assign n2709 = n2707 | n2708 ;
  assign n2710 = n2616 & n2709 ;
  assign n2711 = n761 & ~n2710 ;
  assign n2712 = ~n742 & n750 ;
  assign n2713 = n742 & ~n750 ;
  assign n2714 = n2712 | n2713 ;
  assign n2715 = ~n2709 & n2714 ;
  assign n2716 = n2616 & n2715 ;
  assign n2717 = n750 & ~n761 ;
  assign n2718 = ~n750 & n761 ;
  assign n2719 = n2717 | n2718 ;
  assign n2720 = n2709 & ~n2719 ;
  assign n2721 = n2614 & n2720 ;
  assign n2722 = n2716 | n2721 ;
  assign n2723 = ~n2614 & n2616 ;
  assign n2724 = n2614 & ~n2616 ;
  assign n2725 = n2723 | n2724 ;
  assign n2726 = n2709 & n2719 ;
  assign n2727 = n2725 & n2726 ;
  assign n2728 = n2722 | n2727 ;
  assign n2729 = n761 | n2728 ;
  assign n2730 = n761 & n2728 ;
  assign n2731 = n2729 & ~n2730 ;
  assign n2732 = n2711 & n2731 ;
  assign n2733 = n2711 | n2731 ;
  assign n2734 = ~n2732 & n2733 ;
  assign n2735 = ~n2609 & n2693 ;
  assign n2736 = n2605 & n2690 ;
  assign n2737 = n2602 & n2685 ;
  assign n2738 = n2736 | n2737 ;
  assign n2739 = n2735 | n2738 ;
  assign n2740 = n2621 & ~n2624 ;
  assign n2741 = n2622 & ~n2625 ;
  assign n2742 = n2740 | n2741 ;
  assign n2743 = n2697 & n2742 ;
  assign n2744 = n2739 | n2743 ;
  assign n2745 = n969 | n2744 ;
  assign n2746 = n969 & n2744 ;
  assign n2747 = n2745 & ~n2746 ;
  assign n2748 = n2614 & n2690 ;
  assign n2749 = n2616 & ~n2692 ;
  assign n2750 = n2681 & n2749 ;
  assign n2751 = n2748 | n2750 ;
  assign n2752 = ~n2609 & n2684 ;
  assign n2753 = ~n2681 & n2752 ;
  assign n2754 = n2751 | n2753 ;
  assign n2755 = n2609 & ~n2724 ;
  assign n2756 = ~n2609 & n2724 ;
  assign n2757 = n2755 | n2756 ;
  assign n2758 = ( n2697 & n2753 ) | ( n2697 & ~n2757 ) | ( n2753 & ~n2757 );
  assign n2759 = ~n2697 & n2757 ;
  assign n2760 = ( n2751 & n2758 ) | ( n2751 & ~n2759 ) | ( n2758 & ~n2759 );
  assign n2761 = n2754 | n2760 ;
  assign n2762 = n969 | n2761 ;
  assign n2763 = n969 & n2761 ;
  assign n2764 = n2762 & ~n2763 ;
  assign n2765 = n2616 & n2690 ;
  assign n2766 = n2614 & n2684 ;
  assign n2767 = ~n2681 & n2766 ;
  assign n2768 = n2765 | n2767 ;
  assign n2769 = n2684 & n2725 ;
  assign n2770 = n2681 & n2769 ;
  assign n2771 = n969 | n2770 ;
  assign n2772 = n2768 | n2771 ;
  assign n2773 = ~n969 & n2772 ;
  assign n2774 = n2616 & n2684 ;
  assign n2775 = n969 & ~n2774 ;
  assign n2776 = n2772 & n2775 ;
  assign n2777 = n2768 | n2770 ;
  assign n2778 = n2775 & ~n2777 ;
  assign n2779 = ( n2773 & n2776 ) | ( n2773 & n2778 ) | ( n2776 & n2778 );
  assign n2780 = n2710 & n2779 ;
  assign n2781 = n2764 & n2780 ;
  assign n2782 = n2710 & ~n2781 ;
  assign n2783 = n2618 & ~n2620 ;
  assign n2784 = n2611 | n2621 ;
  assign n2785 = ~n2783 & n2784 ;
  assign n2786 = n2697 & ~n2785 ;
  assign n2787 = ~n2609 & n2690 ;
  assign n2788 = n2605 & n2685 ;
  assign n2789 = n2614 & n2693 ;
  assign n2790 = n2788 | n2789 ;
  assign n2791 = n2787 | n2790 ;
  assign n2792 = n2786 | n2791 ;
  assign n2793 = n969 & ~n2792 ;
  assign n2794 = n969 & ~n2793 ;
  assign n2795 = ( n2792 & n2793 ) | ( n2792 & ~n2794 ) | ( n2793 & ~n2794 );
  assign n2796 = ~n2781 & n2795 ;
  assign n2797 = n2764 & n2779 ;
  assign n2798 = n2795 & n2797 ;
  assign n2799 = ( n2782 & n2796 ) | ( n2782 & n2798 ) | ( n2796 & n2798 );
  assign n2800 = n2781 | n2799 ;
  assign n2801 = ( n2734 & n2747 ) | ( n2734 & n2800 ) | ( n2747 & n2800 );
  assign n2802 = n2625 | n2627 ;
  assign n2803 = ~n2628 & n2802 ;
  assign n2804 = n2697 & n2803 ;
  assign n2805 = n2597 & n2685 ;
  assign n2806 = n2605 & n2693 ;
  assign n2807 = n2602 & n2690 ;
  assign n2808 = n2806 | n2807 ;
  assign n2809 = n2805 | n2808 ;
  assign n2810 = n2804 | n2809 ;
  assign n2811 = n969 & n2810 ;
  assign n2812 = n2810 & ~n2811 ;
  assign n2813 = n969 & ~n2811 ;
  assign n2814 = n2812 | n2813 ;
  assign n2815 = ~n2609 & n2715 ;
  assign n2816 = n2605 & n2720 ;
  assign n2817 = ~n2709 & n2719 ;
  assign n2818 = ~n2714 & n2817 ;
  assign n2819 = n2614 & n2818 ;
  assign n2820 = n2816 | n2819 ;
  assign n2821 = n2815 | n2820 ;
  assign n2822 = n2726 & ~n2785 ;
  assign n2823 = n2821 | n2822 ;
  assign n2824 = n761 & n2823 ;
  assign n2825 = n761 | n2823 ;
  assign n2826 = ~n2824 & n2825 ;
  assign n2827 = n587 & ~n761 ;
  assign n2828 = ~n587 & n761 ;
  assign n2829 = n2827 | n2828 ;
  assign n2830 = n2616 & n2829 ;
  assign n2831 = ~n2609 & n2720 ;
  assign n2832 = n2616 & n2818 ;
  assign n2833 = n2614 & n2715 ;
  assign n2834 = n2832 | n2833 ;
  assign n2835 = n2831 | n2834 ;
  assign n2836 = n2726 & ~n2757 ;
  assign n2837 = n2835 | n2836 ;
  assign n2838 = n761 | n2837 ;
  assign n2839 = n761 & n2837 ;
  assign n2840 = n2838 & ~n2839 ;
  assign n2841 = n2732 & n2840 ;
  assign n2842 = ( n2826 & n2830 ) | ( n2826 & n2841 ) | ( n2830 & n2841 );
  assign n2843 = n587 & ~n599 ;
  assign n2844 = ~n587 & n599 ;
  assign n2845 = n2843 | n2844 ;
  assign n2846 = ~n2829 & n2845 ;
  assign n2847 = n2616 & n2846 ;
  assign n2848 = ~n2008 & n2829 ;
  assign n2849 = n2614 & n2848 ;
  assign n2850 = n2847 | n2849 ;
  assign n2851 = n2008 & n2829 ;
  assign n2852 = n2725 & n2851 ;
  assign n2853 = n2850 | n2852 ;
  assign n2854 = n516 & ~n2853 ;
  assign n2855 = n516 & ~n2854 ;
  assign n2856 = ( n2853 & n2854 ) | ( n2853 & ~n2855 ) | ( n2854 & ~n2855 );
  assign n2857 = n516 & n2856 ;
  assign n2858 = ~n2830 & n2857 ;
  assign n2859 = n516 | n2856 ;
  assign n2860 = ( ~n2830 & n2856 ) | ( ~n2830 & n2859 ) | ( n2856 & n2859 );
  assign n2861 = ~n2858 & n2860 ;
  assign n2862 = ~n2609 & n2818 ;
  assign n2863 = n2605 & n2715 ;
  assign n2864 = n2602 & n2720 ;
  assign n2865 = n2863 | n2864 ;
  assign n2866 = n2862 | n2865 ;
  assign n2867 = n2726 & n2742 ;
  assign n2868 = n2866 | n2867 ;
  assign n2869 = n761 | n2868 ;
  assign n2870 = n761 & n2868 ;
  assign n2871 = n2869 & ~n2870 ;
  assign n2872 = ( n2842 & n2861 ) | ( n2842 & n2871 ) | ( n2861 & n2871 );
  assign n2873 = ( n2861 & n2871 ) | ( n2861 & ~n2872 ) | ( n2871 & ~n2872 );
  assign n2874 = ( n2842 & ~n2872 ) | ( n2842 & n2873 ) | ( ~n2872 & n2873 );
  assign n2875 = n2597 & n2693 ;
  assign n2876 = n2593 & n2690 ;
  assign n2877 = n2875 | n2876 ;
  assign n2878 = ~n2590 & n2685 ;
  assign n2879 = n2877 | n2878 ;
  assign n2880 = n2631 & ~n2633 ;
  assign n2881 = ~n2631 & n2633 ;
  assign n2882 = n2880 | n2881 ;
  assign n2883 = n2697 & ~n2882 ;
  assign n2884 = n2879 | n2883 ;
  assign n2885 = n969 & n2884 ;
  assign n2886 = n2884 & ~n2885 ;
  assign n2887 = n969 & ~n2885 ;
  assign n2888 = n2886 | n2887 ;
  assign n2889 = ( n2826 & n2830 ) | ( n2826 & ~n2842 ) | ( n2830 & ~n2842 );
  assign n2890 = ( n2841 & ~n2842 ) | ( n2841 & n2889 ) | ( ~n2842 & n2889 );
  assign n2891 = n2593 & n2685 ;
  assign n2892 = n2602 & n2693 ;
  assign n2893 = n2597 & n2690 ;
  assign n2894 = n2892 | n2893 ;
  assign n2895 = n2891 | n2894 ;
  assign n2896 = n2600 & n2629 ;
  assign n2897 = n2600 | n2629 ;
  assign n2898 = ~n2896 & n2897 ;
  assign n2899 = n2697 & n2898 ;
  assign n2900 = n2895 | n2899 ;
  assign n2901 = n969 | n2900 ;
  assign n2902 = n969 & n2900 ;
  assign n2903 = n2901 & ~n2902 ;
  assign n2904 = n2890 & n2903 ;
  assign n2905 = ( n2874 & n2888 ) | ( n2874 & n2904 ) | ( n2888 & n2904 );
  assign n2906 = n2890 & ~n2903 ;
  assign n2907 = ( n2903 & ~n2904 ) | ( n2903 & n2906 ) | ( ~n2904 & n2906 );
  assign n2908 = n2874 | n2888 ;
  assign n2909 = ( n2905 & n2907 ) | ( n2905 & n2908 ) | ( n2907 & n2908 );
  assign n2910 = ( n2814 & n2905 ) | ( n2814 & n2909 ) | ( n2905 & n2909 );
  assign n2911 = n2732 | n2840 ;
  assign n2912 = ~n2841 & n2911 ;
  assign n2913 = ( n2905 & n2909 ) | ( n2905 & n2912 ) | ( n2909 & n2912 );
  assign n2914 = ( n2801 & n2910 ) | ( n2801 & n2913 ) | ( n2910 & n2913 );
  assign n2915 = ~n2609 & n2846 ;
  assign n2916 = n2605 & n2848 ;
  assign n2917 = n2008 & ~n2829 ;
  assign n2918 = ~n2845 & n2917 ;
  assign n2919 = n2614 & n2918 ;
  assign n2920 = n2916 | n2919 ;
  assign n2921 = n2915 | n2920 ;
  assign n2922 = ~n2785 & n2851 ;
  assign n2923 = n2921 | n2922 ;
  assign n2924 = n516 & n2923 ;
  assign n2925 = n2923 & ~n2924 ;
  assign n2926 = n516 & ~n2924 ;
  assign n2927 = n2925 | n2926 ;
  assign n2928 = n516 & n2616 ;
  assign n2929 = ~n2609 & n2848 ;
  assign n2930 = n2616 & n2918 ;
  assign n2931 = n2614 & n2846 ;
  assign n2932 = n2930 | n2931 ;
  assign n2933 = n2929 | n2932 ;
  assign n2934 = ~n2757 & n2851 ;
  assign n2935 = n2933 | n2934 ;
  assign n2936 = n516 | n2935 ;
  assign n2937 = n516 & n2935 ;
  assign n2938 = n2936 & ~n2937 ;
  assign n2939 = n2858 & n2938 ;
  assign n2940 = ( n2927 & n2928 ) | ( n2927 & n2939 ) | ( n2928 & n2939 );
  assign n2941 = ( n2927 & n2928 ) | ( n2927 & ~n2940 ) | ( n2928 & ~n2940 );
  assign n2942 = n2726 & n2898 ;
  assign n2943 = n2593 & n2720 ;
  assign n2944 = n2602 & n2818 ;
  assign n2945 = n2597 & n2715 ;
  assign n2946 = n2944 | n2945 ;
  assign n2947 = n2943 | n2946 ;
  assign n2948 = n2942 | n2947 ;
  assign n2949 = n761 & n2948 ;
  assign n2950 = n761 | n2948 ;
  assign n2951 = ~n2949 & n2950 ;
  assign n2952 = ~n2940 & n2951 ;
  assign n2953 = n2938 & n2951 ;
  assign n2954 = n2858 & n2953 ;
  assign n2955 = ( n2941 & n2952 ) | ( n2941 & n2954 ) | ( n2952 & n2954 );
  assign n2956 = n2940 & ~n2951 ;
  assign n2957 = n2938 | n2951 ;
  assign n2958 = ( n2858 & n2951 ) | ( n2858 & n2957 ) | ( n2951 & n2957 );
  assign n2959 = ( n2941 & ~n2956 ) | ( n2941 & n2958 ) | ( ~n2956 & n2958 );
  assign n2960 = ~n2955 & n2959 ;
  assign n2961 = n2858 | n2938 ;
  assign n2962 = ~n2939 & n2961 ;
  assign n2963 = n2597 & n2720 ;
  assign n2964 = n2605 & n2818 ;
  assign n2965 = n2602 & n2715 ;
  assign n2966 = n2964 | n2965 ;
  assign n2967 = n2963 | n2966 ;
  assign n2968 = n2726 & n2803 ;
  assign n2969 = n2967 | n2968 ;
  assign n2970 = n761 | n2969 ;
  assign n2971 = n761 & n2969 ;
  assign n2972 = n2970 & ~n2971 ;
  assign n2973 = n2962 & n2972 ;
  assign n2974 = n2962 | n2972 ;
  assign n2975 = ~n2973 & n2974 ;
  assign n2976 = n2872 | n2973 ;
  assign n2977 = ( n2973 & n2975 ) | ( n2973 & n2976 ) | ( n2975 & n2976 );
  assign n2978 = n2960 | n2977 ;
  assign n2979 = n2960 & n2977 ;
  assign n2980 = n2978 & ~n2979 ;
  assign n2981 = n2584 & n2685 ;
  assign n2982 = ~n2590 & n2690 ;
  assign n2983 = n2593 & n2693 ;
  assign n2984 = n2982 | n2983 ;
  assign n2985 = n2981 | n2984 ;
  assign n2986 = n2635 & ~n2640 ;
  assign n2987 = ~n2635 & n2640 ;
  assign n2988 = n2986 | n2987 ;
  assign n2989 = n2697 & ~n2988 ;
  assign n2990 = n2985 | n2989 ;
  assign n2991 = n969 | n2990 ;
  assign n2992 = n969 & n2990 ;
  assign n2993 = n2991 & ~n2992 ;
  assign n2994 = n2872 | n2975 ;
  assign n2995 = n2872 & n2975 ;
  assign n2996 = n2994 & ~n2995 ;
  assign n2997 = n2993 & n2996 ;
  assign n2998 = n2993 & ~n2997 ;
  assign n2999 = ~n2993 & n2996 ;
  assign n3000 = n2997 | n2999 ;
  assign n3001 = n2998 | n3000 ;
  assign n3002 = ( n2706 & ~n2980 ) | ( n2706 & n3001 ) | ( ~n2980 & n3001 );
  assign n3003 = ( n2706 & ~n2980 ) | ( n2706 & n2997 ) | ( ~n2980 & n2997 );
  assign n3004 = ( n2914 & n3002 ) | ( n2914 & n3003 ) | ( n3002 & n3003 );
  assign n3005 = ( n2914 & n2997 ) | ( n2914 & n3001 ) | ( n2997 & n3001 );
  assign n3006 = ( n2706 & ~n3004 ) | ( n2706 & n3005 ) | ( ~n3004 & n3005 );
  assign n3007 = ~n1238 & n1291 ;
  assign n3008 = n1238 & ~n1291 ;
  assign n3009 = n3007 | n3008 ;
  assign n3010 = n32 & ~n1356 ;
  assign n3011 = ~n32 & n1356 ;
  assign n3012 = n3010 | n3011 ;
  assign n3013 = ~n3009 & n3012 ;
  assign n3014 = n2567 & n3013 ;
  assign n3015 = n1291 & ~n1356 ;
  assign n3016 = ~n1291 & n1356 ;
  assign n3017 = n3015 | n3016 ;
  assign n3018 = n3009 & ~n3012 ;
  assign n3019 = ~n3017 & n3018 ;
  assign n3020 = n2574 & n3019 ;
  assign n3021 = ~n3012 & n3017 ;
  assign n3022 = ~n2570 & n3021 ;
  assign n3023 = n3020 | n3022 ;
  assign n3024 = n3014 | n3023 ;
  assign n3025 = n2648 & ~n2650 ;
  assign n3026 = ~n2648 & n2650 ;
  assign n3027 = n3025 | n3026 ;
  assign n3028 = n3009 & n3012 ;
  assign n3029 = ~n3027 & n3028 ;
  assign n3030 = n3024 | n3029 ;
  assign n3031 = n1238 & n3030 ;
  assign n3032 = n1238 | n3030 ;
  assign n3033 = ~n3031 & n3032 ;
  assign n3034 = n3004 & n3033 ;
  assign n3035 = n2980 & n3033 ;
  assign n3036 = ( ~n3006 & n3034 ) | ( ~n3006 & n3035 ) | ( n3034 & n3035 );
  assign n3037 = n3004 | n3033 ;
  assign n3038 = n2980 | n3033 ;
  assign n3039 = ( ~n3006 & n3037 ) | ( ~n3006 & n3038 ) | ( n3037 & n3038 );
  assign n3040 = ~n3036 & n3039 ;
  assign n3041 = n2998 | n2999 ;
  assign n3042 = n2914 & n3041 ;
  assign n3043 = n2914 | n3041 ;
  assign n3044 = ~n3042 & n3043 ;
  assign n3045 = ~n2874 & n2888 ;
  assign n3046 = ( ~n2888 & n2908 ) | ( ~n2888 & n3045 ) | ( n2908 & n3045 );
  assign n3047 = ( n2890 & n2903 ) | ( n2890 & n2912 ) | ( n2903 & n2912 );
  assign n3048 = ~n2801 & n3046 ;
  assign n3049 = ( n2814 & n2890 ) | ( n2814 & n2903 ) | ( n2890 & n2903 );
  assign n3050 = n3046 & ~n3049 ;
  assign n3051 = ( ~n3047 & n3048 ) | ( ~n3047 & n3050 ) | ( n3048 & n3050 );
  assign n3052 = n3046 & ~n3051 ;
  assign n3053 = n2574 & n3013 ;
  assign n3054 = n2584 & n3019 ;
  assign n3055 = n2580 & n3021 ;
  assign n3056 = n3054 | n3055 ;
  assign n3057 = n3053 | n3056 ;
  assign n3058 = n2585 | n2587 ;
  assign n3059 = n2644 | n3058 ;
  assign n3060 = ~n2645 & n3059 ;
  assign n3061 = n3028 & n3060 ;
  assign n3062 = n3057 | n3061 ;
  assign n3063 = n1238 | n3062 ;
  assign n3064 = n1238 & n3062 ;
  assign n3065 = n3063 & ~n3064 ;
  assign n3066 = n3051 & n3065 ;
  assign n3067 = ( n2801 & n3047 ) | ( n2801 & n3049 ) | ( n3047 & n3049 );
  assign n3068 = n3065 & n3067 ;
  assign n3069 = ( ~n3052 & n3066 ) | ( ~n3052 & n3068 ) | ( n3066 & n3068 );
  assign n3070 = n3051 | n3065 ;
  assign n3071 = n3065 | n3067 ;
  assign n3072 = ( ~n3052 & n3070 ) | ( ~n3052 & n3071 ) | ( n3070 & n3071 );
  assign n3073 = ~n3069 & n3072 ;
  assign n3074 = ( n2801 & n2814 ) | ( n2801 & n2912 ) | ( n2814 & n2912 );
  assign n3075 = n2907 & ~n3074 ;
  assign n3076 = n2907 & n3074 ;
  assign n3077 = ( n3074 & n3075 ) | ( n3074 & ~n3076 ) | ( n3075 & ~n3076 );
  assign n3078 = n2580 & n3013 ;
  assign n3079 = n2584 & n3021 ;
  assign n3080 = ~n2590 & n3019 ;
  assign n3081 = n3079 | n3080 ;
  assign n3082 = n3078 | n3081 ;
  assign n3083 = n2701 & n3028 ;
  assign n3084 = n3082 | n3083 ;
  assign n3085 = n1238 | n3084 ;
  assign n3086 = n1238 & n3084 ;
  assign n3087 = n3085 & ~n3086 ;
  assign n3088 = ~n2988 & n3028 ;
  assign n3089 = ( n2814 & n2912 ) | ( n2814 & ~n3074 ) | ( n2912 & ~n3074 );
  assign n3090 = ( n2801 & ~n3074 ) | ( n2801 & n3089 ) | ( ~n3074 & n3089 );
  assign n3091 = n2584 & n3013 ;
  assign n3092 = ~n2590 & n3021 ;
  assign n3093 = n2593 & ~n3017 ;
  assign n3094 = n3018 & n3093 ;
  assign n3095 = n3092 | n3094 ;
  assign n3096 = n3091 | n3095 ;
  assign n3097 = ( n1238 & n3090 ) | ( n1238 & n3096 ) | ( n3090 & n3096 );
  assign n3098 = n1238 | n3090 ;
  assign n3099 = ( n3088 & n3097 ) | ( n3088 & n3098 ) | ( n3097 & n3098 );
  assign n3100 = n3088 | n3096 ;
  assign n3101 = ( n3090 & ~n3099 ) | ( n3090 & n3100 ) | ( ~n3099 & n3100 );
  assign n3102 = ( n1238 & ~n3099 ) | ( n1238 & n3101 ) | ( ~n3099 & n3101 );
  assign n3103 = ( ~n2734 & n2747 ) | ( ~n2734 & n2800 ) | ( n2747 & n2800 );
  assign n3104 = ( n2734 & ~n2800 ) | ( n2734 & n3103 ) | ( ~n2800 & n3103 );
  assign n3105 = ( ~n2747 & n3103 ) | ( ~n2747 & n3104 ) | ( n3103 & n3104 );
  assign n3106 = ~n2590 & n3013 ;
  assign n3107 = n2593 & n3021 ;
  assign n3108 = n2597 & ~n3017 ;
  assign n3109 = n3018 & n3108 ;
  assign n3110 = n3107 | n3109 ;
  assign n3111 = n3106 | n3110 ;
  assign n3112 = ~n2882 & n3028 ;
  assign n3113 = n3111 | n3112 ;
  assign n3114 = n1238 & n3113 ;
  assign n3115 = n1238 | n3113 ;
  assign n3116 = ~n3114 & n3115 ;
  assign n3117 = n3105 & n3116 ;
  assign n3118 = n3102 & n3117 ;
  assign n3119 = n2597 & n3013 ;
  assign n3120 = n2605 & n3019 ;
  assign n3121 = n2602 & n3021 ;
  assign n3122 = n3120 | n3121 ;
  assign n3123 = n3119 | n3122 ;
  assign n3124 = n2803 & n3028 ;
  assign n3125 = n3123 | n3124 ;
  assign n3126 = n1238 & n3125 ;
  assign n3127 = n1238 | n3125 ;
  assign n3128 = ~n3126 & n3127 ;
  assign n3129 = n2764 | n2779 ;
  assign n3130 = ~n2797 & n3129 ;
  assign n3131 = n3128 & n3130 ;
  assign n3132 = n3128 | n3130 ;
  assign n3133 = ~n3131 & n3132 ;
  assign n3134 = n2772 | n2775 ;
  assign n3135 = ~n2775 & n2777 ;
  assign n3136 = ( n2773 & n3134 ) | ( n2773 & ~n3135 ) | ( n3134 & ~n3135 );
  assign n3137 = ~n2779 & n3136 ;
  assign n3138 = ~n2609 & n3019 ;
  assign n3139 = n2605 & n3021 ;
  assign n3140 = n2602 & n3013 ;
  assign n3141 = n3139 | n3140 ;
  assign n3142 = n3138 | n3141 ;
  assign n3143 = n2742 & n3028 ;
  assign n3144 = n3142 | n3143 ;
  assign n3145 = n1238 | n3144 ;
  assign n3146 = n1238 & n3144 ;
  assign n3147 = n3145 & ~n3146 ;
  assign n3148 = n3137 & n3147 ;
  assign n3149 = n3137 | n3147 ;
  assign n3150 = ~n3148 & n3149 ;
  assign n3151 = n2614 & n3021 ;
  assign n3152 = n2616 & ~n3017 ;
  assign n3153 = n3018 & n3152 ;
  assign n3154 = n3151 | n3153 ;
  assign n3155 = ~n2609 & n3013 ;
  assign n3156 = n3154 | n3155 ;
  assign n3157 = ( ~n2757 & n3028 ) | ( ~n2757 & n3155 ) | ( n3028 & n3155 );
  assign n3158 = n2757 & ~n3028 ;
  assign n3159 = ( n3154 & n3157 ) | ( n3154 & ~n3158 ) | ( n3157 & ~n3158 );
  assign n3160 = n3156 | n3159 ;
  assign n3161 = n1238 | n3160 ;
  assign n3162 = n1238 & n3160 ;
  assign n3163 = n3161 & ~n3162 ;
  assign n3164 = ~n2609 & n3021 ;
  assign n3165 = n2605 & n3013 ;
  assign n3166 = n2614 & n3019 ;
  assign n3167 = n3165 | n3166 ;
  assign n3168 = n3164 | n3167 ;
  assign n3169 = ~n2785 & n3028 ;
  assign n3170 = n3168 | n3169 ;
  assign n3171 = n1238 & n3170 ;
  assign n3172 = n1238 | n3170 ;
  assign n3173 = ~n3171 & n3172 ;
  assign n3174 = n2616 & n3021 ;
  assign n3175 = n2614 & n3013 ;
  assign n3176 = n3174 | n3175 ;
  assign n3177 = n2725 & n3028 ;
  assign n3178 = n1238 & ~n3177 ;
  assign n3179 = ~n3176 & n3178 ;
  assign n3180 = n1238 & ~n3179 ;
  assign n3181 = n1238 & ~n2616 ;
  assign n3182 = ( n1238 & ~n3012 ) | ( n1238 & n3181 ) | ( ~n3012 & n3181 );
  assign n3183 = n3179 & n3182 ;
  assign n3184 = n3176 | n3177 ;
  assign n3185 = n3182 & n3184 ;
  assign n3186 = ( ~n3180 & n3183 ) | ( ~n3180 & n3185 ) | ( n3183 & n3185 );
  assign n3187 = ( n2774 & n3173 ) | ( n2774 & n3186 ) | ( n3173 & n3186 );
  assign n3188 = n2774 & n3173 ;
  assign n3189 = ( n3163 & n3187 ) | ( n3163 & n3188 ) | ( n3187 & n3188 );
  assign n3190 = n3150 & n3189 ;
  assign n3191 = n3131 | n3190 ;
  assign n3192 = n3131 | n3148 ;
  assign n3193 = ( n3133 & n3191 ) | ( n3133 & n3192 ) | ( n3191 & n3192 );
  assign n3194 = n3105 | n3116 ;
  assign n3195 = ~n3117 & n3194 ;
  assign n3196 = n2781 & ~n2795 ;
  assign n3197 = n2795 | n2797 ;
  assign n3198 = ( n2782 & ~n3196 ) | ( n2782 & n3197 ) | ( ~n3196 & n3197 );
  assign n3199 = ~n2799 & n3198 ;
  assign n3200 = n3195 & n3199 ;
  assign n3201 = n2593 & n3013 ;
  assign n3202 = n2602 & n3019 ;
  assign n3203 = n2597 & n3021 ;
  assign n3204 = n3202 | n3203 ;
  assign n3205 = n3201 | n3204 ;
  assign n3206 = ( n2898 & n3028 ) | ( n2898 & n3205 ) | ( n3028 & n3205 );
  assign n3207 = ( n1238 & ~n3028 ) | ( n1238 & n3205 ) | ( ~n3028 & n3205 );
  assign n3208 = ( n1238 & ~n2898 ) | ( n1238 & n3207 ) | ( ~n2898 & n3207 );
  assign n3209 = n3206 | n3208 ;
  assign n3210 = ~n3205 & n3208 ;
  assign n3211 = ( ~n1238 & n3209 ) | ( ~n1238 & n3210 ) | ( n3209 & n3210 );
  assign n3212 = n3195 & n3211 ;
  assign n3213 = ( n3193 & n3200 ) | ( n3193 & n3212 ) | ( n3200 & n3212 );
  assign n3214 = ( n3102 & n3118 ) | ( n3102 & n3213 ) | ( n3118 & n3213 );
  assign n3215 = n1238 & n3100 ;
  assign n3216 = n3099 & ~n3215 ;
  assign n3217 = n3214 | n3216 ;
  assign n3218 = ( n3077 & n3087 ) | ( n3077 & n3217 ) | ( n3087 & n3217 );
  assign n3219 = n3069 | n3218 ;
  assign n3220 = ( n3069 & n3073 ) | ( n3069 & n3219 ) | ( n3073 & n3219 );
  assign n3221 = ~n2570 & n3013 ;
  assign n3222 = n2580 & n3019 ;
  assign n3223 = n2574 & n3021 ;
  assign n3224 = n3222 | n3223 ;
  assign n3225 = n3221 | n3224 ;
  assign n3226 = ~n2577 & n2646 ;
  assign n3227 = n2577 & ~n2646 ;
  assign n3228 = n3226 | n3227 ;
  assign n3229 = n3028 & ~n3228 ;
  assign n3230 = n3225 | n3229 ;
  assign n3231 = n1238 & n3230 ;
  assign n3232 = n1238 | n3230 ;
  assign n3233 = ~n3231 & n3232 ;
  assign n3234 = ( n3044 & n3220 ) | ( n3044 & n3233 ) | ( n3220 & n3233 );
  assign n3235 = n3040 & n3234 ;
  assign n3236 = n3040 | n3234 ;
  assign n3237 = ~n3235 & n3236 ;
  assign n3238 = n2547 & n2555 ;
  assign n3239 = n2551 & n2655 ;
  assign n3240 = ~n2550 & n2556 ;
  assign n3241 = n3239 | n3240 ;
  assign n3242 = n3238 | n3241 ;
  assign n3243 = ~n2550 & n2555 ;
  assign n3244 = ( n2550 & ~n2555 ) | ( n2550 & n2656 ) | ( ~n2555 & n2656 );
  assign n3245 = ( n2665 & ~n3243 ) | ( n2665 & n3244 ) | ( ~n3243 & n3244 );
  assign n3246 = n2656 | n2665 ;
  assign n3247 = ( n2550 & ~n3245 ) | ( n2550 & n3246 ) | ( ~n3245 & n3246 );
  assign n3248 = ( n2555 & n3245 ) | ( n2555 & ~n3247 ) | ( n3245 & ~n3247 );
  assign n3249 = n2673 & ~n3248 ;
  assign n3250 = n3242 | n3249 ;
  assign n3251 = n32 | n3250 ;
  assign n3252 = n32 & n3250 ;
  assign n3253 = n3251 & ~n3252 ;
  assign n3254 = n3237 & n3253 ;
  assign n3255 = ~n3237 & n3253 ;
  assign n3256 = ( n3237 & ~n3254 ) | ( n3237 & n3255 ) | ( ~n3254 & n3255 );
  assign n3257 = n2547 & ~n2550 ;
  assign n3258 = n2551 & n2567 ;
  assign n3259 = n2556 & n2655 ;
  assign n3260 = n3258 | n3259 ;
  assign n3261 = n3257 | n3260 ;
  assign n3262 = ( n2652 & n2659 ) | ( n2652 & n2662 ) | ( n2659 & n2662 );
  assign n3263 = n2658 & ~n3262 ;
  assign n3264 = n2665 | n3263 ;
  assign n3265 = n2673 & ~n3264 ;
  assign n3266 = n3261 | n3265 ;
  assign n3267 = n32 | n3266 ;
  assign n3268 = n32 & n3266 ;
  assign n3269 = n3267 & ~n3268 ;
  assign n3270 = ( n3044 & ~n3220 ) | ( n3044 & n3233 ) | ( ~n3220 & n3233 );
  assign n3271 = ( n3220 & ~n3234 ) | ( n3220 & n3270 ) | ( ~n3234 & n3270 );
  assign n3272 = ( ~n3077 & n3087 ) | ( ~n3077 & n3217 ) | ( n3087 & n3217 );
  assign n3273 = ( n3077 & ~n3218 ) | ( n3077 & n3272 ) | ( ~n3218 & n3272 );
  assign n3274 = ~n29 & n2580 ;
  assign n3275 = n2546 & n3274 ;
  assign n3276 = pi0 & ~n3228 ;
  assign n3277 = n2556 & n2574 ;
  assign n3278 = ( n2546 & n3276 ) | ( n2546 & n3277 ) | ( n3276 & n3277 );
  assign n3279 = n2546 | n3276 ;
  assign n3280 = ( n3275 & n3278 ) | ( n3275 & n3279 ) | ( n3278 & n3279 );
  assign n3281 = pi0 & ~n2570 ;
  assign n3282 = ( ~n2546 & n3277 ) | ( ~n2546 & n3281 ) | ( n3277 & n3281 );
  assign n3283 = n2546 & ~n3281 ;
  assign n3284 = ( n3275 & n3282 ) | ( n3275 & ~n3283 ) | ( n3282 & ~n3283 );
  assign n3285 = n3280 | n3284 ;
  assign n3286 = ~n32 & n3285 ;
  assign n3287 = n32 & ~n3285 ;
  assign n3288 = n3286 | n3287 ;
  assign n3289 = n3102 | n3117 ;
  assign n3290 = n3213 | n3289 ;
  assign n3291 = ~n3214 & n3290 ;
  assign n3292 = n3195 | n3199 ;
  assign n3293 = n3195 | n3211 ;
  assign n3294 = ( n3193 & n3292 ) | ( n3193 & n3293 ) | ( n3292 & n3293 );
  assign n3295 = ~n3213 & n3294 ;
  assign n3296 = ( n3288 & n3291 ) | ( n3288 & n3295 ) | ( n3291 & n3295 );
  assign n3297 = pi0 & n2544 ;
  assign n3298 = n3060 & n3297 ;
  assign n3299 = n2556 & n2580 ;
  assign n3300 = pi0 & n2574 ;
  assign n3301 = ( ~n2546 & n3299 ) | ( ~n2546 & n3300 ) | ( n3299 & n3300 );
  assign n3302 = ~n29 & n2584 ;
  assign n3303 = ( n2546 & n3299 ) | ( n2546 & n3302 ) | ( n3299 & n3302 );
  assign n3304 = n3301 | n3303 ;
  assign n3305 = n32 | n3304 ;
  assign n3306 = n2673 | n3305 ;
  assign n3307 = ( n3060 & n3305 ) | ( n3060 & n3306 ) | ( n3305 & n3306 );
  assign n3308 = ~n3298 & n3307 ;
  assign n3309 = n32 & n3304 ;
  assign n3310 = n3308 & ~n3309 ;
  assign n3311 = ( n3288 & n3291 ) | ( n3288 & n3310 ) | ( n3291 & n3310 );
  assign n3312 = n2556 & n2593 ;
  assign n3313 = pi0 & ~n2590 ;
  assign n3314 = ( ~n2546 & n3312 ) | ( ~n2546 & n3313 ) | ( n3312 & n3313 );
  assign n3315 = ~n29 & n2597 ;
  assign n3316 = ( n2546 & n3312 ) | ( n2546 & n3315 ) | ( n3312 & n3315 );
  assign n3317 = n3314 | n3316 ;
  assign n3318 = n2673 | n3317 ;
  assign n3319 = ( ~n2882 & n3317 ) | ( ~n2882 & n3318 ) | ( n3317 & n3318 );
  assign n3320 = n32 | n3319 ;
  assign n3321 = ~n32 & n3319 ;
  assign n3322 = ( ~n3319 & n3320 ) | ( ~n3319 & n3321 ) | ( n3320 & n3321 );
  assign n3323 = n2673 & n2898 ;
  assign n3324 = n2556 & n2597 ;
  assign n3325 = pi0 & n2593 ;
  assign n3326 = ( ~n2546 & n3324 ) | ( ~n2546 & n3325 ) | ( n3324 & n3325 );
  assign n3327 = ~n29 & n2602 ;
  assign n3328 = ( n2546 & n3324 ) | ( n2546 & n3327 ) | ( n3324 & n3327 );
  assign n3329 = n3326 | n3328 ;
  assign n3330 = n3323 | n3329 ;
  assign n3331 = n3163 & n3186 ;
  assign n3332 = n3163 | n3186 ;
  assign n3333 = ~n3331 & n3332 ;
  assign n3334 = n2898 & n3297 ;
  assign n3335 = n3179 | n3182 ;
  assign n3336 = n3182 | n3184 ;
  assign n3337 = ( ~n3180 & n3335 ) | ( ~n3180 & n3336 ) | ( n3335 & n3336 );
  assign n3338 = ~n3186 & n3337 ;
  assign n3339 = n2616 & n3012 ;
  assign n3340 = pi0 & ~n2785 ;
  assign n3341 = n2546 & n3340 ;
  assign n3342 = pi0 & n2605 ;
  assign n3343 = n2556 & ~n2609 ;
  assign n3344 = ( ~n2546 & n3342 ) | ( ~n2546 & n3343 ) | ( n3342 & n3343 );
  assign n3345 = n2546 & ~n3342 ;
  assign n3346 = ( n3341 & n3344 ) | ( n3341 & ~n3345 ) | ( n3344 & ~n3345 );
  assign n3347 = ~n29 & n2614 ;
  assign n3348 = ( n2546 & n3343 ) | ( n2546 & n3347 ) | ( n3343 & n3347 );
  assign n3349 = n2546 | n3347 ;
  assign n3350 = ( n3341 & n3348 ) | ( n3341 & n3349 ) | ( n3348 & n3349 );
  assign n3351 = n3346 | n3350 ;
  assign n3352 = n32 & n3351 ;
  assign n3353 = n32 | n3351 ;
  assign n3354 = ~n3352 & n3353 ;
  assign n3355 = pi0 & n2614 ;
  assign n3356 = ~n2546 & n3355 ;
  assign n3357 = n32 & ~n2616 ;
  assign n3358 = ( n32 & ~n2556 ) | ( n32 & n3357 ) | ( ~n2556 & n3357 );
  assign n3359 = ~n3356 & n3358 ;
  assign n3360 = n2547 & ~n2609 ;
  assign n3361 = n2551 & n2616 ;
  assign n3362 = n2556 & n2614 ;
  assign n3363 = n3361 | n3362 ;
  assign n3364 = n3360 | n3363 ;
  assign n3365 = n32 & n3364 ;
  assign n3366 = pi0 & n2725 ;
  assign n3367 = n2544 & n3366 ;
  assign n3368 = n3365 | n3367 ;
  assign n3369 = n2616 | n2757 ;
  assign n3370 = n2544 & ~n3369 ;
  assign n3371 = ( pi0 & n2616 ) | ( pi0 & n3370 ) | ( n2616 & n3370 );
  assign n3372 = n3368 | n3371 ;
  assign n3373 = n3359 & ~n3372 ;
  assign n3374 = ( n3339 & n3354 ) | ( n3339 & n3373 ) | ( n3354 & n3373 );
  assign n3375 = n29 | n2609 ;
  assign n3376 = n2546 & ~n3375 ;
  assign n3377 = n2556 & n2605 ;
  assign n3378 = pi0 & n2602 ;
  assign n3379 = ~n2546 & n3378 ;
  assign n3380 = n3377 | n3379 ;
  assign n3381 = ( ~n32 & n3376 ) | ( ~n32 & n3380 ) | ( n3376 & n3380 );
  assign n3382 = n32 & ~n3375 ;
  assign n3383 = n2546 & n3382 ;
  assign n3384 = pi0 & n2742 ;
  assign n3385 = n2546 & n3384 ;
  assign n3386 = ( n32 & ~n3383 ) | ( n32 & n3385 ) | ( ~n3383 & n3385 );
  assign n3387 = ~n3380 & n3386 ;
  assign n3388 = ( n3381 & ~n3383 ) | ( n3381 & n3387 ) | ( ~n3383 & n3387 );
  assign n3389 = n2544 & n3384 ;
  assign n3390 = n3388 & ~n3389 ;
  assign n3391 = ( n3338 & n3374 ) | ( n3338 & n3390 ) | ( n3374 & n3390 );
  assign n3392 = ~n3334 & n3391 ;
  assign n3393 = n2547 & n2597 ;
  assign n3394 = n2551 & n2605 ;
  assign n3395 = n2556 & n2602 ;
  assign n3396 = n3394 | n3395 ;
  assign n3397 = n3393 | n3396 ;
  assign n3398 = n2673 & n2803 ;
  assign n3399 = n3397 | n3398 ;
  assign n3400 = n32 & ~n3399 ;
  assign n3401 = ( ~n32 & n3399 ) | ( ~n32 & n3400 ) | ( n3399 & n3400 );
  assign n3402 = n3400 | n3401 ;
  assign n3403 = ~n3334 & n3402 ;
  assign n3404 = ( n3333 & n3392 ) | ( n3333 & n3403 ) | ( n3392 & n3403 );
  assign n3405 = ( n32 & n3330 ) | ( n32 & n3404 ) | ( n3330 & n3404 );
  assign n3406 = ( n32 & n3330 ) | ( n32 & ~n3334 ) | ( n3330 & ~n3334 );
  assign n3407 = ( ~n2774 & n3173 ) | ( ~n2774 & n3186 ) | ( n3173 & n3186 );
  assign n3408 = ~n2774 & n3173 ;
  assign n3409 = ( n3163 & n3407 ) | ( n3163 & n3408 ) | ( n3407 & n3408 );
  assign n3410 = ( n2774 & ~n3331 ) | ( n2774 & n3409 ) | ( ~n3331 & n3409 );
  assign n3411 = ( ~n3173 & n3409 ) | ( ~n3173 & n3410 ) | ( n3409 & n3410 );
  assign n3412 = ( n3405 & n3406 ) | ( n3405 & n3411 ) | ( n3406 & n3411 );
  assign n3413 = ( n32 & n3329 ) | ( n32 & ~n3404 ) | ( n3329 & ~n3404 );
  assign n3414 = ( n32 & n3329 ) | ( n32 & n3334 ) | ( n3329 & n3334 );
  assign n3415 = ( ~n3411 & n3413 ) | ( ~n3411 & n3414 ) | ( n3413 & n3414 );
  assign n3416 = n3412 & ~n3415 ;
  assign n3417 = n3322 & n3391 ;
  assign n3418 = n3322 & n3402 ;
  assign n3419 = ( n3333 & n3417 ) | ( n3333 & n3418 ) | ( n3417 & n3418 );
  assign n3420 = n3411 & n3419 ;
  assign n3421 = ( n3322 & n3416 ) | ( n3322 & n3420 ) | ( n3416 & n3420 );
  assign n3422 = n3150 | n3189 ;
  assign n3423 = ~n3190 & n3422 ;
  assign n3424 = n3322 | n3391 ;
  assign n3425 = n3322 | n3402 ;
  assign n3426 = ( n3333 & n3424 ) | ( n3333 & n3425 ) | ( n3424 & n3425 );
  assign n3427 = ( n3322 & n3411 ) | ( n3322 & n3426 ) | ( n3411 & n3426 );
  assign n3428 = n3423 & n3427 ;
  assign n3429 = ( n3416 & n3423 ) | ( n3416 & n3428 ) | ( n3423 & n3428 );
  assign n3430 = n3421 | n3429 ;
  assign n3431 = ( n3193 & n3199 ) | ( n3193 & n3211 ) | ( n3199 & n3211 );
  assign n3432 = ( n3193 & n3199 ) | ( n3193 & ~n3431 ) | ( n3199 & ~n3431 );
  assign n3433 = n2701 & n3297 ;
  assign n3434 = n2556 & n2584 ;
  assign n3435 = n29 | n2590 ;
  assign n3436 = ( n2546 & n3434 ) | ( n2546 & ~n3435 ) | ( n3434 & ~n3435 );
  assign n3437 = pi0 & n2580 ;
  assign n3438 = ( ~n2546 & n3434 ) | ( ~n2546 & n3437 ) | ( n3434 & n3437 );
  assign n3439 = n3436 | n3438 ;
  assign n3440 = n2673 | n3439 ;
  assign n3441 = ( n2701 & n3439 ) | ( n2701 & n3440 ) | ( n3439 & n3440 );
  assign n3442 = ( n32 & ~n3433 ) | ( n32 & n3441 ) | ( ~n3433 & n3441 );
  assign n3443 = ( n32 & n3297 ) | ( n32 & n3439 ) | ( n3297 & n3439 );
  assign n3444 = n32 & n3439 ;
  assign n3445 = ( n2701 & n3443 ) | ( n2701 & n3444 ) | ( n3443 & n3444 );
  assign n3446 = n3442 & ~n3445 ;
  assign n3447 = ( n3133 & n3148 ) | ( n3133 & n3190 ) | ( n3148 & n3190 );
  assign n3448 = n3148 | n3190 ;
  assign n3449 = n3133 | n3448 ;
  assign n3450 = ~n3447 & n3449 ;
  assign n3451 = ( ~n3431 & n3446 ) | ( ~n3431 & n3450 ) | ( n3446 & n3450 );
  assign n3452 = ( n3211 & n3446 ) | ( n3211 & n3450 ) | ( n3446 & n3450 );
  assign n3453 = ( n3432 & n3451 ) | ( n3432 & n3452 ) | ( n3451 & n3452 );
  assign n3454 = ~n2988 & n3297 ;
  assign n3455 = n2556 & ~n2590 ;
  assign n3456 = pi0 & n2584 ;
  assign n3457 = ( ~n2546 & n3455 ) | ( ~n2546 & n3456 ) | ( n3455 & n3456 );
  assign n3458 = ~n29 & n2593 ;
  assign n3459 = ( n2546 & n3455 ) | ( n2546 & n3458 ) | ( n3455 & n3458 );
  assign n3460 = n3457 | n3459 ;
  assign n3461 = n2673 | n3460 ;
  assign n3462 = ( ~n2988 & n3460 ) | ( ~n2988 & n3461 ) | ( n3460 & n3461 );
  assign n3463 = ( n32 & ~n3454 ) | ( n32 & n3462 ) | ( ~n3454 & n3462 );
  assign n3464 = ( n32 & n3297 ) | ( n32 & n3460 ) | ( n3297 & n3460 );
  assign n3465 = n32 & n3460 ;
  assign n3466 = ( ~n2988 & n3464 ) | ( ~n2988 & n3465 ) | ( n3464 & n3465 );
  assign n3467 = n3463 & ~n3466 ;
  assign n3468 = ( ~n3431 & n3446 ) | ( ~n3431 & n3467 ) | ( n3446 & n3467 );
  assign n3469 = ( n3211 & n3446 ) | ( n3211 & n3467 ) | ( n3446 & n3467 );
  assign n3470 = ( n3432 & n3468 ) | ( n3432 & n3469 ) | ( n3468 & n3469 );
  assign n3471 = ( n3430 & n3453 ) | ( n3430 & n3470 ) | ( n3453 & n3470 );
  assign n3472 = ( n3296 & n3311 ) | ( n3296 & n3471 ) | ( n3311 & n3471 );
  assign n3473 = n2673 & ~n3027 ;
  assign n3474 = n2547 & n2567 ;
  assign n3475 = n2551 & n2574 ;
  assign n3476 = n2556 & ~n2570 ;
  assign n3477 = n3475 | n3476 ;
  assign n3478 = n3474 | n3477 ;
  assign n3479 = n3473 | n3478 ;
  assign n3480 = n32 | n3479 ;
  assign n3481 = n32 & n3479 ;
  assign n3482 = n3480 & ~n3481 ;
  assign n3483 = ( n3273 & n3472 ) | ( n3273 & n3482 ) | ( n3472 & n3482 );
  assign n3484 = n3073 & n3218 ;
  assign n3485 = n3073 | n3218 ;
  assign n3486 = ~n3484 & n3485 ;
  assign n3487 = n2547 & n2655 ;
  assign n3488 = n2551 & ~n2570 ;
  assign n3489 = n2556 & n2567 ;
  assign n3490 = n3488 | n3489 ;
  assign n3491 = n3487 | n3490 ;
  assign n3492 = n2652 & n2661 ;
  assign n3493 = n2652 | n2661 ;
  assign n3494 = ~n3492 & n3493 ;
  assign n3495 = n2673 & n3494 ;
  assign n3496 = n3491 | n3495 ;
  assign n3497 = n32 & ~n3496 ;
  assign n3498 = ( ~n32 & n3496 ) | ( ~n32 & n3497 ) | ( n3496 & n3497 );
  assign n3499 = n3497 | n3498 ;
  assign n3500 = ( n3483 & n3486 ) | ( n3483 & n3499 ) | ( n3486 & n3499 );
  assign n3501 = ( n3269 & n3271 ) | ( n3269 & n3500 ) | ( n3271 & n3500 );
  assign n3502 = n3256 & n3501 ;
  assign n3503 = n3254 | n3502 ;
  assign n3504 = ~n2609 & n2918 ;
  assign n3505 = n2605 & n2846 ;
  assign n3506 = n2602 & n2848 ;
  assign n3507 = n3505 | n3506 ;
  assign n3508 = n3504 | n3507 ;
  assign n3509 = n2742 & n2851 ;
  assign n3510 = n3508 | n3509 ;
  assign n3511 = n516 & n3510 ;
  assign n3512 = n516 & n2614 ;
  assign n3513 = ~n3511 & n3512 ;
  assign n3514 = n3512 & ~n3513 ;
  assign n3515 = ( n516 & n3510 ) | ( n516 & ~n3513 ) | ( n3510 & ~n3513 );
  assign n3516 = ( ~n3511 & n3514 ) | ( ~n3511 & n3515 ) | ( n3514 & n3515 );
  assign n3517 = n2726 & ~n2882 ;
  assign n3518 = ~n2590 & n2720 ;
  assign n3519 = n2597 & n2818 ;
  assign n3520 = n2593 & n2715 ;
  assign n3521 = n3519 | n3520 ;
  assign n3522 = n3518 | n3521 ;
  assign n3523 = n3517 | n3522 ;
  assign n3524 = n761 & n3523 ;
  assign n3525 = n761 | n3523 ;
  assign n3526 = ~n3524 & n3525 ;
  assign n3527 = ( n2940 & n3516 ) | ( n2940 & ~n3526 ) | ( n3516 & ~n3526 );
  assign n3528 = ( ~n2940 & n3526 ) | ( ~n2940 & n3527 ) | ( n3526 & n3527 );
  assign n3529 = ( ~n3516 & n3527 ) | ( ~n3516 & n3528 ) | ( n3527 & n3528 );
  assign n3530 = n2955 | n2979 ;
  assign n3531 = ~n3529 & n3530 ;
  assign n3532 = n3529 & ~n3530 ;
  assign n3533 = n3531 | n3532 ;
  assign n3534 = n2574 & n2685 ;
  assign n3535 = n2584 & n2693 ;
  assign n3536 = n2580 & n2690 ;
  assign n3537 = n3535 | n3536 ;
  assign n3538 = n3534 | n3537 ;
  assign n3539 = n2697 & n3060 ;
  assign n3540 = n3538 | n3539 ;
  assign n3541 = n969 | n3540 ;
  assign n3542 = n969 & n3540 ;
  assign n3543 = n3541 & ~n3542 ;
  assign n3544 = n3533 & n3543 ;
  assign n3545 = n3533 | n3543 ;
  assign n3546 = ~n3544 & n3545 ;
  assign n3547 = n2706 | n2980 ;
  assign n3548 = n3546 & n3547 ;
  assign n3549 = n2706 & n2980 ;
  assign n3550 = n3546 & n3549 ;
  assign n3551 = ( n2706 & n2980 ) | ( n2706 & ~n2997 ) | ( n2980 & ~n2997 );
  assign n3552 = n3547 & ~n3551 ;
  assign n3553 = ( n3546 & n3550 ) | ( n3546 & n3552 ) | ( n3550 & n3552 );
  assign n3554 = ( n3041 & n3548 ) | ( n3041 & n3553 ) | ( n3548 & n3553 );
  assign n3555 = n3548 & n3553 ;
  assign n3556 = ( n2914 & n3554 ) | ( n2914 & n3555 ) | ( n3554 & n3555 );
  assign n3557 = n3546 | n3547 ;
  assign n3558 = n3546 | n3549 ;
  assign n3559 = n3552 | n3558 ;
  assign n3560 = ( n3041 & n3557 ) | ( n3041 & n3559 ) | ( n3557 & n3559 );
  assign n3561 = n3557 & n3559 ;
  assign n3562 = ( n2914 & n3560 ) | ( n2914 & n3561 ) | ( n3560 & n3561 );
  assign n3563 = ~n3556 & n3562 ;
  assign n3564 = n2655 & n3013 ;
  assign n3565 = ~n2570 & n3019 ;
  assign n3566 = n2567 & n3021 ;
  assign n3567 = n3565 | n3566 ;
  assign n3568 = n3564 | n3567 ;
  assign n3569 = n3028 & n3494 ;
  assign n3570 = n3568 | n3569 ;
  assign n3571 = n1238 & n3570 ;
  assign n3572 = n1238 | n3570 ;
  assign n3573 = ~n3571 & n3572 ;
  assign n3574 = n3563 & n3573 ;
  assign n3575 = n3563 | n3573 ;
  assign n3576 = ~n3574 & n3575 ;
  assign n3577 = n3036 | n3235 ;
  assign n3578 = n3576 | n3577 ;
  assign n3579 = ( n3036 & n3040 ) | ( n3036 & n3576 ) | ( n3040 & n3576 );
  assign n3580 = n3036 & n3576 ;
  assign n3581 = ( n3234 & n3579 ) | ( n3234 & n3580 ) | ( n3579 & n3580 );
  assign n3582 = n3578 & ~n3581 ;
  assign n3583 = ( n2678 & n3503 ) | ( n2678 & n3582 ) | ( n3503 & n3582 );
  assign n3584 = ( ~n2678 & n3503 ) | ( ~n2678 & n3582 ) | ( n3503 & n3582 );
  assign n3585 = ( n2678 & ~n3583 ) | ( n2678 & n3584 ) | ( ~n3583 & n3584 );
  assign n3586 = n186 | n2484 ;
  assign n3587 = n487 | n3586 ;
  assign n3588 = n277 | n3587 ;
  assign n3589 = n131 | n3588 ;
  assign n3590 = n96 | n123 ;
  assign n3591 = n2162 | n3590 ;
  assign n3592 = n265 | n281 ;
  assign n3593 = n191 | n272 ;
  assign n3594 = n3592 | n3593 ;
  assign n3595 = n311 | n322 ;
  assign n3596 = n3594 | n3595 ;
  assign n3597 = n3591 | n3596 ;
  assign n3598 = n222 | n3597 ;
  assign n3599 = n286 | n3598 ;
  assign n3600 = n204 | n3599 ;
  assign n3601 = n190 | n213 ;
  assign n3602 = n3600 | n3601 ;
  assign n3603 = n158 | n397 ;
  assign n3604 = n384 | n3603 ;
  assign n3605 = n3602 | n3604 ;
  assign n3606 = n220 | n3605 ;
  assign n3607 = n233 | n3606 ;
  assign n3608 = n106 | n3607 ;
  assign n3609 = n430 | n3608 ;
  assign n3610 = n361 | n2022 ;
  assign n3611 = n3609 | n3610 ;
  assign n3612 = n2480 | n3611 ;
  assign n3613 = n3589 | n3612 ;
  assign n3614 = n471 | n3613 ;
  assign n3615 = n224 | n3614 ;
  assign n3616 = n183 | n3615 ;
  assign n3617 = n195 | n3616 ;
  assign n3618 = n451 | n3617 ;
  assign n3619 = n423 | n3618 ;
  assign n3620 = n124 | n3619 ;
  assign n3621 = n148 | n3620 ;
  assign n3622 = n234 | n423 ;
  assign n3623 = n240 | n3622 ;
  assign n3624 = n345 | n3623 ;
  assign n3625 = n400 | n3624 ;
  assign n3626 = n669 | n3625 ;
  assign n3627 = n283 | n3626 ;
  assign n3628 = n180 | n3627 ;
  assign n3629 = n184 | n3628 ;
  assign n3630 = n287 | n3629 ;
  assign n3631 = n271 | n459 ;
  assign n3632 = n3630 | n3631 ;
  assign n3633 = n148 | n321 ;
  assign n3634 = n3632 | n3633 ;
  assign n3635 = n398 | n1098 ;
  assign n3636 = n260 | n3635 ;
  assign n3637 = n2026 | n3636 ;
  assign n3638 = n158 | n214 ;
  assign n3639 = n245 | n548 ;
  assign n3640 = n3638 | n3639 ;
  assign n3641 = n3637 | n3640 ;
  assign n3642 = n169 | n312 ;
  assign n3643 = n384 | n3642 ;
  assign n3644 = n657 | n3643 ;
  assign n3645 = n189 | n3644 ;
  assign n3646 = n3641 | n3645 ;
  assign n3647 = n389 | n3646 ;
  assign n3648 = n2373 | n3647 ;
  assign n3649 = n3634 | n3648 ;
  assign n3650 = n199 | n2191 ;
  assign n3651 = n129 | n3650 ;
  assign n3652 = n290 | n3651 ;
  assign n3653 = n3649 | n3652 ;
  assign n3654 = n134 | n315 ;
  assign n3655 = n109 | n3654 ;
  assign n3656 = n549 | n3655 ;
  assign n3657 = n347 | n3656 ;
  assign n3658 = n161 | n3657 ;
  assign n3659 = n3653 | n3658 ;
  assign n3660 = n3256 | n3501 ;
  assign n3661 = ~n3502 & n3660 ;
  assign n3662 = n3269 & n3271 ;
  assign n3663 = n3269 & ~n3271 ;
  assign n3664 = ( n3271 & ~n3662 ) | ( n3271 & n3663 ) | ( ~n3662 & n3663 );
  assign n3665 = ~n3500 & n3664 ;
  assign n3666 = n291 | n2157 ;
  assign n3667 = n221 | n2213 ;
  assign n3668 = n3666 | n3667 ;
  assign n3669 = n162 | n1362 ;
  assign n3670 = n3668 | n3669 ;
  assign n3671 = n335 | n2341 ;
  assign n3672 = n2334 | n3671 ;
  assign n3673 = n422 | n3672 ;
  assign n3674 = n663 | n2021 ;
  assign n3675 = n199 | n3674 ;
  assign n3676 = n263 | n3675 ;
  assign n3677 = n3673 | n3676 ;
  assign n3678 = n3670 | n3677 ;
  assign n3679 = n2287 | n3678 ;
  assign n3680 = n215 | n3679 ;
  assign n3681 = n180 | n3680 ;
  assign n3682 = n259 | n3681 ;
  assign n3683 = n190 | n3682 ;
  assign n3684 = n292 | n3683 ;
  assign n3685 = n213 | n3684 ;
  assign n3686 = n115 | n3685 ;
  assign n3687 = ( ~n3664 & n3665 ) | ( ~n3664 & n3686 ) | ( n3665 & n3686 );
  assign n3688 = ( n3500 & n3665 ) | ( n3500 & n3687 ) | ( n3665 & n3687 );
  assign n3689 = ( n3659 & n3661 ) | ( n3659 & n3688 ) | ( n3661 & n3688 );
  assign n3690 = ( n3585 & ~n3621 ) | ( n3585 & n3689 ) | ( ~n3621 & n3689 );
  assign n3691 = ( n3585 & n3621 ) | ( n3585 & ~n3689 ) | ( n3621 & ~n3689 );
  assign n3692 = ( ~n3585 & n3690 ) | ( ~n3585 & n3691 ) | ( n3690 & n3691 );
  assign n3693 = n1046 | n3590 ;
  assign n3694 = n669 | n3693 ;
  assign n3695 = n1366 | n3694 ;
  assign n3696 = n2221 | n3695 ;
  assign n3697 = n382 | n3696 ;
  assign n3698 = n413 | n3697 ;
  assign n3699 = n2480 | n3698 ;
  assign n3700 = n214 | n3699 ;
  assign n3701 = n126 | n3700 ;
  assign n3702 = n241 | n3701 ;
  assign n3703 = n279 | n474 ;
  assign n3704 = n3590 | n3703 ;
  assign n3705 = n195 | n287 ;
  assign n3706 = n289 | n3705 ;
  assign n3707 = n3704 | n3706 ;
  assign n3708 = n312 | n344 ;
  assign n3709 = n3707 | n3708 ;
  assign n3710 = n343 | n442 ;
  assign n3711 = n2017 | n3710 ;
  assign n3712 = n3709 | n3711 ;
  assign n3713 = n247 | n3712 ;
  assign n3714 = n1094 & ~n3713 ;
  assign n3715 = n222 | n259 ;
  assign n3716 = n150 | n3715 ;
  assign n3717 = n213 | n3716 ;
  assign n3718 = n383 | n3717 ;
  assign n3719 = n3714 & ~n3718 ;
  assign n3720 = n358 | n430 ;
  assign n3721 = n311 | n3720 ;
  assign n3722 = n3719 & ~n3721 ;
  assign n3723 = n2538 & n3722 ;
  assign n3724 = n3722 & ~n3723 ;
  assign n3725 = ( n2538 & ~n3723 ) | ( n2538 & n3724 ) | ( ~n3723 & n3724 );
  assign n3726 = n2547 & ~n3725 ;
  assign n3727 = n2551 & n2555 ;
  assign n3728 = n2540 & n2556 ;
  assign n3729 = n3727 | n3728 ;
  assign n3730 = n3726 | n3729 ;
  assign n3731 = ~n2540 & n3725 ;
  assign n3732 = n2540 & ~n3725 ;
  assign n3733 = n3731 | n3732 ;
  assign n3734 = n2561 | n2669 ;
  assign n3735 = n3733 | n3734 ;
  assign n3736 = n2561 | n2670 ;
  assign n3737 = n3733 | n3736 ;
  assign n3738 = ( n2665 & n3735 ) | ( n2665 & n3737 ) | ( n3735 & n3737 );
  assign n3739 = ~n3733 & n3738 ;
  assign n3740 = ( n2665 & n3734 ) | ( n2665 & n3736 ) | ( n3734 & n3736 );
  assign n3741 = ( n3738 & n3739 ) | ( n3738 & ~n3740 ) | ( n3739 & ~n3740 );
  assign n3742 = n2673 & ~n3741 ;
  assign n3743 = n3730 | n3742 ;
  assign n3744 = n32 & n3743 ;
  assign n3745 = n3743 & ~n3744 ;
  assign n3746 = n32 & ~n3744 ;
  assign n3747 = n3745 | n3746 ;
  assign n3748 = ~n2570 & n2685 ;
  assign n3749 = n2574 & n2690 ;
  assign n3750 = n2580 & n2693 ;
  assign n3751 = n3749 | n3750 ;
  assign n3752 = n3748 | n3751 ;
  assign n3753 = n2697 & ~n3228 ;
  assign n3754 = n3752 | n3753 ;
  assign n3755 = n969 & n3754 ;
  assign n3756 = n3754 & ~n3755 ;
  assign n3757 = n969 & ~n3755 ;
  assign n3758 = n3756 | n3757 ;
  assign n3759 = n2940 | n3516 ;
  assign n3760 = n2955 & n3529 ;
  assign n3761 = ( n2979 & n3529 ) | ( n2979 & n3760 ) | ( n3529 & n3760 );
  assign n3762 = ( ~n3527 & n3759 ) | ( ~n3527 & n3761 ) | ( n3759 & n3761 );
  assign n3763 = n2584 & n2720 ;
  assign n3764 = n2593 & n2818 ;
  assign n3765 = ~n2590 & n2715 ;
  assign n3766 = n3764 | n3765 ;
  assign n3767 = n3763 | n3766 ;
  assign n3768 = n2726 & ~n2988 ;
  assign n3769 = n3767 | n3768 ;
  assign n3770 = n761 | n3769 ;
  assign n3771 = n761 & n3769 ;
  assign n3772 = n3770 & ~n3771 ;
  assign n3773 = n3513 | n3516 ;
  assign n3774 = n516 & n2609 ;
  assign n3775 = n2597 & n2848 ;
  assign n3776 = n2605 & n2918 ;
  assign n3777 = n2602 & n2846 ;
  assign n3778 = n3776 | n3777 ;
  assign n3779 = n3775 | n3778 ;
  assign n3780 = n2803 & n2851 ;
  assign n3781 = n3779 | n3780 ;
  assign n3782 = n3774 & n3781 ;
  assign n3783 = n3774 | n3781 ;
  assign n3784 = ~n3782 & n3783 ;
  assign n3785 = n2940 & n3784 ;
  assign n3786 = n3513 & n3784 ;
  assign n3787 = ( n3773 & n3785 ) | ( n3773 & n3786 ) | ( n3785 & n3786 );
  assign n3788 = n2940 | n3784 ;
  assign n3789 = n3513 | n3784 ;
  assign n3790 = ( n3773 & n3788 ) | ( n3773 & n3789 ) | ( n3788 & n3789 );
  assign n3791 = ~n3787 & n3790 ;
  assign n3792 = ( n3759 & n3772 ) | ( n3759 & n3791 ) | ( n3772 & n3791 );
  assign n3793 = ( ~n3527 & n3772 ) | ( ~n3527 & n3791 ) | ( n3772 & n3791 );
  assign n3794 = ( n3761 & n3792 ) | ( n3761 & n3793 ) | ( n3792 & n3793 );
  assign n3795 = ( n3772 & n3791 ) | ( n3772 & ~n3794 ) | ( n3791 & ~n3794 );
  assign n3796 = ( n3762 & ~n3794 ) | ( n3762 & n3795 ) | ( ~n3794 & n3795 );
  assign n3797 = n3758 & n3796 ;
  assign n3798 = n3758 & ~n3797 ;
  assign n3799 = ~n3758 & n3796 ;
  assign n3800 = n3798 | n3799 ;
  assign n3801 = n3544 | n3550 ;
  assign n3802 = n3544 | n3546 ;
  assign n3803 = ( n3552 & n3801 ) | ( n3552 & n3802 ) | ( n3801 & n3802 );
  assign n3804 = n3800 & n3803 ;
  assign n3805 = ( n3544 & n3547 ) | ( n3544 & n3802 ) | ( n3547 & n3802 );
  assign n3806 = n3799 & n3805 ;
  assign n3807 = ( n3798 & n3805 ) | ( n3798 & n3806 ) | ( n3805 & n3806 );
  assign n3808 = ( n3042 & n3804 ) | ( n3042 & n3807 ) | ( n3804 & n3807 );
  assign n3809 = ( n3041 & n3803 ) | ( n3041 & n3805 ) | ( n3803 & n3805 );
  assign n3810 = n3803 & n3805 ;
  assign n3811 = ( n2914 & n3809 ) | ( n2914 & n3810 ) | ( n3809 & n3810 );
  assign n3812 = n3800 | n3811 ;
  assign n3813 = ~n3808 & n3812 ;
  assign n3814 = n3574 | n3581 ;
  assign n3815 = ~n2550 & n3013 ;
  assign n3816 = n2567 & n3019 ;
  assign n3817 = n2655 & n3021 ;
  assign n3818 = n3816 | n3817 ;
  assign n3819 = n3815 | n3818 ;
  assign n3820 = n3028 & ~n3264 ;
  assign n3821 = n3819 | n3820 ;
  assign n3822 = n1238 | n3821 ;
  assign n3823 = n1238 & n3821 ;
  assign n3824 = n3822 & ~n3823 ;
  assign n3825 = ( ~n3813 & n3814 ) | ( ~n3813 & n3824 ) | ( n3814 & n3824 );
  assign n3826 = ( n3814 & n3824 ) | ( n3814 & ~n3825 ) | ( n3824 & ~n3825 );
  assign n3827 = ( n3813 & n3825 ) | ( n3813 & ~n3826 ) | ( n3825 & ~n3826 );
  assign n3828 = n3747 & n3827 ;
  assign n3829 = n3747 & ~n3828 ;
  assign n3830 = ~n3747 & n3827 ;
  assign n3831 = n3583 & n3830 ;
  assign n3832 = ( n3583 & n3829 ) | ( n3583 & n3831 ) | ( n3829 & n3831 );
  assign n3833 = n3583 | n3830 ;
  assign n3834 = n3829 | n3833 ;
  assign n3835 = ~n3832 & n3834 ;
  assign n3836 = n3702 | n3835 ;
  assign n3837 = n3702 & n3835 ;
  assign n3838 = n3836 & ~n3837 ;
  assign n3839 = ( n3585 & n3621 ) | ( n3585 & n3689 ) | ( n3621 & n3689 );
  assign n3840 = n3838 & n3839 ;
  assign n3841 = n3838 | n3839 ;
  assign n3842 = ~n3840 & n3841 ;
  assign n3843 = n3692 & n3842 ;
  assign n3844 = n3842 & ~n3843 ;
  assign n3845 = ( n3692 & ~n3843 ) | ( n3692 & n3844 ) | ( ~n3843 & n3844 );
  assign n3846 = pi22 & ~pi23 ;
  assign n3847 = ~pi22 & pi23 ;
  assign n3848 = n3846 | n3847 ;
  assign n3849 = n3845 & n3848 ;
  assign n3850 = n375 | n2251 ;
  assign n3851 = n2187 | n3850 ;
  assign n3852 = n683 | n3851 ;
  assign n3853 = n196 | n284 ;
  assign n3854 = n236 | n3853 ;
  assign n3855 = n101 | n3854 ;
  assign n3856 = n3852 | n3855 ;
  assign n3857 = n2480 | n3856 ;
  assign n3858 = n3605 | n3857 ;
  assign n3859 = n267 | n2486 ;
  assign n3860 = n3858 | n3859 ;
  assign n3861 = n263 | n3860 ;
  assign n3862 = n290 | n3861 ;
  assign n3863 = n157 | n3862 ;
  assign n3864 = n451 | n3863 ;
  assign n3865 = n312 | n3864 ;
  assign n3866 = n121 | n548 ;
  assign n3867 = n2162 | n2334 ;
  assign n3868 = n327 | n3867 ;
  assign n3869 = n683 | n3868 ;
  assign n3870 = n418 | n3869 ;
  assign n3871 = n451 | n3870 ;
  assign n3872 = n131 | n3871 ;
  assign n3873 = n488 | n853 ;
  assign n3874 = n665 | n3873 ;
  assign n3875 = n1364 & ~n1376 ;
  assign n3876 = ~n3874 & n3875 ;
  assign n3877 = ~n346 & n3876 ;
  assign n3878 = ( n2354 & ~n3872 ) | ( n2354 & n3877 ) | ( ~n3872 & n3877 );
  assign n3879 = ~n2354 & n3878 ;
  assign n3880 = ~n3866 & n3879 ;
  assign n3881 = ~n347 & n3880 ;
  assign n3882 = ~n146 & n3881 ;
  assign n3883 = ~n394 & n3882 ;
  assign n3884 = ~n3723 & n3883 ;
  assign n3885 = n3723 & ~n3883 ;
  assign n3886 = n3884 | n3885 ;
  assign n3887 = n3725 | n3886 ;
  assign n3888 = n3725 & n3886 ;
  assign n3889 = n3887 & ~n3888 ;
  assign n3890 = ~n3732 & n3733 ;
  assign n3891 = ( n2540 & n2561 ) | ( n2540 & ~n3725 ) | ( n2561 & ~n3725 );
  assign n3892 = ( n2670 & ~n3890 ) | ( n2670 & n3891 ) | ( ~n3890 & n3891 );
  assign n3893 = ( n2669 & ~n3890 ) | ( n2669 & n3891 ) | ( ~n3890 & n3891 );
  assign n3894 = ( n2665 & n3892 ) | ( n2665 & n3893 ) | ( n3892 & n3893 );
  assign n3895 = n3889 | n3894 ;
  assign n3896 = n3889 & n3894 ;
  assign n3897 = n3895 & ~n3896 ;
  assign n3898 = n2673 & n3897 ;
  assign n3899 = n2547 & ~n3886 ;
  assign n3900 = n2540 & n2551 ;
  assign n3901 = n2556 & ~n3725 ;
  assign n3902 = n3900 | n3901 ;
  assign n3903 = n3899 | n3902 ;
  assign n3904 = n3898 | n3903 ;
  assign n3905 = n32 & n3904 ;
  assign n3906 = n3904 & ~n3905 ;
  assign n3907 = n32 & ~n3905 ;
  assign n3908 = n3906 | n3907 ;
  assign n3909 = n2697 & ~n3027 ;
  assign n3910 = n2567 & n2685 ;
  assign n3911 = n2574 & n2693 ;
  assign n3912 = ~n2570 & n2690 ;
  assign n3913 = n3911 | n3912 ;
  assign n3914 = n3910 | n3913 ;
  assign n3915 = n3909 | n3914 ;
  assign n3916 = n969 & n3915 ;
  assign n3917 = n3915 & ~n3916 ;
  assign n3918 = n969 & ~n3916 ;
  assign n3919 = n3917 | n3918 ;
  assign n3920 = n2580 & n2720 ;
  assign n3921 = ~n2590 & n2818 ;
  assign n3922 = n2584 & n2715 ;
  assign n3923 = n3921 | n3922 ;
  assign n3924 = n3920 | n3923 ;
  assign n3925 = n2701 & n2726 ;
  assign n3926 = n3924 | n3925 ;
  assign n3927 = n761 | n3926 ;
  assign n3928 = n761 & n3926 ;
  assign n3929 = n3927 & ~n3928 ;
  assign n3930 = n2593 & n2848 ;
  assign n3931 = n2602 & n2918 ;
  assign n3932 = n2597 & n2846 ;
  assign n3933 = n3931 | n3932 ;
  assign n3934 = n3930 | n3933 ;
  assign n3935 = n2851 & n2898 ;
  assign n3936 = n3934 | n3935 ;
  assign n3937 = n516 & ~n2605 ;
  assign n3938 = n3936 & n3937 ;
  assign n3939 = n3936 | n3937 ;
  assign n3940 = ~n3938 & n3939 ;
  assign n3941 = n516 & ~n2609 ;
  assign n3942 = ~n3781 & n3941 ;
  assign n3943 = n3784 | n3942 ;
  assign n3944 = ( n2940 & n3942 ) | ( n2940 & n3943 ) | ( n3942 & n3943 );
  assign n3945 = n3513 | n3942 ;
  assign n3946 = ( n3784 & n3942 ) | ( n3784 & n3945 ) | ( n3942 & n3945 );
  assign n3947 = ( n3773 & n3944 ) | ( n3773 & n3946 ) | ( n3944 & n3946 );
  assign n3948 = ~n3940 & n3947 ;
  assign n3949 = ( n2940 & n3513 ) | ( n2940 & n3773 ) | ( n3513 & n3773 );
  assign n3950 = n3929 & n3940 ;
  assign n3951 = ~n3943 & n3950 ;
  assign n3952 = n3929 & ~n3942 ;
  assign n3953 = n3940 & n3952 ;
  assign n3954 = ( ~n3949 & n3951 ) | ( ~n3949 & n3953 ) | ( n3951 & n3953 );
  assign n3955 = ( n3929 & n3948 ) | ( n3929 & n3954 ) | ( n3948 & n3954 );
  assign n3956 = n3940 & ~n3947 ;
  assign n3957 = n3948 | n3956 ;
  assign n3958 = ~n3929 & n3957 ;
  assign n3959 = ( n3929 & ~n3955 ) | ( n3929 & n3958 ) | ( ~n3955 & n3958 );
  assign n3960 = n3794 | n3959 ;
  assign n3961 = ~n3794 & n3960 ;
  assign n3962 = ( ~n3959 & n3960 ) | ( ~n3959 & n3961 ) | ( n3960 & n3961 );
  assign n3963 = n3919 & n3962 ;
  assign n3964 = n3919 & ~n3963 ;
  assign n3965 = ~n3919 & n3962 ;
  assign n3966 = n3964 | n3965 ;
  assign n3967 = n3797 & n3965 ;
  assign n3968 = ( n3797 & n3964 ) | ( n3797 & n3967 ) | ( n3964 & n3967 );
  assign n3969 = ( n3804 & n3966 ) | ( n3804 & n3968 ) | ( n3966 & n3968 );
  assign n3970 = ( n3807 & n3966 ) | ( n3807 & n3968 ) | ( n3966 & n3968 );
  assign n3971 = ( n3042 & n3969 ) | ( n3042 & n3970 ) | ( n3969 & n3970 );
  assign n3972 = n3797 | n3965 ;
  assign n3973 = n3964 | n3972 ;
  assign n3974 = n3804 | n3973 ;
  assign n3975 = n3807 | n3973 ;
  assign n3976 = ( n3042 & n3974 ) | ( n3042 & n3975 ) | ( n3974 & n3975 );
  assign n3977 = ~n3971 & n3976 ;
  assign n3978 = n2555 & n3013 ;
  assign n3979 = n2655 & n3019 ;
  assign n3980 = ~n2550 & n3021 ;
  assign n3981 = n3979 | n3980 ;
  assign n3982 = n3978 | n3981 ;
  assign n3983 = n3028 & ~n3248 ;
  assign n3984 = n3982 | n3983 ;
  assign n3985 = n1238 | n3984 ;
  assign n3986 = n1238 & n3984 ;
  assign n3987 = n3985 & ~n3986 ;
  assign n3988 = ~n3977 & n3987 ;
  assign n3989 = n3977 & n3987 ;
  assign n3990 = n3977 & ~n3989 ;
  assign n3991 = ( n3574 & n3813 ) | ( n3574 & n3824 ) | ( n3813 & n3824 );
  assign n3992 = n3988 & n3991 ;
  assign n3993 = ( n3990 & n3991 ) | ( n3990 & n3992 ) | ( n3991 & n3992 );
  assign n3994 = n3813 | n3824 ;
  assign n3995 = n3988 & n3994 ;
  assign n3996 = ( n3990 & n3994 ) | ( n3990 & n3995 ) | ( n3994 & n3995 );
  assign n3997 = ( n3581 & n3993 ) | ( n3581 & n3996 ) | ( n3993 & n3996 );
  assign n3998 = ( n3581 & n3991 ) | ( n3581 & n3994 ) | ( n3991 & n3994 );
  assign n3999 = ( n3977 & ~n3987 ) | ( n3977 & n3998 ) | ( ~n3987 & n3998 );
  assign n4000 = ( n3988 & ~n3997 ) | ( n3988 & n3999 ) | ( ~n3997 & n3999 );
  assign n4001 = n3908 & n4000 ;
  assign n4002 = n3908 & ~n4001 ;
  assign n4003 = ~n3908 & n4000 ;
  assign n4004 = n4002 | n4003 ;
  assign n4005 = n3828 | n3832 ;
  assign n4006 = n4004 | n4005 ;
  assign n4007 = n4004 & n4005 ;
  assign n4008 = n4006 & ~n4007 ;
  assign n4009 = n3865 | n4008 ;
  assign n4010 = n3865 & n4008 ;
  assign n4011 = n4009 & ~n4010 ;
  assign n4012 = n3689 | n3702 ;
  assign n4013 = n3621 | n3702 ;
  assign n4014 = ( n3585 & n4012 ) | ( n3585 & n4013 ) | ( n4012 & n4013 );
  assign n4015 = ( n3835 & n3839 ) | ( n3835 & n4014 ) | ( n3839 & n4014 );
  assign n4016 = ( n3837 & n3838 ) | ( n3837 & n4015 ) | ( n3838 & n4015 );
  assign n4017 = n4011 & n4016 ;
  assign n4018 = n4011 | n4016 ;
  assign n4019 = ~n4017 & n4018 ;
  assign n4020 = n3843 & n4019 ;
  assign n4021 = n3843 | n4019 ;
  assign n4022 = ~n4020 & n4021 ;
  assign n4023 = n3849 & ~n4022 ;
  assign n4024 = ~n3849 & n4022 ;
  assign n4025 = n4023 | n4024 ;
  assign n4026 = n216 | n425 ;
  assign n4027 = n654 | n4026 ;
  assign n4028 = n206 | n2037 ;
  assign n4029 = n224 | n4028 ;
  assign n4030 = n281 | n4029 ;
  assign n4031 = n321 | n4030 ;
  assign n4032 = n358 | n4031 ;
  assign n4033 = n4027 | n4032 ;
  assign n4034 = n3670 | n4033 ;
  assign n4035 = n287 | n4034 ;
  assign n4036 = n142 | n4035 ;
  assign n4037 = n112 | n4036 ;
  assign n4038 = n389 | n4037 ;
  assign n4039 = n315 | n4038 ;
  assign n4040 = n234 | n4039 ;
  assign n4041 = n394 | n4040 ;
  assign n4042 = n4010 | n4016 ;
  assign n4043 = ( n4010 & n4011 ) | ( n4010 & n4042 ) | ( n4011 & n4042 );
  assign n4044 = n2697 & n3494 ;
  assign n4045 = n2655 & n2685 ;
  assign n4046 = ~n2570 & n2693 ;
  assign n4047 = n2567 & n2690 ;
  assign n4048 = n4046 | n4047 ;
  assign n4049 = n4045 | n4048 ;
  assign n4050 = n4044 | n4049 ;
  assign n4051 = n969 & n4050 ;
  assign n4052 = n4050 & ~n4051 ;
  assign n4053 = n969 & ~n4051 ;
  assign n4054 = n4052 | n4053 ;
  assign n4055 = ~n2590 & n2848 ;
  assign n4056 = n2597 & n2918 ;
  assign n4057 = n2593 & n2846 ;
  assign n4058 = n4056 | n4057 ;
  assign n4059 = n4055 | n4058 ;
  assign n4060 = n2851 & ~n2882 ;
  assign n4061 = n4059 | n4060 ;
  assign n4062 = n516 & ~n2602 ;
  assign n4063 = n4061 & n4062 ;
  assign n4064 = n4061 | n4062 ;
  assign n4065 = ~n4063 & n4064 ;
  assign n4066 = n516 & ~n3936 ;
  assign n4067 = n2605 & n4066 ;
  assign n4068 = n3940 | n4067 ;
  assign n4069 = ( n3943 & n4067 ) | ( n3943 & n4068 ) | ( n4067 & n4068 );
  assign n4070 = n4065 & n4069 ;
  assign n4071 = n3942 | n4067 ;
  assign n4072 = ( n3940 & n4067 ) | ( n3940 & n4071 ) | ( n4067 & n4071 );
  assign n4073 = n4065 & n4072 ;
  assign n4074 = ( n3949 & n4070 ) | ( n3949 & n4073 ) | ( n4070 & n4073 );
  assign n4075 = n4065 & ~n4074 ;
  assign n4076 = n2574 & n2720 ;
  assign n4077 = n2584 & n2818 ;
  assign n4078 = n2580 & n2715 ;
  assign n4079 = n4077 | n4078 ;
  assign n4080 = n4076 | n4079 ;
  assign n4081 = n2726 & n3060 ;
  assign n4082 = n4080 | n4081 ;
  assign n4083 = n761 | n4082 ;
  assign n4084 = n761 & n4082 ;
  assign n4085 = n4083 & ~n4084 ;
  assign n4086 = ~n4074 & n4085 ;
  assign n4087 = n4069 & n4085 ;
  assign n4088 = n4072 & n4085 ;
  assign n4089 = ( n3949 & n4087 ) | ( n3949 & n4088 ) | ( n4087 & n4088 );
  assign n4090 = ( n4075 & n4086 ) | ( n4075 & n4089 ) | ( n4086 & n4089 );
  assign n4091 = n4074 & ~n4085 ;
  assign n4092 = n4069 | n4085 ;
  assign n4093 = n4072 | n4085 ;
  assign n4094 = ( n3949 & n4092 ) | ( n3949 & n4093 ) | ( n4092 & n4093 );
  assign n4095 = ( n4075 & ~n4091 ) | ( n4075 & n4094 ) | ( ~n4091 & n4094 );
  assign n4096 = ~n4090 & n4095 ;
  assign n4097 = n3929 | n3955 ;
  assign n4098 = n3958 | n4097 ;
  assign n4099 = n4096 & n4098 ;
  assign n4100 = n3955 & n4096 ;
  assign n4101 = ( n3794 & n4099 ) | ( n3794 & n4100 ) | ( n4099 & n4100 );
  assign n4102 = ( n3794 & n3955 ) | ( n3794 & n4098 ) | ( n3955 & n4098 );
  assign n4103 = n4096 | n4102 ;
  assign n4104 = ~n4101 & n4103 ;
  assign n4105 = n4054 & n4104 ;
  assign n4106 = n4054 & ~n4105 ;
  assign n4107 = ~n4054 & n4104 ;
  assign n4108 = n4106 | n4107 ;
  assign n4109 = n3963 | n3968 ;
  assign n4110 = n3963 | n3965 ;
  assign n4111 = n3964 | n4110 ;
  assign n4112 = ( n3804 & n4109 ) | ( n3804 & n4111 ) | ( n4109 & n4111 );
  assign n4113 = ( n3807 & n4109 ) | ( n3807 & n4111 ) | ( n4109 & n4111 );
  assign n4114 = ( n3042 & n4112 ) | ( n3042 & n4113 ) | ( n4112 & n4113 );
  assign n4115 = n4108 | n4114 ;
  assign n4116 = n4108 & n4114 ;
  assign n4117 = n4115 & ~n4116 ;
  assign n4118 = n2540 & n3013 ;
  assign n4119 = ~n2550 & n3019 ;
  assign n4120 = n2555 & n3021 ;
  assign n4121 = n4119 | n4120 ;
  assign n4122 = n4118 | n4121 ;
  assign n4123 = n2672 & n3028 ;
  assign n4124 = n4122 | n4123 ;
  assign n4125 = n1238 | n4124 ;
  assign n4126 = n1238 & n4124 ;
  assign n4127 = n4125 & ~n4126 ;
  assign n4128 = ~n4117 & n4127 ;
  assign n4129 = n4117 & ~n4127 ;
  assign n4130 = n4128 | n4129 ;
  assign n4131 = n3989 & ~n4130 ;
  assign n4132 = ( n3993 & ~n4130 ) | ( n3993 & n4131 ) | ( ~n4130 & n4131 );
  assign n4133 = ( n3996 & ~n4130 ) | ( n3996 & n4131 ) | ( ~n4130 & n4131 );
  assign n4134 = ( n3581 & n4132 ) | ( n3581 & n4133 ) | ( n4132 & n4133 );
  assign n4135 = n3989 | n3997 ;
  assign n4136 = n4130 | n4134 ;
  assign n4137 = ( n4134 & ~n4135 ) | ( n4134 & n4136 ) | ( ~n4135 & n4136 );
  assign n4138 = n4001 | n4007 ;
  assign n4139 = n2551 & ~n3725 ;
  assign n4140 = n2556 & ~n3886 ;
  assign n4141 = n4139 | n4140 ;
  assign n4142 = ( n3886 & n3887 ) | ( n3886 & ~n3896 ) | ( n3887 & ~n3896 );
  assign n4143 = n3886 & ~n3896 ;
  assign n4144 = n4142 & ~n4143 ;
  assign n4145 = n2673 & n4144 ;
  assign n4146 = n4141 | n4145 ;
  assign n4147 = n32 & n4146 ;
  assign n4148 = n4146 & ~n4147 ;
  assign n4149 = n32 & ~n4147 ;
  assign n4150 = n4148 | n4149 ;
  assign n4151 = ( ~n4137 & n4138 ) | ( ~n4137 & n4150 ) | ( n4138 & n4150 );
  assign n4152 = ( n4138 & n4150 ) | ( n4138 & ~n4151 ) | ( n4150 & ~n4151 );
  assign n4153 = ( n4137 & n4151 ) | ( n4137 & ~n4152 ) | ( n4151 & ~n4152 );
  assign n4154 = ( n4041 & n4043 ) | ( n4041 & ~n4153 ) | ( n4043 & ~n4153 );
  assign n4155 = ( ~n4043 & n4153 ) | ( ~n4043 & n4154 ) | ( n4153 & n4154 );
  assign n4156 = ( ~n4041 & n4154 ) | ( ~n4041 & n4155 ) | ( n4154 & n4155 );
  assign n4157 = n4020 | n4156 ;
  assign n4158 = n4020 & n4156 ;
  assign n4159 = n4157 & ~n4158 ;
  assign n4160 = n3845 | n4022 ;
  assign n4161 = n3848 & n4160 ;
  assign n4162 = ~n4159 & n4161 ;
  assign n4163 = n4159 & ~n4161 ;
  assign n4164 = n4162 | n4163 ;
  assign n4165 = n4159 | n4160 ;
  assign n4166 = n3848 & n4165 ;
  assign n4167 = n4041 | n4153 ;
  assign n4168 = n4041 & n4153 ;
  assign n4169 = ( n3865 & n4041 ) | ( n3865 & n4153 ) | ( n4041 & n4153 );
  assign n4170 = ( n4008 & n4168 ) | ( n4008 & n4169 ) | ( n4168 & n4169 );
  assign n4171 = ( n4016 & n4167 ) | ( n4016 & n4170 ) | ( n4167 & n4170 );
  assign n4172 = n4167 & n4169 ;
  assign n4173 = n4167 & n4168 ;
  assign n4174 = ( n4008 & n4172 ) | ( n4008 & n4173 ) | ( n4172 & n4173 );
  assign n4175 = ( n4011 & n4171 ) | ( n4011 & n4174 ) | ( n4171 & n4174 );
  assign n4176 = n2251 | n3625 ;
  assign n4177 = n291 | n4176 ;
  assign n4178 = n900 | n4177 ;
  assign n4179 = n2086 | n4178 ;
  assign n4180 = n1375 | n4179 ;
  assign n4181 = n713 | n4180 ;
  assign n4182 = n444 | n4181 ;
  assign n4183 = n259 | n4182 ;
  assign n4184 = n267 | n4183 ;
  assign n4185 = n333 | n4184 ;
  assign n4186 = n124 | n4185 ;
  assign n4187 = n101 | n4186 ;
  assign n4188 = n2551 & ~n3886 ;
  assign n4189 = n2673 & ~n4142 ;
  assign n4190 = n4188 | n4189 ;
  assign n4191 = n32 & n4190 ;
  assign n4192 = n4190 & ~n4191 ;
  assign n4193 = n32 & ~n4191 ;
  assign n4194 = n4192 | n4193 ;
  assign n4195 = n4090 | n4101 ;
  assign n4196 = ~n2570 & n2720 ;
  assign n4197 = n2580 & n2818 ;
  assign n4198 = n2574 & n2715 ;
  assign n4199 = n4197 | n4198 ;
  assign n4200 = n4196 | n4199 ;
  assign n4201 = n2726 & ~n3228 ;
  assign n4202 = n4200 | n4201 ;
  assign n4203 = n761 | n4202 ;
  assign n4204 = n761 & n4202 ;
  assign n4205 = n4203 & ~n4204 ;
  assign n4206 = n516 & ~n4061 ;
  assign n4207 = n2602 & n4206 ;
  assign n4208 = n4065 | n4207 ;
  assign n4209 = ( n4069 & n4207 ) | ( n4069 & n4208 ) | ( n4207 & n4208 );
  assign n4210 = ( n4072 & n4207 ) | ( n4072 & n4208 ) | ( n4207 & n4208 );
  assign n4211 = ( n3949 & n4209 ) | ( n3949 & n4210 ) | ( n4209 & n4210 );
  assign n4212 = n516 & ~n2597 ;
  assign n4213 = n2584 & n2848 ;
  assign n4214 = n2593 & n2918 ;
  assign n4215 = ~n2590 & n2846 ;
  assign n4216 = n4214 | n4215 ;
  assign n4217 = n4213 | n4216 ;
  assign n4218 = n2851 & ~n2988 ;
  assign n4219 = n4217 | n4218 ;
  assign n4220 = n4212 & n4219 ;
  assign n4221 = n4212 | n4219 ;
  assign n4222 = ~n4220 & n4221 ;
  assign n4223 = n4208 & n4222 ;
  assign n4224 = n4207 & n4222 ;
  assign n4225 = ( n4069 & n4223 ) | ( n4069 & n4224 ) | ( n4223 & n4224 );
  assign n4226 = ( n4072 & n4223 ) | ( n4072 & n4224 ) | ( n4223 & n4224 );
  assign n4227 = ( n3949 & n4225 ) | ( n3949 & n4226 ) | ( n4225 & n4226 );
  assign n4228 = n4211 & ~n4227 ;
  assign n4229 = n4222 & ~n4224 ;
  assign n4230 = ~n4208 & n4222 ;
  assign n4231 = ( ~n4069 & n4229 ) | ( ~n4069 & n4230 ) | ( n4229 & n4230 );
  assign n4232 = ( ~n4072 & n4229 ) | ( ~n4072 & n4230 ) | ( n4229 & n4230 );
  assign n4233 = ( ~n3949 & n4231 ) | ( ~n3949 & n4232 ) | ( n4231 & n4232 );
  assign n4234 = n4205 & n4233 ;
  assign n4235 = ( n4205 & n4228 ) | ( n4205 & n4234 ) | ( n4228 & n4234 );
  assign n4236 = n4205 | n4233 ;
  assign n4237 = n4228 | n4236 ;
  assign n4238 = ~n4235 & n4237 ;
  assign n4239 = n4195 | n4238 ;
  assign n4240 = n4195 & n4238 ;
  assign n4241 = n4239 & ~n4240 ;
  assign n4242 = ~n2550 & n2685 ;
  assign n4243 = n2567 & n2693 ;
  assign n4244 = n2655 & n2690 ;
  assign n4245 = n4243 | n4244 ;
  assign n4246 = n4242 | n4245 ;
  assign n4247 = n2697 & ~n3264 ;
  assign n4248 = n4246 | n4247 ;
  assign n4249 = n969 & n4248 ;
  assign n4250 = n4248 & ~n4249 ;
  assign n4251 = n969 & ~n4249 ;
  assign n4252 = n4250 | n4251 ;
  assign n4253 = n4241 & ~n4252 ;
  assign n4254 = ~n4241 & n4252 ;
  assign n4255 = n4253 | n4254 ;
  assign n4256 = n4054 | n4255 ;
  assign n4257 = n4104 | n4255 ;
  assign n4258 = ( n4114 & n4256 ) | ( n4114 & n4257 ) | ( n4256 & n4257 );
  assign n4259 = n4054 & n4255 ;
  assign n4260 = n4104 & n4255 ;
  assign n4261 = ( n4114 & n4259 ) | ( n4114 & n4260 ) | ( n4259 & n4260 );
  assign n4262 = n4258 & ~n4261 ;
  assign n4263 = n3028 & ~n3738 ;
  assign n4264 = n3028 & n3740 ;
  assign n4265 = ( ~n3739 & n4263 ) | ( ~n3739 & n4264 ) | ( n4263 & n4264 );
  assign n4266 = n3013 & ~n3725 ;
  assign n4267 = n2555 & n3019 ;
  assign n4268 = n2540 & n3021 ;
  assign n4269 = n4267 | n4268 ;
  assign n4270 = n4266 | n4269 ;
  assign n4271 = n1238 | n4270 ;
  assign n4272 = n4265 | n4271 ;
  assign n4273 = n1238 & n4270 ;
  assign n4274 = ( n1238 & n4265 ) | ( n1238 & n4273 ) | ( n4265 & n4273 );
  assign n4275 = n4272 & ~n4274 ;
  assign n4276 = n4262 & n4275 ;
  assign n4277 = n4262 | n4275 ;
  assign n4278 = ~n4276 & n4277 ;
  assign n4279 = n4194 & n4278 ;
  assign n4280 = n4194 | n4278 ;
  assign n4281 = ~n4279 & n4280 ;
  assign n4282 = ( n3989 & n4117 ) | ( n3989 & n4127 ) | ( n4117 & n4127 );
  assign n4283 = n4117 | n4127 ;
  assign n4284 = ( n3997 & n4282 ) | ( n3997 & n4283 ) | ( n4282 & n4283 );
  assign n4285 = n4281 & n4284 ;
  assign n4286 = n4281 | n4284 ;
  assign n4287 = ~n4285 & n4286 ;
  assign n4288 = ( n4134 & n4138 ) | ( n4134 & n4150 ) | ( n4138 & n4150 );
  assign n4289 = ( ~n3989 & n4138 ) | ( ~n3989 & n4150 ) | ( n4138 & n4150 );
  assign n4290 = n4138 & n4150 ;
  assign n4291 = ( ~n3997 & n4289 ) | ( ~n3997 & n4290 ) | ( n4289 & n4290 );
  assign n4292 = ( n4136 & n4288 ) | ( n4136 & n4291 ) | ( n4288 & n4291 );
  assign n4293 = n4287 | n4292 ;
  assign n4294 = n4287 & n4292 ;
  assign n4295 = n4293 & ~n4294 ;
  assign n4296 = n123 | n4295 ;
  assign n4297 = n4187 | n4296 ;
  assign n4298 = n123 & n4295 ;
  assign n4299 = ( n4187 & n4295 ) | ( n4187 & n4298 ) | ( n4295 & n4298 );
  assign n4300 = n4297 & ~n4299 ;
  assign n4301 = n4175 | n4300 ;
  assign n4302 = n4175 & ~n4300 ;
  assign n4303 = ( ~n4175 & n4301 ) | ( ~n4175 & n4302 ) | ( n4301 & n4302 );
  assign n4304 = n4020 & n4303 ;
  assign n4305 = n4156 & n4304 ;
  assign n4306 = n4020 | n4303 ;
  assign n4307 = ( n4156 & n4303 ) | ( n4156 & n4306 ) | ( n4303 & n4306 );
  assign n4308 = ~n4305 & n4307 ;
  assign n4309 = n4166 & n4308 ;
  assign n4310 = n4166 | n4308 ;
  assign n4311 = ~n4309 & n4310 ;
  assign n4312 = n550 | n2037 ;
  assign n4313 = n659 | n4312 ;
  assign n4314 = n954 | n4313 ;
  assign n4315 = n2383 | n4314 ;
  assign n4316 = n357 | n729 ;
  assign n4317 = n4315 | n4316 ;
  assign n4318 = n247 | n264 ;
  assign n4319 = n4317 | n4318 ;
  assign n4320 = n262 | n4319 ;
  assign n4321 = n143 | n4320 ;
  assign n4322 = n2580 & n2848 ;
  assign n4323 = ~n2590 & n2918 ;
  assign n4324 = n2584 & n2846 ;
  assign n4325 = n4323 | n4324 ;
  assign n4326 = n4322 | n4325 ;
  assign n4327 = n2701 & n2851 ;
  assign n4328 = n4326 | n4327 ;
  assign n4329 = n516 & ~n4328 ;
  assign n4330 = n516 & ~n4329 ;
  assign n4331 = ( n4328 & n4329 ) | ( n4328 & ~n4330 ) | ( n4329 & ~n4330 );
  assign n4332 = n32 & n516 ;
  assign n4333 = n2593 & n4332 ;
  assign n4334 = n32 & ~n4333 ;
  assign n4335 = n2593 & ~n4333 ;
  assign n4336 = n516 & n4335 ;
  assign n4337 = n4334 | n4336 ;
  assign n4338 = n4331 & n4337 ;
  assign n4339 = n4331 & ~n4338 ;
  assign n4340 = n4337 & ~n4338 ;
  assign n4341 = n4339 | n4340 ;
  assign n4342 = n516 & n2597 ;
  assign n4343 = ( ~n4219 & n4227 ) | ( ~n4219 & n4342 ) | ( n4227 & n4342 );
  assign n4344 = n2567 & n2720 ;
  assign n4345 = n2574 & n2818 ;
  assign n4346 = ~n2570 & n2715 ;
  assign n4347 = n4345 | n4346 ;
  assign n4348 = n4344 | n4347 ;
  assign n4349 = n2726 & ~n3027 ;
  assign n4350 = n4348 | n4349 ;
  assign n4351 = n761 & n4350 ;
  assign n4352 = n761 | n4350 ;
  assign n4353 = ~n4351 & n4352 ;
  assign n4354 = ( n4227 & n4341 ) | ( n4227 & ~n4353 ) | ( n4341 & ~n4353 );
  assign n4355 = ~n4341 & n4353 ;
  assign n4356 = ( n4343 & n4354 ) | ( n4343 & ~n4355 ) | ( n4354 & ~n4355 );
  assign n4357 = n4227 | n4343 ;
  assign n4358 = ( n4353 & n4356 ) | ( n4353 & ~n4357 ) | ( n4356 & ~n4357 );
  assign n4359 = ( ~n4341 & n4356 ) | ( ~n4341 & n4358 ) | ( n4356 & n4358 );
  assign n4360 = n4090 | n4235 ;
  assign n4361 = ( n4235 & n4238 ) | ( n4235 & n4360 ) | ( n4238 & n4360 );
  assign n4362 = ~n4359 & n4361 ;
  assign n4363 = n4235 | n4238 ;
  assign n4364 = ~n4359 & n4363 ;
  assign n4365 = ( n4101 & n4362 ) | ( n4101 & n4364 ) | ( n4362 & n4364 );
  assign n4366 = n4359 | n4365 ;
  assign n4367 = n2555 & n2685 ;
  assign n4368 = n2655 & n2693 ;
  assign n4369 = ~n2550 & n2690 ;
  assign n4370 = n4368 | n4369 ;
  assign n4371 = n4367 | n4370 ;
  assign n4372 = n2697 & ~n3245 ;
  assign n4373 = ~n2555 & n2697 ;
  assign n4374 = ( n3247 & n4372 ) | ( n3247 & n4373 ) | ( n4372 & n4373 );
  assign n4375 = n4371 | n4374 ;
  assign n4376 = n969 & ~n4371 ;
  assign n4377 = ~n4374 & n4376 ;
  assign n4378 = n969 & ~n4376 ;
  assign n4379 = ( n969 & n4374 ) | ( n969 & n4378 ) | ( n4374 & n4378 );
  assign n4380 = ( n4375 & n4377 ) | ( n4375 & ~n4379 ) | ( n4377 & ~n4379 );
  assign n4381 = n4365 & n4380 ;
  assign n4382 = ~n4361 & n4380 ;
  assign n4383 = ~n4363 & n4380 ;
  assign n4384 = ( ~n4101 & n4382 ) | ( ~n4101 & n4383 ) | ( n4382 & n4383 );
  assign n4385 = ( n4366 & n4381 ) | ( n4366 & n4384 ) | ( n4381 & n4384 );
  assign n4386 = n4365 | n4380 ;
  assign n4387 = ( n4101 & n4361 ) | ( n4101 & n4363 ) | ( n4361 & n4363 );
  assign n4388 = ~n4380 & n4387 ;
  assign n4389 = ( n4366 & n4386 ) | ( n4366 & ~n4388 ) | ( n4386 & ~n4388 );
  assign n4390 = ~n4385 & n4389 ;
  assign n4391 = n4241 | n4390 ;
  assign n4392 = ( n4252 & n4390 ) | ( n4252 & n4391 ) | ( n4390 & n4391 );
  assign n4393 = n4260 | n4392 ;
  assign n4394 = n4259 | n4392 ;
  assign n4395 = ( n4114 & n4393 ) | ( n4114 & n4394 ) | ( n4393 & n4394 );
  assign n4396 = n4105 | n4107 ;
  assign n4397 = n4106 | n4396 ;
  assign n4398 = ( n4241 & n4252 ) | ( n4241 & n4397 ) | ( n4252 & n4397 );
  assign n4399 = n4390 & n4398 ;
  assign n4400 = ( n4105 & n4241 ) | ( n4105 & n4252 ) | ( n4241 & n4252 );
  assign n4401 = n4390 & n4400 ;
  assign n4402 = ( n4114 & n4399 ) | ( n4114 & n4401 ) | ( n4399 & n4401 );
  assign n4403 = n4395 & ~n4402 ;
  assign n4404 = n3013 & ~n3886 ;
  assign n4405 = n2540 & n3019 ;
  assign n4406 = n3021 & ~n3725 ;
  assign n4407 = n4405 | n4406 ;
  assign n4408 = n4404 | n4407 ;
  assign n4409 = n3028 & n3897 ;
  assign n4410 = n4408 | n4409 ;
  assign n4411 = n1238 & n4410 ;
  assign n4412 = n1238 | n4410 ;
  assign n4413 = ~n4411 & n4412 ;
  assign n4414 = n4403 & n4413 ;
  assign n4415 = n4403 | n4413 ;
  assign n4416 = ~n4414 & n4415 ;
  assign n4417 = n4194 | n4276 ;
  assign n4418 = ( n4276 & n4278 ) | ( n4276 & n4417 ) | ( n4278 & n4417 );
  assign n4419 = n4416 & n4418 ;
  assign n4420 = n4416 | n4418 ;
  assign n4421 = ~n4419 & n4420 ;
  assign n4422 = n4285 | n4421 ;
  assign n4423 = n4287 | n4422 ;
  assign n4424 = ( n4292 & n4422 ) | ( n4292 & n4423 ) | ( n4422 & n4423 );
  assign n4425 = ( n4285 & n4287 ) | ( n4285 & n4421 ) | ( n4287 & n4421 );
  assign n4426 = n4285 & n4421 ;
  assign n4427 = ( n4292 & n4425 ) | ( n4292 & n4426 ) | ( n4425 & n4426 );
  assign n4428 = n4424 & ~n4427 ;
  assign n4429 = n4321 | n4428 ;
  assign n4430 = n4321 & n4428 ;
  assign n4431 = n4429 & ~n4430 ;
  assign n4432 = n123 | n4187 ;
  assign n4433 = ( n4168 & n4295 ) | ( n4168 & n4432 ) | ( n4295 & n4432 );
  assign n4434 = n4431 | n4433 ;
  assign n4435 = ( n4167 & n4295 ) | ( n4167 & n4432 ) | ( n4295 & n4432 );
  assign n4436 = n4434 | n4435 ;
  assign n4437 = n4433 & n4435 ;
  assign n4438 = n4431 | n4437 ;
  assign n4439 = ( n3865 & n4433 ) | ( n3865 & n4435 ) | ( n4433 & n4435 );
  assign n4440 = n4431 | n4439 ;
  assign n4441 = ( n4008 & n4438 ) | ( n4008 & n4440 ) | ( n4438 & n4440 );
  assign n4442 = ( n4016 & n4436 ) | ( n4016 & n4441 ) | ( n4436 & n4441 );
  assign n4443 = n4436 & n4440 ;
  assign n4444 = n4436 & n4438 ;
  assign n4445 = ( n4008 & n4443 ) | ( n4008 & n4444 ) | ( n4443 & n4444 );
  assign n4446 = ( n4011 & n4442 ) | ( n4011 & n4445 ) | ( n4442 & n4445 );
  assign n4447 = n4431 & n4433 ;
  assign n4448 = ( n4431 & n4435 ) | ( n4431 & n4447 ) | ( n4435 & n4447 );
  assign n4449 = n4431 & n4437 ;
  assign n4450 = n4431 & n4439 ;
  assign n4451 = ( n4008 & n4449 ) | ( n4008 & n4450 ) | ( n4449 & n4450 );
  assign n4452 = ( n4016 & n4448 ) | ( n4016 & n4451 ) | ( n4448 & n4451 );
  assign n4453 = n4448 & n4450 ;
  assign n4454 = n4448 & n4449 ;
  assign n4455 = ( n4008 & n4453 ) | ( n4008 & n4454 ) | ( n4453 & n4454 );
  assign n4456 = ( n4011 & n4452 ) | ( n4011 & n4455 ) | ( n4452 & n4455 );
  assign n4457 = n4446 & ~n4456 ;
  assign n4458 = n4305 | n4457 ;
  assign n4459 = ( ~n4020 & n4303 ) | ( ~n4020 & n4457 ) | ( n4303 & n4457 );
  assign n4460 = n4303 | n4457 ;
  assign n4461 = ( ~n4156 & n4459 ) | ( ~n4156 & n4460 ) | ( n4459 & n4460 );
  assign n4462 = n4158 & n4461 ;
  assign n4463 = n4458 & ~n4462 ;
  assign n4464 = n3848 & n4308 ;
  assign n4465 = ( n3848 & n4165 ) | ( n3848 & n4464 ) | ( n4165 & n4464 );
  assign n4466 = ~n4463 & n4465 ;
  assign n4467 = n4463 & ~n4465 ;
  assign n4468 = n4466 | n4467 ;
  assign n4469 = n4165 | n4308 ;
  assign n4470 = n3848 & n4463 ;
  assign n4471 = ( n3848 & n4469 ) | ( n3848 & n4470 ) | ( n4469 & n4470 );
  assign n4472 = n346 | n3872 ;
  assign n4473 = n186 | n668 ;
  assign n4474 = n259 | n459 ;
  assign n4475 = n170 | n4474 ;
  assign n4476 = n4473 | n4475 ;
  assign n4477 = n2227 | n4476 ;
  assign n4478 = n288 | n4477 ;
  assign n4479 = n4472 | n4478 ;
  assign n4480 = n2498 | n4479 ;
  assign n4481 = n3855 | n4480 ;
  assign n4482 = n2024 | n4481 ;
  assign n4483 = n264 | n4482 ;
  assign n4484 = n189 | n4483 ;
  assign n4485 = n203 | n4484 ;
  assign n4486 = n96 | n4485 ;
  assign n4487 = n4419 | n4427 ;
  assign n4488 = n4402 | n4414 ;
  assign n4489 = n2726 & n3494 ;
  assign n4490 = n2655 & n2720 ;
  assign n4491 = ~n2570 & n2818 ;
  assign n4492 = n2567 & n2715 ;
  assign n4493 = n4491 | n4492 ;
  assign n4494 = n4490 | n4493 ;
  assign n4495 = n4489 | n4494 ;
  assign n4496 = n761 | n4495 ;
  assign n4497 = n761 & n4495 ;
  assign n4498 = n4496 & ~n4497 ;
  assign n4499 = n4333 | n4338 ;
  assign n4500 = ~n2590 & n4332 ;
  assign n4501 = n32 & ~n4500 ;
  assign n4502 = n2590 | n4500 ;
  assign n4503 = n516 & ~n4502 ;
  assign n4504 = n4501 | n4503 ;
  assign n4505 = n4499 & n4504 ;
  assign n4506 = n4499 & ~n4505 ;
  assign n4507 = n4504 & ~n4505 ;
  assign n4508 = n4506 | n4507 ;
  assign n4509 = n2574 & n2848 ;
  assign n4510 = n2584 & n2918 ;
  assign n4511 = n2580 & n2846 ;
  assign n4512 = n4510 | n4511 ;
  assign n4513 = n4509 | n4512 ;
  assign n4514 = n2851 & n3060 ;
  assign n4515 = n4513 | n4514 ;
  assign n4516 = n516 | n4515 ;
  assign n4517 = n516 & n4515 ;
  assign n4518 = n4516 & ~n4517 ;
  assign n4519 = ( ~n4498 & n4508 ) | ( ~n4498 & n4518 ) | ( n4508 & n4518 );
  assign n4520 = ( n4498 & n4508 ) | ( n4498 & n4518 ) | ( n4508 & n4518 );
  assign n4521 = ( n4498 & n4519 ) | ( n4498 & ~n4520 ) | ( n4519 & ~n4520 );
  assign n4522 = ~n4219 & n4342 ;
  assign n4523 = n4227 | n4522 ;
  assign n4524 = ( n4341 & n4353 ) | ( n4341 & n4523 ) | ( n4353 & n4523 );
  assign n4525 = n2672 & n2697 ;
  assign n4526 = n2540 & n2685 ;
  assign n4527 = ~n2550 & n2693 ;
  assign n4528 = n2555 & n2690 ;
  assign n4529 = n4527 | n4528 ;
  assign n4530 = n4526 | n4529 ;
  assign n4531 = n4525 | n4530 ;
  assign n4532 = n969 & ~n4531 ;
  assign n4533 = n969 & ~n4532 ;
  assign n4534 = ( n4531 & n4532 ) | ( n4531 & ~n4533 ) | ( n4532 & ~n4533 );
  assign n4535 = ( n4521 & ~n4524 ) | ( n4521 & n4534 ) | ( ~n4524 & n4534 );
  assign n4536 = ( n4521 & n4524 ) | ( n4521 & ~n4534 ) | ( n4524 & ~n4534 );
  assign n4537 = ( ~n4521 & n4535 ) | ( ~n4521 & n4536 ) | ( n4535 & n4536 );
  assign n4538 = ( n4100 & n4361 ) | ( n4100 & n4363 ) | ( n4361 & n4363 );
  assign n4539 = ( n4099 & n4361 ) | ( n4099 & n4363 ) | ( n4361 & n4363 );
  assign n4540 = ( n3794 & n4538 ) | ( n3794 & n4539 ) | ( n4538 & n4539 );
  assign n4541 = n4359 & n4540 ;
  assign n4542 = n4385 | n4541 ;
  assign n4543 = n3019 & ~n3725 ;
  assign n4544 = n3021 & ~n3886 ;
  assign n4545 = n4543 | n4544 ;
  assign n4546 = n3028 & n4144 ;
  assign n4547 = n4545 | n4546 ;
  assign n4548 = n1238 | n4547 ;
  assign n4549 = n1238 & n4547 ;
  assign n4550 = n4548 & ~n4549 ;
  assign n4551 = ( n4537 & n4542 ) | ( n4537 & n4550 ) | ( n4542 & n4550 );
  assign n4552 = ( ~n4537 & n4542 ) | ( ~n4537 & n4550 ) | ( n4542 & n4550 );
  assign n4553 = ( n4537 & ~n4551 ) | ( n4537 & n4552 ) | ( ~n4551 & n4552 );
  assign n4554 = n4488 & n4553 ;
  assign n4555 = n4488 | n4553 ;
  assign n4556 = ~n4554 & n4555 ;
  assign n4557 = n4487 & n4556 ;
  assign n4558 = n4487 | n4556 ;
  assign n4559 = ~n4557 & n4558 ;
  assign n4560 = n4486 | n4559 ;
  assign n4561 = n4486 & n4559 ;
  assign n4562 = n4560 & ~n4561 ;
  assign n4563 = n4430 | n4431 ;
  assign n4564 = ( n4430 & n4433 ) | ( n4430 & n4563 ) | ( n4433 & n4563 );
  assign n4565 = n4562 & n4564 ;
  assign n4566 = ( n4430 & n4435 ) | ( n4430 & n4563 ) | ( n4435 & n4563 );
  assign n4567 = n4562 & n4566 ;
  assign n4568 = n4565 | n4567 ;
  assign n4569 = ( n3865 & n4565 ) | ( n3865 & n4567 ) | ( n4565 & n4567 );
  assign n4570 = n4565 & n4567 ;
  assign n4571 = ( n4008 & n4569 ) | ( n4008 & n4570 ) | ( n4569 & n4570 );
  assign n4572 = ( n4016 & n4568 ) | ( n4016 & n4571 ) | ( n4568 & n4571 );
  assign n4573 = n4568 & n4570 ;
  assign n4574 = n4568 & n4569 ;
  assign n4575 = ( n4008 & n4573 ) | ( n4008 & n4574 ) | ( n4573 & n4574 );
  assign n4576 = ( n4011 & n4572 ) | ( n4011 & n4575 ) | ( n4572 & n4575 );
  assign n4577 = n4562 | n4564 ;
  assign n4578 = n4566 | n4577 ;
  assign n4579 = n4564 & n4566 ;
  assign n4580 = n4562 | n4579 ;
  assign n4581 = ( n3865 & n4564 ) | ( n3865 & n4566 ) | ( n4564 & n4566 );
  assign n4582 = n4562 | n4581 ;
  assign n4583 = ( n4008 & n4580 ) | ( n4008 & n4582 ) | ( n4580 & n4582 );
  assign n4584 = ( n4016 & n4578 ) | ( n4016 & n4583 ) | ( n4578 & n4583 );
  assign n4585 = n4578 & n4582 ;
  assign n4586 = n4578 & n4580 ;
  assign n4587 = ( n4008 & n4585 ) | ( n4008 & n4586 ) | ( n4585 & n4586 );
  assign n4588 = ( n4011 & n4584 ) | ( n4011 & n4587 ) | ( n4584 & n4587 );
  assign n4589 = ~n4576 & n4588 ;
  assign n4590 = n4457 & n4589 ;
  assign n4591 = n4305 & n4590 ;
  assign n4592 = n4462 | n4589 ;
  assign n4593 = ~n4591 & n4592 ;
  assign n4594 = n4471 & ~n4593 ;
  assign n4595 = n4471 | n4593 ;
  assign n4596 = ( ~n4471 & n4594 ) | ( ~n4471 & n4595 ) | ( n4594 & n4595 );
  assign n4597 = n4463 | n4593 ;
  assign n4598 = ( n3848 & n4465 ) | ( n3848 & n4597 ) | ( n4465 & n4597 );
  assign n4599 = n853 | n1027 ;
  assign n4600 = n477 | n4599 ;
  assign n4601 = n2345 | n4600 ;
  assign n4602 = n2251 | n4601 ;
  assign n4603 = n460 | n4602 ;
  assign n4604 = n2024 | n4603 ;
  assign n4605 = n121 | n4604 ;
  assign n4606 = n235 | n4605 ;
  assign n4607 = n947 | n3609 ;
  assign n4608 = n2377 | n4607 ;
  assign n4609 = n2523 | n4608 ;
  assign n4610 = n4606 | n4609 ;
  assign n4611 = n293 | n4610 ;
  assign n4612 = n180 | n4611 ;
  assign n4613 = n156 | n4612 ;
  assign n4614 = n418 | n4613 ;
  assign n4615 = n127 | n4614 ;
  assign n4616 = n126 | n4615 ;
  assign n4617 = n3019 & ~n3886 ;
  assign n4618 = n3028 & ~n4142 ;
  assign n4619 = n4617 | n4618 ;
  assign n4620 = ~n1238 & n4619 ;
  assign n4621 = n1238 & ~n4619 ;
  assign n4622 = n4620 | n4621 ;
  assign n4623 = n4524 & n4622 ;
  assign n4624 = n4534 & n4622 ;
  assign n4625 = ( n4521 & n4623 ) | ( n4521 & n4624 ) | ( n4623 & n4624 );
  assign n4626 = n4524 | n4622 ;
  assign n4627 = n4534 | n4622 ;
  assign n4628 = ( n4521 & n4626 ) | ( n4521 & n4627 ) | ( n4626 & n4627 );
  assign n4629 = ~n4625 & n4628 ;
  assign n4630 = n2685 & ~n3725 ;
  assign n4631 = n2555 & n2693 ;
  assign n4632 = n2540 & n2690 ;
  assign n4633 = n4631 | n4632 ;
  assign n4634 = n4630 | n4633 ;
  assign n4635 = ( n2697 & ~n3741 ) | ( n2697 & n4634 ) | ( ~n3741 & n4634 );
  assign n4636 = ( n969 & n4634 ) | ( n969 & ~n4635 ) | ( n4634 & ~n4635 );
  assign n4637 = n4635 | n4636 ;
  assign n4638 = ~n4634 & n4636 ;
  assign n4639 = ( ~n969 & n4637 ) | ( ~n969 & n4638 ) | ( n4637 & n4638 );
  assign n4640 = n2726 & ~n3264 ;
  assign n4641 = ~n2550 & n2720 ;
  assign n4642 = n2567 & n2818 ;
  assign n4643 = n2655 & n2715 ;
  assign n4644 = n4642 | n4643 ;
  assign n4645 = n4641 | n4644 ;
  assign n4646 = n4640 | n4645 ;
  assign n4647 = n761 | n4646 ;
  assign n4648 = n761 & n4646 ;
  assign n4649 = n4647 & ~n4648 ;
  assign n4650 = n4500 | n4505 ;
  assign n4651 = n2584 & n4332 ;
  assign n4652 = n32 & ~n4651 ;
  assign n4653 = n2584 & ~n4651 ;
  assign n4654 = n516 & n4653 ;
  assign n4655 = n4652 | n4654 ;
  assign n4656 = n4650 & n4655 ;
  assign n4657 = n4650 & ~n4656 ;
  assign n4658 = n4655 & ~n4656 ;
  assign n4659 = n4657 | n4658 ;
  assign n4660 = ~n2570 & n2848 ;
  assign n4661 = n2580 & n2918 ;
  assign n4662 = n2574 & n2846 ;
  assign n4663 = n4661 | n4662 ;
  assign n4664 = n4660 | n4663 ;
  assign n4665 = n2851 & ~n3228 ;
  assign n4666 = n4664 | n4665 ;
  assign n4667 = n516 | n4666 ;
  assign n4668 = n516 & n4666 ;
  assign n4669 = n4667 & ~n4668 ;
  assign n4670 = ( ~n4649 & n4659 ) | ( ~n4649 & n4669 ) | ( n4659 & n4669 );
  assign n4671 = ( n4649 & n4659 ) | ( n4649 & n4669 ) | ( n4659 & n4669 );
  assign n4672 = ( n4649 & n4670 ) | ( n4649 & ~n4671 ) | ( n4670 & ~n4671 );
  assign n4673 = ( n4520 & ~n4639 ) | ( n4520 & n4672 ) | ( ~n4639 & n4672 );
  assign n4674 = ( n4639 & ~n4672 ) | ( n4639 & n4673 ) | ( ~n4672 & n4673 );
  assign n4675 = ( ~n4520 & n4673 ) | ( ~n4520 & n4674 ) | ( n4673 & n4674 );
  assign n4676 = n4629 & n4675 ;
  assign n4677 = n4629 | n4675 ;
  assign n4678 = ~n4676 & n4677 ;
  assign n4679 = n4551 & n4678 ;
  assign n4680 = n4551 | n4678 ;
  assign n4681 = ~n4679 & n4680 ;
  assign n4682 = n4487 | n4488 ;
  assign n4683 = ( n4487 & n4553 ) | ( n4487 & n4682 ) | ( n4553 & n4682 );
  assign n4684 = ( n4554 & n4556 ) | ( n4554 & n4683 ) | ( n4556 & n4683 );
  assign n4685 = n4681 & n4684 ;
  assign n4686 = n4681 | n4684 ;
  assign n4687 = ~n4685 & n4686 ;
  assign n4688 = n4616 | n4687 ;
  assign n4689 = n4616 & n4687 ;
  assign n4690 = n4688 & ~n4689 ;
  assign n4691 = n4561 & n4690 ;
  assign n4692 = ( n4576 & n4690 ) | ( n4576 & n4691 ) | ( n4690 & n4691 );
  assign n4693 = n4561 | n4690 ;
  assign n4694 = n4576 | n4693 ;
  assign n4695 = ~n4692 & n4694 ;
  assign n4696 = n4590 & n4695 ;
  assign n4697 = n4305 & n4696 ;
  assign n4698 = n4590 | n4695 ;
  assign n4699 = ( n4305 & n4695 ) | ( n4305 & n4698 ) | ( n4695 & n4698 );
  assign n4700 = ~n4697 & n4699 ;
  assign n4701 = n4465 & ~n4700 ;
  assign n4702 = n3848 & ~n4700 ;
  assign n4703 = ( n4597 & n4701 ) | ( n4597 & n4702 ) | ( n4701 & n4702 );
  assign n4704 = n4465 | n4700 ;
  assign n4705 = n3848 | n4700 ;
  assign n4706 = ( n4597 & n4704 ) | ( n4597 & n4705 ) | ( n4704 & n4705 );
  assign n4707 = ( ~n4598 & n4703 ) | ( ~n4598 & n4706 ) | ( n4703 & n4706 );
  assign n4708 = n882 | n2173 ;
  assign n4709 = n4475 | n4708 ;
  assign n4710 = n144 | n4709 ;
  assign n4711 = n4606 | n4710 ;
  assign n4712 = n224 | n4711 ;
  assign n4713 = n262 | n4712 ;
  assign n4714 = n199 | n4713 ;
  assign n4715 = n213 | n4714 ;
  assign n4716 = n1043 | n4715 ;
  assign n4717 = n346 | n4716 ;
  assign n4718 = n312 | n4717 ;
  assign n4719 = n2685 & ~n3886 ;
  assign n4720 = n2540 & n2693 ;
  assign n4721 = n2690 & ~n3725 ;
  assign n4722 = n4720 | n4721 ;
  assign n4723 = n4719 | n4722 ;
  assign n4724 = n2697 & n3897 ;
  assign n4725 = n4723 | n4724 ;
  assign n4726 = n969 | n4725 ;
  assign n4727 = n969 & n4725 ;
  assign n4728 = n4726 & ~n4727 ;
  assign n4729 = n4639 & n4728 ;
  assign n4730 = n4518 & n4728 ;
  assign n4731 = n4508 & n4728 ;
  assign n4732 = ( n4498 & n4730 ) | ( n4498 & n4731 ) | ( n4730 & n4731 );
  assign n4733 = ( n4672 & n4729 ) | ( n4672 & n4732 ) | ( n4729 & n4732 );
  assign n4734 = n4639 | n4728 ;
  assign n4735 = n4518 | n4728 ;
  assign n4736 = n4508 | n4728 ;
  assign n4737 = ( n4498 & n4735 ) | ( n4498 & n4736 ) | ( n4735 & n4736 );
  assign n4738 = ( n4672 & n4734 ) | ( n4672 & n4737 ) | ( n4734 & n4737 );
  assign n4739 = ~n4733 & n4738 ;
  assign n4740 = n516 & n2580 ;
  assign n4741 = n32 | n1238 ;
  assign n4742 = n32 & n1238 ;
  assign n4743 = n4741 & ~n4742 ;
  assign n4744 = n4740 & n4743 ;
  assign n4745 = n4740 | n4743 ;
  assign n4746 = ~n4744 & n4745 ;
  assign n4747 = n4651 | n4656 ;
  assign n4748 = n2567 & n2848 ;
  assign n4749 = n2574 & n2918 ;
  assign n4750 = ~n2570 & n2846 ;
  assign n4751 = n4749 | n4750 ;
  assign n4752 = n4748 | n4751 ;
  assign n4753 = n2851 & ~n3027 ;
  assign n4754 = n4752 | n4753 ;
  assign n4755 = n516 & n4754 ;
  assign n4756 = n4754 & ~n4755 ;
  assign n4757 = n516 & ~n4755 ;
  assign n4758 = n4756 | n4757 ;
  assign n4759 = ( n4746 & n4747 ) | ( n4746 & n4758 ) | ( n4747 & n4758 );
  assign n4760 = ( ~n4746 & n4747 ) | ( ~n4746 & n4758 ) | ( n4747 & n4758 );
  assign n4761 = ( n4746 & ~n4759 ) | ( n4746 & n4760 ) | ( ~n4759 & n4760 );
  assign n4762 = n2555 & n2720 ;
  assign n4763 = n2655 & n2818 ;
  assign n4764 = ~n2550 & n2715 ;
  assign n4765 = n4763 | n4764 ;
  assign n4766 = n4762 | n4765 ;
  assign n4767 = n2726 & ~n3248 ;
  assign n4768 = n4766 | n4767 ;
  assign n4769 = n761 | n4768 ;
  assign n4770 = n761 & n4768 ;
  assign n4771 = n4769 & ~n4770 ;
  assign n4772 = ( n4671 & n4761 ) | ( n4671 & n4771 ) | ( n4761 & n4771 );
  assign n4773 = ( n4761 & n4771 ) | ( n4761 & ~n4772 ) | ( n4771 & ~n4772 );
  assign n4774 = ( n4671 & ~n4772 ) | ( n4671 & n4773 ) | ( ~n4772 & n4773 );
  assign n4775 = n4625 | n4629 ;
  assign n4776 = ( n4625 & n4675 ) | ( n4625 & n4775 ) | ( n4675 & n4775 );
  assign n4777 = ( n4739 & n4774 ) | ( n4739 & n4776 ) | ( n4774 & n4776 );
  assign n4778 = ( n4774 & n4776 ) | ( n4774 & ~n4777 ) | ( n4776 & ~n4777 );
  assign n4779 = ( n4739 & ~n4777 ) | ( n4739 & n4778 ) | ( ~n4777 & n4778 );
  assign n4780 = n4679 | n4685 ;
  assign n4781 = n4779 | n4780 ;
  assign n4782 = ( n4679 & n4685 ) | ( n4679 & n4779 ) | ( n4685 & n4779 );
  assign n4783 = n4781 & ~n4782 ;
  assign n4784 = n4718 & n4783 ;
  assign n4785 = n4718 | n4783 ;
  assign n4786 = ~n4784 & n4785 ;
  assign n4787 = n4689 | n4692 ;
  assign n4788 = n4786 & n4787 ;
  assign n4789 = n4786 | n4787 ;
  assign n4790 = ~n4788 & n4789 ;
  assign n4791 = n4697 & n4790 ;
  assign n4792 = n4697 | n4790 ;
  assign n4793 = ~n4791 & n4792 ;
  assign n4794 = n4469 | n4700 ;
  assign n4795 = n4597 | n4794 ;
  assign n4796 = n3848 & n4795 ;
  assign n4797 = ~n4793 & n4796 ;
  assign n4798 = n4793 & ~n4796 ;
  assign n4799 = n4797 | n4798 ;
  assign n4800 = n200 | n206 ;
  assign n4801 = n289 | n4800 ;
  assign n4802 = n236 | n4801 ;
  assign n4803 = n322 | n4802 ;
  assign n4804 = n394 | n4803 ;
  assign n4805 = n344 | n4804 ;
  assign n4806 = n401 | n2109 ;
  assign n4807 = n470 | n4806 ;
  assign n4808 = n286 | n4807 ;
  assign n4809 = n469 | n4808 ;
  assign n4810 = n190 | n4809 ;
  assign n4811 = n277 | n4810 ;
  assign n4812 = n191 | n4811 ;
  assign n4813 = n134 | n4812 ;
  assign n4814 = n124 | n4813 ;
  assign n4815 = n430 | n4814 ;
  assign n4816 = n924 | n2253 ;
  assign n4817 = n918 | n4816 ;
  assign n4818 = ( ~n3647 & n4815 ) | ( ~n3647 & n4817 ) | ( n4815 & n4817 );
  assign n4819 = n3647 | n4818 ;
  assign n4820 = n4805 | n4819 ;
  assign n4821 = n2693 & ~n3725 ;
  assign n4822 = n2690 & ~n3886 ;
  assign n4823 = n4821 | n4822 ;
  assign n4824 = ( n2697 & n4144 ) | ( n2697 & n4823 ) | ( n4144 & n4823 );
  assign n4825 = ( n969 & n4823 ) | ( n969 & ~n4824 ) | ( n4823 & ~n4824 );
  assign n4826 = n4824 | n4825 ;
  assign n4827 = ~n4823 & n4825 ;
  assign n4828 = ( ~n969 & n4826 ) | ( ~n969 & n4827 ) | ( n4826 & n4827 );
  assign n4829 = n2655 & n2848 ;
  assign n4830 = ~n2570 & n2918 ;
  assign n4831 = n2567 & n2846 ;
  assign n4832 = n4830 | n4831 ;
  assign n4833 = n4829 | n4832 ;
  assign n4834 = n2851 & n3494 ;
  assign n4835 = n4833 | n4834 ;
  assign n4836 = n516 | n4835 ;
  assign n4837 = n516 & n4835 ;
  assign n4838 = n4836 & ~n4837 ;
  assign n4839 = n516 & n2574 ;
  assign n4840 = ~n4740 & n4741 ;
  assign n4841 = ( n4741 & ~n4743 ) | ( n4741 & n4840 ) | ( ~n4743 & n4840 );
  assign n4842 = ( ~n4838 & n4839 ) | ( ~n4838 & n4841 ) | ( n4839 & n4841 );
  assign n4843 = ( n4839 & n4841 ) | ( n4839 & ~n4842 ) | ( n4841 & ~n4842 );
  assign n4844 = ( n4838 & n4842 ) | ( n4838 & ~n4843 ) | ( n4842 & ~n4843 );
  assign n4845 = n2540 & n2720 ;
  assign n4846 = ~n2550 & n2818 ;
  assign n4847 = n2555 & n2715 ;
  assign n4848 = n4846 | n4847 ;
  assign n4849 = n4845 | n4848 ;
  assign n4850 = n2672 & n2726 ;
  assign n4851 = n4849 | n4850 ;
  assign n4852 = n761 & n4851 ;
  assign n4853 = n761 | n4851 ;
  assign n4854 = ~n4852 & n4853 ;
  assign n4855 = ( n4759 & n4844 ) | ( n4759 & n4854 ) | ( n4844 & n4854 );
  assign n4856 = ( n4759 & ~n4844 ) | ( n4759 & n4854 ) | ( ~n4844 & n4854 );
  assign n4857 = ( n4844 & ~n4855 ) | ( n4844 & n4856 ) | ( ~n4855 & n4856 );
  assign n4858 = ( n4772 & ~n4828 ) | ( n4772 & n4857 ) | ( ~n4828 & n4857 );
  assign n4859 = ( n4828 & ~n4857 ) | ( n4828 & n4858 ) | ( ~n4857 & n4858 );
  assign n4860 = n4733 | n4738 ;
  assign n4861 = ( n4733 & ~n4772 ) | ( n4733 & n4860 ) | ( ~n4772 & n4860 );
  assign n4862 = ( n4671 & n4733 ) | ( n4671 & n4860 ) | ( n4733 & n4860 );
  assign n4863 = ( n4773 & n4861 ) | ( n4773 & n4862 ) | ( n4861 & n4862 );
  assign n4864 = n4858 & n4863 ;
  assign n4865 = ~n4772 & n4863 ;
  assign n4866 = ( n4859 & n4864 ) | ( n4859 & n4865 ) | ( n4864 & n4865 );
  assign n4867 = n4858 | n4863 ;
  assign n4868 = n4772 & ~n4863 ;
  assign n4869 = ( n4859 & n4867 ) | ( n4859 & ~n4868 ) | ( n4867 & ~n4868 );
  assign n4870 = ~n4866 & n4869 ;
  assign n4871 = n4739 & ~n4772 ;
  assign n4872 = n4671 & n4739 ;
  assign n4873 = ( n4773 & n4871 ) | ( n4773 & n4872 ) | ( n4871 & n4872 );
  assign n4874 = ( n4777 & n4782 ) | ( n4777 & ~n4873 ) | ( n4782 & ~n4873 );
  assign n4875 = n4870 | n4874 ;
  assign n4876 = n4777 & n4870 ;
  assign n4877 = n4870 & ~n4873 ;
  assign n4878 = ( n4782 & n4876 ) | ( n4782 & n4877 ) | ( n4876 & n4877 );
  assign n4879 = n4875 & ~n4878 ;
  assign n4880 = n4820 | n4879 ;
  assign n4881 = n4820 & n4879 ;
  assign n4882 = n4880 & ~n4881 ;
  assign n4883 = n4784 | n4787 ;
  assign n4884 = ( n4784 & n4786 ) | ( n4784 & n4883 ) | ( n4786 & n4883 );
  assign n4885 = n4882 & n4884 ;
  assign n4886 = n4882 | n4884 ;
  assign n4887 = ~n4885 & n4886 ;
  assign n4888 = n4791 | n4887 ;
  assign n4889 = n4791 & n4887 ;
  assign n4890 = n4888 & ~n4889 ;
  assign n4891 = n4793 | n4795 ;
  assign n4892 = n3848 & n4891 ;
  assign n4893 = ~n4890 & n4892 ;
  assign n4894 = n4890 & ~n4892 ;
  assign n4895 = n4893 | n4894 ;
  assign n4907 = n4866 | n4878 ;
  assign n4908 = n4759 & ~n4844 ;
  assign n4909 = ( n4844 & n4854 ) | ( n4844 & n4908 ) | ( n4854 & n4908 );
  assign n4910 = n2693 & ~n3886 ;
  assign n4911 = n2697 & ~n4142 ;
  assign n4912 = n4910 | n4911 ;
  assign n4913 = n969 & ~n4912 ;
  assign n4914 = ~n969 & n4912 ;
  assign n4915 = n4913 | n4914 ;
  assign n4916 = n4758 & n4915 ;
  assign n4917 = n4747 & n4915 ;
  assign n4918 = ( n4746 & n4916 ) | ( n4746 & n4917 ) | ( n4916 & n4917 );
  assign n4919 = n4844 & n4918 ;
  assign n4920 = ( n4908 & n4915 ) | ( n4908 & n4919 ) | ( n4915 & n4919 );
  assign n4921 = ~n4758 & n4915 ;
  assign n4922 = ~n4747 & n4915 ;
  assign n4923 = ( ~n4746 & n4921 ) | ( ~n4746 & n4922 ) | ( n4921 & n4922 );
  assign n4924 = ( n4844 & n4915 ) | ( n4844 & n4923 ) | ( n4915 & n4923 );
  assign n4925 = ( n4909 & n4920 ) | ( n4909 & n4924 ) | ( n4920 & n4924 );
  assign n4926 = n4854 | n4915 ;
  assign n4927 = n4758 | n4915 ;
  assign n4928 = n4747 | n4915 ;
  assign n4929 = ( n4746 & n4927 ) | ( n4746 & n4928 ) | ( n4927 & n4928 );
  assign n4930 = ( n4844 & n4926 ) | ( n4844 & n4929 ) | ( n4926 & n4929 );
  assign n4931 = ~n4925 & n4930 ;
  assign n4932 = n516 & ~n2577 ;
  assign n4933 = ~n2550 & n2848 ;
  assign n4934 = n2567 & n2918 ;
  assign n4935 = n2655 & n2846 ;
  assign n4936 = n4934 | n4935 ;
  assign n4937 = n4933 | n4936 ;
  assign n4938 = n2851 & ~n3264 ;
  assign n4939 = n4937 | n4938 ;
  assign n4940 = n516 & n4939 ;
  assign n4941 = n4939 & ~n4940 ;
  assign n4942 = n516 & ~n4940 ;
  assign n4943 = n4941 | n4942 ;
  assign n4944 = n4932 | n4943 ;
  assign n4945 = n4932 & n4943 ;
  assign n4946 = n4944 & ~n4945 ;
  assign n4947 = n2720 & ~n3725 ;
  assign n4948 = n2555 & n2818 ;
  assign n4949 = n2540 & n2715 ;
  assign n4950 = n4948 | n4949 ;
  assign n4951 = n4947 | n4950 ;
  assign n4952 = n2726 & ~n3741 ;
  assign n4953 = n4951 | n4952 ;
  assign n4954 = n761 | n4953 ;
  assign n4955 = n761 & n4953 ;
  assign n4956 = n4954 & ~n4955 ;
  assign n4957 = ( n4842 & n4946 ) | ( n4842 & ~n4956 ) | ( n4946 & ~n4956 );
  assign n4958 = ( ~n4842 & n4946 ) | ( ~n4842 & n4956 ) | ( n4946 & n4956 );
  assign n4959 = ( ~n4946 & n4957 ) | ( ~n4946 & n4958 ) | ( n4957 & n4958 );
  assign n4960 = n4930 & ~n4959 ;
  assign n4961 = ~n4925 & n4960 ;
  assign n4962 = n4930 | n4959 ;
  assign n4963 = ( ~n4925 & n4959 ) | ( ~n4925 & n4962 ) | ( n4959 & n4962 );
  assign n4964 = ( ~n4931 & n4961 ) | ( ~n4931 & n4963 ) | ( n4961 & n4963 );
  assign n4965 = ( n4772 & n4828 ) | ( n4772 & n4857 ) | ( n4828 & n4857 );
  assign n4966 = ( ~n4866 & n4964 ) | ( ~n4866 & n4965 ) | ( n4964 & n4965 );
  assign n4967 = n4964 & n4965 ;
  assign n4968 = ( ~n4878 & n4966 ) | ( ~n4878 & n4967 ) | ( n4966 & n4967 );
  assign n4969 = ( n4964 & n4965 ) | ( n4964 & ~n4967 ) | ( n4965 & ~n4967 );
  assign n4970 = ( n4964 & n4965 ) | ( n4964 & ~n4966 ) | ( n4965 & ~n4966 );
  assign n4971 = ( n4878 & n4969 ) | ( n4878 & n4970 ) | ( n4969 & n4970 );
  assign n4972 = ( n4907 & n4968 ) | ( n4907 & ~n4971 ) | ( n4968 & ~n4971 );
  assign n4896 = n144 | n682 ;
  assign n4897 = n3589 | n4896 ;
  assign n4898 = n2486 | n4897 ;
  assign n4899 = n2354 | n4898 ;
  assign n4900 = n2523 | n4899 ;
  assign n4901 = n293 | n4900 ;
  assign n4902 = n290 | n4901 ;
  assign n4903 = n191 | n4902 ;
  assign n4904 = n271 | n4903 ;
  assign n4905 = n494 | n4904 ;
  assign n4906 = n154 | n4905 ;
  assign n4973 = n4906 & n4972 ;
  assign n4974 = ( n397 & n4972 ) | ( n397 & n4973 ) | ( n4972 & n4973 );
  assign n4975 = n4906 | n4972 ;
  assign n4976 = n397 | n4975 ;
  assign n4977 = ~n4974 & n4976 ;
  assign n4978 = n4881 | n4882 ;
  assign n4979 = ( n4881 & n4884 ) | ( n4881 & n4978 ) | ( n4884 & n4978 );
  assign n4980 = n4977 & n4979 ;
  assign n4981 = n4977 | n4979 ;
  assign n4982 = ~n4980 & n4981 ;
  assign n4983 = n4889 | n4982 ;
  assign n4984 = n4889 & n4982 ;
  assign n4985 = n4983 & ~n4984 ;
  assign n4986 = n4890 | n4891 ;
  assign n4987 = n3848 & n4986 ;
  assign n4988 = ~n4985 & n4987 ;
  assign n4989 = n4985 & ~n4987 ;
  assign n4990 = n4988 | n4989 ;
  assign n5001 = n516 & ~n2570 ;
  assign n5002 = ~n4839 & n5001 ;
  assign n5003 = n4932 & ~n5002 ;
  assign n5004 = ( n4943 & n5002 ) | ( n4943 & ~n5003 ) | ( n5002 & ~n5003 );
  assign n5005 = n516 & n2567 ;
  assign n5006 = ( ~n969 & n4839 ) | ( ~n969 & n5005 ) | ( n4839 & n5005 );
  assign n5007 = ( n969 & ~n5005 ) | ( n969 & n5006 ) | ( ~n5005 & n5006 );
  assign n5008 = ( ~n4839 & n5006 ) | ( ~n4839 & n5007 ) | ( n5006 & n5007 );
  assign n5009 = n5004 & ~n5008 ;
  assign n5010 = ~n5004 & n5008 ;
  assign n5011 = n5009 | n5010 ;
  assign n5012 = n2555 & n2848 ;
  assign n5013 = n2655 & n2918 ;
  assign n5014 = ~n2550 & n2846 ;
  assign n5015 = n5013 | n5014 ;
  assign n5016 = n5012 | n5015 ;
  assign n5017 = n2851 & ~n3248 ;
  assign n5018 = n5016 | n5017 ;
  assign n5019 = n516 & n5018 ;
  assign n5020 = n516 & ~n5019 ;
  assign n5021 = n5018 & ~n5019 ;
  assign n5022 = n5020 | n5021 ;
  assign n5023 = ~n5011 & n5022 ;
  assign n5024 = n5011 & n5022 ;
  assign n5025 = ( n5011 & n5023 ) | ( n5011 & ~n5024 ) | ( n5023 & ~n5024 );
  assign n5026 = n2720 & ~n3886 ;
  assign n5027 = n2540 & n2818 ;
  assign n5028 = n2715 & ~n3725 ;
  assign n5029 = n5027 | n5028 ;
  assign n5030 = n5026 | n5029 ;
  assign n5031 = n2726 & n3897 ;
  assign n5032 = n5030 | n5031 ;
  assign n5033 = n761 | n5032 ;
  assign n5034 = n761 & n5032 ;
  assign n5035 = n5033 & ~n5034 ;
  assign n5036 = n4956 & n5035 ;
  assign n5037 = n4838 & n5035 ;
  assign n5038 = ~n4839 & n5035 ;
  assign n5039 = ( ~n4841 & n5037 ) | ( ~n4841 & n5038 ) | ( n5037 & n5038 );
  assign n5040 = ( ~n4946 & n5036 ) | ( ~n4946 & n5039 ) | ( n5036 & n5039 );
  assign n5041 = n4957 | n5040 ;
  assign n5042 = ~n4956 & n5035 ;
  assign n5043 = ~n4838 & n5035 ;
  assign n5044 = n4839 & n5035 ;
  assign n5045 = ( n4841 & n5043 ) | ( n4841 & n5044 ) | ( n5043 & n5044 );
  assign n5046 = ( n4946 & n5042 ) | ( n4946 & n5045 ) | ( n5042 & n5045 );
  assign n5047 = n5041 & ~n5046 ;
  assign n5048 = n5025 & n5047 ;
  assign n5049 = n5025 | n5047 ;
  assign n5050 = ~n5048 & n5049 ;
  assign n5051 = n4925 | n5050 ;
  assign n5052 = n4930 & n4959 ;
  assign n5053 = ~n4925 & n5052 ;
  assign n5054 = n5051 | n5053 ;
  assign n5055 = ( n4925 & n5050 ) | ( n4925 & n5053 ) | ( n5050 & n5053 );
  assign n5056 = n5054 & ~n5055 ;
  assign n5057 = n4964 | n4965 ;
  assign n5058 = ( n4866 & n4964 ) | ( n4866 & n4965 ) | ( n4964 & n4965 );
  assign n5059 = ( n4878 & n5057 ) | ( n4878 & n5058 ) | ( n5057 & n5058 );
  assign n5060 = n5056 | n5059 ;
  assign n5061 = n5056 & n5058 ;
  assign n5062 = n5056 & n5057 ;
  assign n5063 = ( n4878 & n5061 ) | ( n4878 & n5062 ) | ( n5061 & n5062 );
  assign n5064 = n5060 & ~n5063 ;
  assign n4991 = n368 | n2022 ;
  assign n4992 = n160 | n398 ;
  assign n4993 = n4991 | n4992 ;
  assign n4994 = n2480 | n3634 ;
  assign n4995 = n1057 | n4994 ;
  assign n4996 = n2523 | n4995 ;
  assign n4997 = n4993 | n4996 ;
  assign n4998 = n268 | n922 ;
  assign n4999 = n278 | n4998 ;
  assign n5000 = n4997 | n4999 ;
  assign n5065 = n5000 & n5064 ;
  assign n5066 = ( n553 & n5064 ) | ( n553 & n5065 ) | ( n5064 & n5065 );
  assign n5067 = n5000 | n5064 ;
  assign n5068 = n553 | n5067 ;
  assign n5069 = ~n5066 & n5068 ;
  assign n5070 = n4973 | n4979 ;
  assign n5071 = n4972 | n4979 ;
  assign n5072 = ( n397 & n5070 ) | ( n397 & n5071 ) | ( n5070 & n5071 );
  assign n5073 = ( n4974 & n4977 ) | ( n4974 & n5072 ) | ( n4977 & n5072 );
  assign n5074 = n5069 & n5073 ;
  assign n5075 = n5069 | n5073 ;
  assign n5076 = ~n5074 & n5075 ;
  assign n5077 = n4984 | n5076 ;
  assign n5078 = n4984 & n5076 ;
  assign n5079 = n5077 & ~n5078 ;
  assign n5080 = n4985 | n4986 ;
  assign n5081 = n3848 & n5080 ;
  assign n5082 = ~n5079 & n5081 ;
  assign n5083 = n5079 & ~n5081 ;
  assign n5084 = n5082 | n5083 ;
  assign n5085 = n198 | n320 ;
  assign n5086 = n555 | n949 ;
  assign n5087 = n860 | n5086 ;
  assign n5088 = n3708 | n5087 ;
  assign n5089 = ( ~n432 & n3707 ) | ( ~n432 & n5088 ) | ( n3707 & n5088 );
  assign n5090 = n3707 & n5088 ;
  assign n5091 = ( ~n428 & n5089 ) | ( ~n428 & n5090 ) | ( n5089 & n5090 );
  assign n5092 = n433 | n5091 ;
  assign n5093 = n5085 | n5092 ;
  assign n5094 = n2540 & n2848 ;
  assign n5095 = ~n2550 & n2918 ;
  assign n5096 = n2555 & n2846 ;
  assign n5097 = n5095 | n5096 ;
  assign n5098 = n5094 | n5097 ;
  assign n5099 = n2672 & n2851 ;
  assign n5100 = n5098 | n5099 ;
  assign n5101 = n516 | n5100 ;
  assign n5102 = n516 & n5100 ;
  assign n5103 = n5101 & ~n5102 ;
  assign n5104 = n516 & n2655 ;
  assign n5105 = ( ~n5006 & n5103 ) | ( ~n5006 & n5104 ) | ( n5103 & n5104 );
  assign n5106 = ( n5006 & ~n5104 ) | ( n5006 & n5105 ) | ( ~n5104 & n5105 );
  assign n5107 = ( ~n5103 & n5105 ) | ( ~n5103 & n5106 ) | ( n5105 & n5106 );
  assign n5108 = n5009 | n5022 ;
  assign n5109 = ( n5009 & ~n5011 ) | ( n5009 & n5108 ) | ( ~n5011 & n5108 );
  assign n5110 = ~n5107 & n5109 ;
  assign n5111 = n2726 & n4144 ;
  assign n5112 = n2818 & ~n3725 ;
  assign n5113 = n2715 & ~n3886 ;
  assign n5114 = n5112 | n5113 ;
  assign n5115 = n5111 | n5114 ;
  assign n5116 = n761 & n5115 ;
  assign n5117 = n761 | n5115 ;
  assign n5118 = ~n5116 & n5117 ;
  assign n5119 = ( ~n5107 & n5109 ) | ( ~n5107 & n5118 ) | ( n5109 & n5118 );
  assign n5120 = ~n5110 & n5119 ;
  assign n5121 = n5105 & ~n5118 ;
  assign n5122 = n5103 | n5118 ;
  assign n5123 = ( n5106 & n5121 ) | ( n5106 & ~n5122 ) | ( n5121 & ~n5122 );
  assign n5124 = ( n5109 & ~n5118 ) | ( n5109 & n5123 ) | ( ~n5118 & n5123 );
  assign n5125 = ( ~n5109 & n5110 ) | ( ~n5109 & n5124 ) | ( n5110 & n5124 );
  assign n5126 = n5120 | n5125 ;
  assign n5127 = ~n5040 & n5049 ;
  assign n5128 = n5055 | n5058 ;
  assign n5129 = ( n5055 & n5056 ) | ( n5055 & n5128 ) | ( n5056 & n5128 );
  assign n5130 = ( n5126 & n5127 ) | ( n5126 & ~n5129 ) | ( n5127 & ~n5129 );
  assign n5131 = n5055 | n5057 ;
  assign n5132 = ( n5055 & n5056 ) | ( n5055 & n5131 ) | ( n5056 & n5131 );
  assign n5133 = ( n5126 & n5127 ) | ( n5126 & ~n5132 ) | ( n5127 & ~n5132 );
  assign n5134 = ( ~n4878 & n5130 ) | ( ~n4878 & n5133 ) | ( n5130 & n5133 );
  assign n5135 = ( n4878 & n5129 ) | ( n4878 & n5132 ) | ( n5129 & n5132 );
  assign n5136 = ( ~n5127 & n5134 ) | ( ~n5127 & n5135 ) | ( n5134 & n5135 );
  assign n5137 = ( ~n5126 & n5134 ) | ( ~n5126 & n5136 ) | ( n5134 & n5136 );
  assign n5138 = n5093 | n5137 ;
  assign n5139 = n5093 & n5137 ;
  assign n5140 = n5138 & ~n5139 ;
  assign n5141 = n5066 | n5069 ;
  assign n5142 = ( n5066 & n5073 ) | ( n5066 & n5141 ) | ( n5073 & n5141 );
  assign n5143 = n5140 & n5142 ;
  assign n5144 = n5140 | n5142 ;
  assign n5145 = ~n5143 & n5144 ;
  assign n5146 = n5078 | n5145 ;
  assign n5147 = n5078 & n5145 ;
  assign n5148 = n5146 & ~n5147 ;
  assign n5149 = n5079 | n5080 ;
  assign n5150 = n3848 & n5149 ;
  assign n5151 = ~n5148 & n5150 ;
  assign n5152 = n5148 & ~n5150 ;
  assign n5153 = n5151 | n5152 ;
  assign n5154 = n150 | n184 ;
  assign n5155 = n289 | n5154 ;
  assign n5156 = n494 | n5155 ;
  assign n5157 = n549 | n5156 ;
  assign n5158 = n2273 | n5157 ;
  assign n5159 = n900 | n5158 ;
  assign n5160 = n4032 | n5159 ;
  assign n5161 = n2446 | n5160 ;
  assign n5162 = n283 | n5161 ;
  assign n5163 = n177 | n5162 ;
  assign n5164 = n430 | n5163 ;
  assign n5165 = n2033 | n5164 ;
  assign n5166 = n516 & ~n2550 ;
  assign n5167 = ~n5104 & n5166 ;
  assign n5168 = n5104 & ~n5166 ;
  assign n5169 = n5167 | n5168 ;
  assign n5170 = ( n5006 & n5103 ) | ( n5006 & ~n5104 ) | ( n5103 & ~n5104 );
  assign n5171 = n5169 | n5170 ;
  assign n5172 = n5169 & n5170 ;
  assign n5173 = n5171 & ~n5172 ;
  assign n5174 = n2818 & ~n3886 ;
  assign n5175 = n2726 & ~n4142 ;
  assign n5176 = n5174 | n5175 ;
  assign n5177 = n761 | n5176 ;
  assign n5178 = n761 & n5176 ;
  assign n5179 = n5177 & ~n5178 ;
  assign n5180 = n2848 & ~n3725 ;
  assign n5181 = n2555 & n2918 ;
  assign n5182 = n2540 & n2846 ;
  assign n5183 = n5181 | n5182 ;
  assign n5184 = n5180 | n5183 ;
  assign n5185 = n2851 & ~n3741 ;
  assign n5186 = n5184 | n5185 ;
  assign n5187 = n516 & n5186 ;
  assign n5188 = n516 & ~n5187 ;
  assign n5189 = n5186 & ~n5187 ;
  assign n5190 = n5188 | n5189 ;
  assign n5191 = n5179 & n5190 ;
  assign n5192 = n5190 & ~n5191 ;
  assign n5193 = ( n5179 & ~n5191 ) | ( n5179 & n5192 ) | ( ~n5191 & n5192 );
  assign n5194 = n5173 & ~n5193 ;
  assign n5195 = n5193 | n5194 ;
  assign n5196 = ( ~n5173 & n5194 ) | ( ~n5173 & n5195 ) | ( n5194 & n5195 );
  assign n5197 = ~n5110 & n5196 ;
  assign n5198 = ~n5120 & n5197 ;
  assign n5199 = n5119 & ~n5196 ;
  assign n5200 = n5198 | n5199 ;
  assign n5201 = n5134 & n5200 ;
  assign n5202 = n5126 | n5127 ;
  assign n5203 = n5126 & n5127 ;
  assign n5204 = n5202 & ~n5203 ;
  assign n5205 = n5055 & n5204 ;
  assign n5206 = n5200 | n5202 ;
  assign n5207 = ( n5200 & ~n5205 ) | ( n5200 & n5206 ) | ( ~n5205 & n5206 );
  assign n5208 = ( n5200 & ~n5204 ) | ( n5200 & n5206 ) | ( ~n5204 & n5206 );
  assign n5209 = ( ~n5061 & n5207 ) | ( ~n5061 & n5208 ) | ( n5207 & n5208 );
  assign n5210 = ( ~n5062 & n5207 ) | ( ~n5062 & n5208 ) | ( n5207 & n5208 );
  assign n5211 = ( ~n4878 & n5209 ) | ( ~n4878 & n5210 ) | ( n5209 & n5210 );
  assign n5212 = ~n5201 & n5211 ;
  assign n5213 = ( n5139 & n5165 ) | ( n5139 & n5212 ) | ( n5165 & n5212 );
  assign n5214 = ( n5138 & n5165 ) | ( n5138 & n5212 ) | ( n5165 & n5212 );
  assign n5215 = ( n5142 & n5213 ) | ( n5142 & n5214 ) | ( n5213 & n5214 );
  assign n5216 = ( ~n5139 & n5165 ) | ( ~n5139 & n5212 ) | ( n5165 & n5212 );
  assign n5217 = ( ~n5138 & n5165 ) | ( ~n5138 & n5212 ) | ( n5165 & n5212 );
  assign n5218 = ( ~n5142 & n5216 ) | ( ~n5142 & n5217 ) | ( n5216 & n5217 );
  assign n5219 = n5139 | n5140 ;
  assign n5220 = ( n5139 & n5142 ) | ( n5139 & n5219 ) | ( n5142 & n5219 );
  assign n5221 = ( ~n5215 & n5218 ) | ( ~n5215 & n5220 ) | ( n5218 & n5220 );
  assign n5222 = n5147 | n5221 ;
  assign n5223 = n5147 & n5221 ;
  assign n5224 = n5222 & ~n5223 ;
  assign n5225 = n5148 | n5149 ;
  assign n5226 = n3848 & n5225 ;
  assign n5227 = ~n5224 & n5226 ;
  assign n5228 = n5224 & ~n5226 ;
  assign n5229 = n5227 | n5228 ;
  assign n5230 = n260 | n262 ;
  assign n5231 = n214 | n334 ;
  assign n5232 = n5230 | n5231 ;
  assign n5233 = n451 | n460 ;
  assign n5234 = n3855 | n5233 ;
  assign n5235 = n5232 | n5234 ;
  assign n5236 = n1042 | n2102 ;
  assign n5237 = n2191 | n5236 ;
  assign n5238 = n5235 | n5237 ;
  assign n5239 = n304 | n5238 ;
  assign n5240 = n3670 | n5239 ;
  assign n5241 = n200 | n323 ;
  assign n5242 = n418 | n5241 ;
  assign n5243 = n321 | n5242 ;
  assign n5244 = n347 | n5243 ;
  assign n5245 = n414 | n5244 ;
  assign n5246 = n5240 | n5245 ;
  assign n5247 = n2848 & ~n3886 ;
  assign n5248 = n2540 & n2918 ;
  assign n5249 = n2846 & ~n3725 ;
  assign n5250 = n5248 | n5249 ;
  assign n5251 = n5247 | n5250 ;
  assign n5252 = n2851 & n3897 ;
  assign n5253 = n5251 | n5252 ;
  assign n5254 = n516 & n5253 ;
  assign n5255 = n5253 & ~n5254 ;
  assign n5256 = n516 & ~n5254 ;
  assign n5257 = n5255 | n5256 ;
  assign n5258 = ~n5168 & n5169 ;
  assign n5259 = n516 & n2555 ;
  assign n5260 = ~n761 & n5166 ;
  assign n5261 = n761 & ~n5166 ;
  assign n5262 = n5260 | n5261 ;
  assign n5263 = n5259 & ~n5262 ;
  assign n5264 = ~n5259 & n5262 ;
  assign n5265 = n5263 | n5264 ;
  assign n5266 = ( n5170 & n5257 ) | ( n5170 & ~n5265 ) | ( n5257 & ~n5265 );
  assign n5267 = ( n5168 & n5257 ) | ( n5168 & ~n5265 ) | ( n5257 & ~n5265 );
  assign n5268 = ( ~n5258 & n5266 ) | ( ~n5258 & n5267 ) | ( n5266 & n5267 );
  assign n5269 = ( n5168 & n5170 ) | ( n5168 & ~n5258 ) | ( n5170 & ~n5258 );
  assign n5270 = ( n5265 & n5268 ) | ( n5265 & ~n5269 ) | ( n5268 & ~n5269 );
  assign n5271 = ( ~n5257 & n5268 ) | ( ~n5257 & n5270 ) | ( n5268 & n5270 );
  assign n5272 = ~n5173 & n5193 ;
  assign n5273 = n5191 & ~n5268 ;
  assign n5274 = n5191 & n5257 ;
  assign n5275 = ( ~n5270 & n5273 ) | ( ~n5270 & n5274 ) | ( n5273 & n5274 );
  assign n5276 = ( ~n5271 & n5272 ) | ( ~n5271 & n5275 ) | ( n5272 & n5275 );
  assign n5277 = ~n5191 & n5268 ;
  assign n5278 = n5191 | n5257 ;
  assign n5279 = ( n5270 & n5277 ) | ( n5270 & ~n5278 ) | ( n5277 & ~n5278 );
  assign n5280 = ~n5272 & n5279 ;
  assign n5281 = n5276 | n5280 ;
  assign n5282 = n5199 & ~n5281 ;
  assign n5283 = ( n5211 & n5281 ) | ( n5211 & ~n5282 ) | ( n5281 & ~n5282 );
  assign n5284 = ~n5199 & n5281 ;
  assign n5285 = n5211 & n5284 ;
  assign n5286 = n5283 & ~n5285 ;
  assign n5287 = n5246 & n5286 ;
  assign n5288 = n5246 | n5286 ;
  assign n5289 = ~n5287 & n5288 ;
  assign n5290 = n5214 & ~n5289 ;
  assign n5291 = n5213 & ~n5289 ;
  assign n5292 = ( n5142 & n5290 ) | ( n5142 & n5291 ) | ( n5290 & n5291 );
  assign n5293 = ~n5214 & n5289 ;
  assign n5294 = ~n5213 & n5289 ;
  assign n5295 = ( ~n5142 & n5293 ) | ( ~n5142 & n5294 ) | ( n5293 & n5294 );
  assign n5296 = n5292 | n5295 ;
  assign n5297 = n5221 & n5296 ;
  assign n5298 = n5147 & n5297 ;
  assign n5299 = n5221 | n5296 ;
  assign n5300 = ( n5147 & n5296 ) | ( n5147 & n5299 ) | ( n5296 & n5299 );
  assign n5301 = ~n5298 & n5300 ;
  assign n5302 = n5224 | n5225 ;
  assign n5303 = n3848 & n5302 ;
  assign n5304 = ~n5301 & n5303 ;
  assign n5305 = n5301 & ~n5303 ;
  assign n5306 = n5304 | n5305 ;
  assign n5307 = n5287 | n5289 ;
  assign n5308 = n2273 | n2334 ;
  assign n5309 = n2127 | n5308 ;
  assign n5310 = n152 | n5309 ;
  assign n5311 = n1388 | n5310 ;
  assign n5312 = n932 | n5311 ;
  assign n5313 = n2115 | n5312 ;
  assign n5314 = n205 | n2523 ;
  assign n5315 = n225 | n5314 ;
  assign n5316 = n183 | n5315 ;
  assign n5317 = n5313 | n5316 ;
  assign n5318 = n323 | n5317 ;
  assign n5319 = n333 | n5318 ;
  assign n5320 = n198 | n5319 ;
  assign n5321 = n234 | n5320 ;
  assign n5322 = n516 & n2540 ;
  assign n5323 = n5259 | n5260 ;
  assign n5324 = ( n5260 & ~n5262 ) | ( n5260 & n5323 ) | ( ~n5262 & n5323 );
  assign n5325 = n2846 & ~n3886 ;
  assign n5326 = n2845 | n3725 ;
  assign n5327 = n2917 & ~n5326 ;
  assign n5328 = n5325 | n5327 ;
  assign n5329 = n2851 & n4144 ;
  assign n5330 = n516 & ~n5329 ;
  assign n5331 = ~n5328 & n5330 ;
  assign n5332 = n516 & ~n5331 ;
  assign n5333 = ( n5322 & n5324 ) | ( n5322 & n5331 ) | ( n5324 & n5331 );
  assign n5334 = n5328 | n5329 ;
  assign n5335 = ( n5322 & n5324 ) | ( n5322 & n5334 ) | ( n5324 & n5334 );
  assign n5336 = ( ~n5332 & n5333 ) | ( ~n5332 & n5335 ) | ( n5333 & n5335 );
  assign n5337 = ( n5322 & n5324 ) | ( n5322 & ~n5336 ) | ( n5324 & ~n5336 );
  assign n5338 = n5268 & n5336 ;
  assign n5339 = ( n5331 & ~n5332 ) | ( n5331 & n5334 ) | ( ~n5332 & n5334 );
  assign n5340 = n5268 & ~n5339 ;
  assign n5341 = ( ~n5337 & n5338 ) | ( ~n5337 & n5340 ) | ( n5338 & n5340 );
  assign n5342 = n5268 | n5336 ;
  assign n5343 = ~n5268 & n5339 ;
  assign n5344 = ( n5337 & ~n5342 ) | ( n5337 & n5343 ) | ( ~n5342 & n5343 );
  assign n5345 = n5341 | n5344 ;
  assign n5346 = n5276 | n5282 ;
  assign n5347 = ~n5276 & n5281 ;
  assign n5348 = ( n5211 & ~n5346 ) | ( n5211 & n5347 ) | ( ~n5346 & n5347 );
  assign n5349 = n5345 | n5348 ;
  assign n5350 = n5345 & n5348 ;
  assign n5351 = n5349 & ~n5350 ;
  assign n5352 = n5321 | n5351 ;
  assign n5353 = n5321 & n5351 ;
  assign n5354 = n5352 & ~n5353 ;
  assign n5355 = n5213 & n5354 ;
  assign n5356 = n5287 & n5354 ;
  assign n5357 = ( n5307 & n5355 ) | ( n5307 & n5356 ) | ( n5355 & n5356 );
  assign n5358 = ( n5287 & n5289 ) | ( n5287 & n5354 ) | ( n5289 & n5354 );
  assign n5359 = ( n5214 & n5356 ) | ( n5214 & n5358 ) | ( n5356 & n5358 );
  assign n5360 = ( n5142 & n5357 ) | ( n5142 & n5359 ) | ( n5357 & n5359 );
  assign n5361 = n5307 | n5354 ;
  assign n5362 = n5287 | n5354 ;
  assign n5363 = ( n5214 & n5361 ) | ( n5214 & n5362 ) | ( n5361 & n5362 );
  assign n5364 = n5213 | n5354 ;
  assign n5365 = ( n5307 & n5362 ) | ( n5307 & n5364 ) | ( n5362 & n5364 );
  assign n5366 = ( n5142 & n5363 ) | ( n5142 & n5365 ) | ( n5363 & n5365 );
  assign n5367 = ~n5360 & n5366 ;
  assign n5368 = n5296 & n5367 ;
  assign n5369 = n5223 & n5368 ;
  assign n5370 = n5298 | n5367 ;
  assign n5371 = ~n5369 & n5370 ;
  assign n5372 = n5301 | n5302 ;
  assign n5373 = n3848 & n5372 ;
  assign n5374 = ~n5371 & n5373 ;
  assign n5375 = n5371 & ~n5373 ;
  assign n5376 = n5374 | n5375 ;
  assign n5377 = n293 | n1109 ;
  assign n5378 = n305 | n5377 ;
  assign n5379 = n1108 | n5378 ;
  assign n5380 = n129 | n5379 ;
  assign n5381 = n947 | n5380 ;
  assign n5382 = n422 | n5157 ;
  assign n5383 = ( ~n2280 & n5381 ) | ( ~n2280 & n5382 ) | ( n5381 & n5382 );
  assign n5384 = n5381 & n5382 ;
  assign n5385 = ( ~n2276 & n5383 ) | ( ~n2276 & n5384 ) | ( n5383 & n5384 );
  assign n5386 = n2281 | n5385 ;
  assign n5387 = n158 | n272 ;
  assign n5388 = n154 | n234 ;
  assign n5389 = n5387 | n5388 ;
  assign n5390 = n240 | n5389 ;
  assign n5391 = n183 | n1020 ;
  assign n5392 = n1019 | n5391 ;
  assign n5393 = n5390 | n5392 ;
  assign n5394 = n5386 | n5393 ;
  assign n5395 = n516 & ~n3733 ;
  assign n5396 = n2851 & ~n4142 ;
  assign n5397 = n2845 | n3886 ;
  assign n5398 = n2917 & ~n5397 ;
  assign n5399 = n5396 | n5398 ;
  assign n5400 = n516 & ~n5399 ;
  assign n5401 = ~n516 & n5399 ;
  assign n5402 = n5400 | n5401 ;
  assign n5403 = ~n5395 & n5402 ;
  assign n5404 = n5395 & ~n5402 ;
  assign n5405 = n5403 | n5404 ;
  assign n5406 = ( ~n5322 & n5324 ) | ( ~n5322 & n5331 ) | ( n5324 & n5331 );
  assign n5407 = ( ~n5322 & n5324 ) | ( ~n5322 & n5334 ) | ( n5324 & n5334 );
  assign n5408 = ( ~n5332 & n5406 ) | ( ~n5332 & n5407 ) | ( n5406 & n5407 );
  assign n5409 = n5405 & ~n5408 ;
  assign n5410 = ~n5405 & n5408 ;
  assign n5411 = n5409 | n5410 ;
  assign n5412 = ~n5341 & n5348 ;
  assign n5413 = ( ~n5341 & n5345 ) | ( ~n5341 & n5412 ) | ( n5345 & n5412 );
  assign n5414 = n5411 & n5413 ;
  assign n5415 = n5411 | n5413 ;
  assign n5416 = ~n5414 & n5415 ;
  assign n5417 = n5394 & n5416 ;
  assign n5418 = n5394 | n5416 ;
  assign n5419 = ~n5417 & n5418 ;
  assign n5420 = n5353 & ~n5417 ;
  assign n5421 = ( n5357 & n5419 ) | ( n5357 & n5420 ) | ( n5419 & n5420 );
  assign n5422 = n5353 & n5419 ;
  assign n5423 = ( n5358 & n5419 ) | ( n5358 & n5422 ) | ( n5419 & n5422 );
  assign n5424 = ( n5356 & n5419 ) | ( n5356 & n5422 ) | ( n5419 & n5422 );
  assign n5425 = ( n5214 & n5423 ) | ( n5214 & n5424 ) | ( n5423 & n5424 );
  assign n5426 = ( n5142 & n5421 ) | ( n5142 & n5425 ) | ( n5421 & n5425 );
  assign n5427 = n5353 | n5419 ;
  assign n5428 = n5359 | n5427 ;
  assign n5429 = n5357 | n5427 ;
  assign n5430 = ( n5142 & n5428 ) | ( n5142 & n5429 ) | ( n5428 & n5429 );
  assign n5431 = ~n5426 & n5430 ;
  assign n5432 = n5368 & n5431 ;
  assign n5433 = n5223 & n5432 ;
  assign n5434 = n5368 | n5431 ;
  assign n5435 = ( n5223 & n5431 ) | ( n5223 & n5434 ) | ( n5431 & n5434 );
  assign n5436 = ~n5433 & n5435 ;
  assign n5437 = n5371 | n5372 ;
  assign n5438 = n3848 & n5437 ;
  assign n5439 = ~n5436 & n5438 ;
  assign n5440 = n5436 & ~n5438 ;
  assign n5441 = n5439 | n5440 ;
  assign n5442 = n451 | n5232 ;
  assign n5443 = n377 | n2178 ;
  assign n5444 = n2223 | n5443 ;
  assign n5445 = n5442 | n5444 ;
  assign n5446 = n159 | n3596 ;
  assign n5447 = n5445 | n5446 ;
  assign n5448 = n282 | n3676 ;
  assign n5449 = n127 | n5448 ;
  assign n5450 = n162 | n5449 ;
  assign n5451 = n5447 | n5450 ;
  assign n5452 = ~n2540 & n3886 ;
  assign n5453 = ( n516 & n2540 ) | ( n516 & n5452 ) | ( n2540 & n5452 );
  assign n5454 = ( ~n3886 & n5452 ) | ( ~n3886 & n5453 ) | ( n5452 & n5453 );
  assign n5455 = n516 & ~n3725 ;
  assign n5456 = ~n5322 & n5455 ;
  assign n5457 = n5395 & ~n5456 ;
  assign n5458 = ( n5402 & n5456 ) | ( n5402 & ~n5457 ) | ( n5456 & ~n5457 );
  assign n5459 = ( n5408 & ~n5454 ) | ( n5408 & n5458 ) | ( ~n5454 & n5458 );
  assign n5460 = ~n5454 & n5458 ;
  assign n5461 = ( ~n5405 & n5459 ) | ( ~n5405 & n5460 ) | ( n5459 & n5460 );
  assign n5462 = n5454 & ~n5458 ;
  assign n5463 = ( n5411 & ~n5461 ) | ( n5411 & n5462 ) | ( ~n5461 & n5462 );
  assign n5464 = ( n5413 & ~n5461 ) | ( n5413 & n5463 ) | ( ~n5461 & n5463 );
  assign n5465 = ~n5410 & n5411 ;
  assign n5466 = ( ~n5410 & n5413 ) | ( ~n5410 & n5465 ) | ( n5413 & n5465 );
  assign n5467 = ( n5458 & n5464 ) | ( n5458 & ~n5466 ) | ( n5464 & ~n5466 );
  assign n5468 = ( ~n5454 & n5464 ) | ( ~n5454 & n5467 ) | ( n5464 & n5467 );
  assign n5469 = n5451 & n5468 ;
  assign n5470 = n5451 | n5468 ;
  assign n5471 = n5417 & n5470 ;
  assign n5472 = ~n5469 & n5471 ;
  assign n5473 = ~n5469 & n5470 ;
  assign n5474 = ( n5425 & n5472 ) | ( n5425 & n5473 ) | ( n5472 & n5473 );
  assign n5475 = ( n5420 & n5472 ) | ( n5420 & n5473 ) | ( n5472 & n5473 );
  assign n5476 = ( n5419 & n5472 ) | ( n5419 & n5473 ) | ( n5472 & n5473 );
  assign n5477 = ( n5357 & n5475 ) | ( n5357 & n5476 ) | ( n5475 & n5476 );
  assign n5478 = ( n5142 & n5474 ) | ( n5142 & n5477 ) | ( n5474 & n5477 );
  assign n5479 = n5417 | n5425 ;
  assign n5480 = n5417 | n5420 ;
  assign n5481 = ( n5357 & n5418 ) | ( n5357 & n5480 ) | ( n5418 & n5480 );
  assign n5482 = ( n5142 & n5479 ) | ( n5142 & n5481 ) | ( n5479 & n5481 );
  assign n5483 = ~n5478 & n5482 ;
  assign n5484 = ~n5471 & n5473 ;
  assign n5485 = ~n5425 & n5484 ;
  assign n5486 = ~n5420 & n5484 ;
  assign n5487 = ~n5419 & n5484 ;
  assign n5488 = ( ~n5357 & n5486 ) | ( ~n5357 & n5487 ) | ( n5486 & n5487 );
  assign n5489 = ( ~n5142 & n5485 ) | ( ~n5142 & n5488 ) | ( n5485 & n5488 );
  assign n5490 = n5483 | n5489 ;
  assign n5491 = n5431 & n5490 ;
  assign n5492 = n5369 & n5491 ;
  assign n5493 = n5433 | n5490 ;
  assign n5494 = ~n5492 & n5493 ;
  assign n5495 = ( n3848 & n5436 ) | ( n3848 & n5438 ) | ( n5436 & n5438 );
  assign n5496 = ~n5494 & n5495 ;
  assign n5497 = n5494 & ~n5495 ;
  assign n5498 = n5496 | n5497 ;
  assign n5499 = n5436 | n5494 ;
  assign n5500 = n5437 | n5499 ;
  assign n5501 = n3848 & n5500 ;
  assign n5502 = n461 | n462 ;
  assign n5503 = n135 | n695 ;
  assign n5504 = n5502 | n5503 ;
  assign n5505 = n2022 | n2498 ;
  assign n5506 = n505 | n5505 ;
  assign n5507 = n5504 | n5506 ;
  assign n5508 = n283 | n2191 ;
  assign n5509 = n289 | n5508 ;
  assign n5510 = n109 | n5509 ;
  assign n5511 = n313 | n5510 ;
  assign n5512 = n5507 | n5511 ;
  assign n5513 = n384 | n5512 ;
  assign n5514 = n5469 & n5513 ;
  assign n5515 = ( n5471 & n5513 ) | ( n5471 & n5514 ) | ( n5513 & n5514 );
  assign n5516 = ( n5473 & n5513 ) | ( n5473 & n5514 ) | ( n5513 & n5514 );
  assign n5517 = ( n5425 & n5515 ) | ( n5425 & n5516 ) | ( n5515 & n5516 );
  assign n5518 = ( n5420 & n5515 ) | ( n5420 & n5516 ) | ( n5515 & n5516 );
  assign n5519 = ( n5419 & n5515 ) | ( n5419 & n5516 ) | ( n5515 & n5516 );
  assign n5520 = ( n5357 & n5518 ) | ( n5357 & n5519 ) | ( n5518 & n5519 );
  assign n5521 = ( n5142 & n5517 ) | ( n5142 & n5520 ) | ( n5517 & n5520 );
  assign n5522 = n5469 | n5513 ;
  assign n5523 = n5471 | n5522 ;
  assign n5524 = n5473 | n5522 ;
  assign n5525 = ( n5425 & n5523 ) | ( n5425 & n5524 ) | ( n5523 & n5524 );
  assign n5526 = ( n5420 & n5523 ) | ( n5420 & n5524 ) | ( n5523 & n5524 );
  assign n5527 = ( n5419 & n5523 ) | ( n5419 & n5524 ) | ( n5523 & n5524 );
  assign n5528 = ( n5357 & n5526 ) | ( n5357 & n5527 ) | ( n5526 & n5527 );
  assign n5529 = ( n5142 & n5525 ) | ( n5142 & n5528 ) | ( n5525 & n5528 );
  assign n5530 = ~n5521 & n5529 ;
  assign n5531 = n5431 & ~n5530 ;
  assign n5532 = n5490 & n5531 ;
  assign n5533 = n5369 & n5532 ;
  assign n5534 = n5530 | n5532 ;
  assign n5535 = ( n5369 & n5530 ) | ( n5369 & n5534 ) | ( n5530 & n5534 );
  assign n5536 = ( ~n5492 & n5533 ) | ( ~n5492 & n5535 ) | ( n5533 & n5535 );
  assign n5537 = n5501 & n5536 ;
  assign n5538 = n5501 | n5536 ;
  assign n5539 = ~n5537 & n5538 ;
  assign n5540 = n5500 | n5536 ;
  assign n5541 = n3848 & n5540 ;
  assign n5542 = n235 | n289 ;
  assign n5543 = n123 | n5542 ;
  assign n5544 = n161 | n473 ;
  assign n5545 = n2093 | n5544 ;
  assign n5546 = n425 | n5545 ;
  assign n5547 = n1083 | n5546 ;
  assign n5548 = n1025 | n5547 ;
  assign n5549 = n927 | n5548 ;
  assign n5550 = n225 | n5549 ;
  assign n5551 = n265 | n5550 ;
  assign n5552 = ( ~n3641 & n3643 ) | ( ~n3641 & n5551 ) | ( n3643 & n5551 );
  assign n5553 = n3641 | n5552 ;
  assign n5554 = n5543 | n5553 ;
  assign n5555 = n5515 | n5554 ;
  assign n5556 = n5516 | n5554 ;
  assign n5557 = ( n5425 & n5555 ) | ( n5425 & n5556 ) | ( n5555 & n5556 );
  assign n5558 = ( n5421 & n5555 ) | ( n5421 & n5556 ) | ( n5555 & n5556 );
  assign n5559 = ( n5142 & n5557 ) | ( n5142 & n5558 ) | ( n5557 & n5558 );
  assign n5560 = n5515 & n5554 ;
  assign n5561 = n5516 & n5554 ;
  assign n5562 = ( n5425 & n5560 ) | ( n5425 & n5561 ) | ( n5560 & n5561 );
  assign n5563 = ( n5421 & n5560 ) | ( n5421 & n5561 ) | ( n5560 & n5561 );
  assign n5564 = ( n5142 & n5562 ) | ( n5142 & n5563 ) | ( n5562 & n5563 );
  assign n5565 = n5559 & ~n5564 ;
  assign n5566 = n5530 | n5565 ;
  assign n5567 = ( n5491 & n5565 ) | ( n5491 & n5566 ) | ( n5565 & n5566 );
  assign n5568 = n5565 & n5566 ;
  assign n5569 = ( n5369 & n5567 ) | ( n5369 & n5568 ) | ( n5567 & n5568 );
  assign n5570 = n5530 & n5559 ;
  assign n5571 = n5569 & ~n5570 ;
  assign n5572 = ( ~n5492 & n5569 ) | ( ~n5492 & n5571 ) | ( n5569 & n5571 );
  assign n5573 = n5541 & ~n5572 ;
  assign n5574 = ~n5541 & n5572 ;
  assign n5575 = n5573 | n5574 ;
  assign n5576 = n5536 | n5572 ;
  assign n5577 = n5500 | n5576 ;
  assign n5578 = n3848 & n5577 ;
  assign n5579 = n5368 & n5570 ;
  assign n5580 = n5223 & n5579 ;
  assign n5581 = n129 | n4475 ;
  assign n5582 = n385 | n5581 ;
  assign n5583 = n5379 | n5582 ;
  assign n5584 = n126 | n891 ;
  assign n5585 = n2065 | n5584 ;
  assign n5586 = n5583 | n5585 ;
  assign n5587 = n181 | n221 ;
  assign n5588 = n282 | n5587 ;
  assign n5589 = n284 | n5588 ;
  assign n5590 = n134 | n5589 ;
  assign n5591 = n389 | n5590 ;
  assign n5592 = n556 | n5591 ;
  assign n5593 = n5586 | n5592 ;
  assign n5594 = n5554 & n5593 ;
  assign n5595 = n5515 & n5594 ;
  assign n5596 = n5516 & n5594 ;
  assign n5597 = ( n5425 & n5595 ) | ( n5425 & n5596 ) | ( n5595 & n5596 );
  assign n5598 = ( n5421 & n5595 ) | ( n5421 & n5596 ) | ( n5595 & n5596 );
  assign n5599 = ( n5142 & n5597 ) | ( n5142 & n5598 ) | ( n5597 & n5598 );
  assign n5600 = n5554 | n5593 ;
  assign n5601 = ( n5515 & n5593 ) | ( n5515 & n5600 ) | ( n5593 & n5600 );
  assign n5602 = ( n5516 & n5593 ) | ( n5516 & n5600 ) | ( n5593 & n5600 );
  assign n5603 = ( n5425 & n5601 ) | ( n5425 & n5602 ) | ( n5601 & n5602 );
  assign n5604 = ( n5421 & n5601 ) | ( n5421 & n5602 ) | ( n5601 & n5602 );
  assign n5605 = ( n5142 & n5603 ) | ( n5142 & n5604 ) | ( n5603 & n5604 );
  assign n5606 = ~n5599 & n5605 ;
  assign n5607 = ~n5491 & n5580 ;
  assign n5608 = ( n5580 & n5606 ) | ( n5580 & n5607 ) | ( n5606 & n5607 );
  assign n5609 = ( n5606 & n5607 ) | ( n5606 & ~n5608 ) | ( n5607 & ~n5608 );
  assign n5610 = ( n5580 & ~n5608 ) | ( n5580 & n5609 ) | ( ~n5608 & n5609 );
  assign n5611 = n5578 & ~n5610 ;
  assign n5612 = ~n5578 & n5610 ;
  assign n5613 = n5611 | n5612 ;
  assign n5614 = n5491 & n5570 ;
  assign n5615 = n186 | n329 ;
  assign n5616 = n559 | n4815 ;
  assign n5617 = n262 | n2024 ;
  assign n5618 = n5616 | n5617 ;
  assign n5619 = n265 | n268 ;
  assign n5620 = n5618 | n5619 ;
  assign n5621 = ( ~n944 & n5615 ) | ( ~n944 & n5620 ) | ( n5615 & n5620 );
  assign n5622 = n213 | n233 ;
  assign n5623 = n106 | n5622 ;
  assign n5624 = n944 | n5623 ;
  assign n5625 = n5621 | n5624 ;
  assign n5626 = n5594 | n5625 ;
  assign n5627 = ( n5515 & n5625 ) | ( n5515 & n5626 ) | ( n5625 & n5626 );
  assign n5628 = n383 | n5627 ;
  assign n5629 = ( n5516 & n5625 ) | ( n5516 & n5626 ) | ( n5625 & n5626 );
  assign n5630 = n383 | n5629 ;
  assign n5631 = ( n5425 & n5628 ) | ( n5425 & n5630 ) | ( n5628 & n5630 );
  assign n5632 = ( n5421 & n5628 ) | ( n5421 & n5630 ) | ( n5628 & n5630 );
  assign n5633 = ( n5142 & n5631 ) | ( n5142 & n5632 ) | ( n5631 & n5632 );
  assign n5634 = ( ~n5570 & n5606 ) | ( ~n5570 & n5633 ) | ( n5606 & n5633 );
  assign n5635 = n5606 | n5633 ;
  assign n5636 = ( ~n5491 & n5634 ) | ( ~n5491 & n5635 ) | ( n5634 & n5635 );
  assign n5637 = n5614 & n5636 ;
  assign n5638 = n5369 & n5637 ;
  assign n5639 = n5594 & n5625 ;
  assign n5640 = n5516 & n5639 ;
  assign n5641 = ( n383 & n5596 ) | ( n383 & n5640 ) | ( n5596 & n5640 );
  assign n5642 = n5515 & n5639 ;
  assign n5643 = ( n383 & n5595 ) | ( n383 & n5642 ) | ( n5595 & n5642 );
  assign n5644 = ( n5425 & n5641 ) | ( n5425 & n5643 ) | ( n5641 & n5643 );
  assign n5645 = ( n5421 & n5641 ) | ( n5421 & n5643 ) | ( n5641 & n5643 );
  assign n5646 = ( n5142 & n5644 ) | ( n5142 & n5645 ) | ( n5644 & n5645 );
  assign n5647 = n5633 & ~n5646 ;
  assign n5648 = n5606 | n5647 ;
  assign n5649 = ( n5570 & n5647 ) | ( n5570 & n5648 ) | ( n5647 & n5648 );
  assign n5650 = ( ~n5369 & n5491 ) | ( ~n5369 & n5649 ) | ( n5491 & n5649 );
  assign n5651 = ( n5369 & n5647 ) | ( n5369 & n5650 ) | ( n5647 & n5650 );
  assign n5652 = ~n5638 & n5651 ;
  assign n5653 = n5577 | n5610 ;
  assign n5654 = n3848 & n5653 ;
  assign n5655 = ~n5652 & n5654 ;
  assign n5656 = n5652 & ~n5654 ;
  assign n5657 = n5655 | n5656 ;
  assign n5658 = ( ~n261 & n351 ) | ( ~n261 & n2530 ) | ( n351 & n2530 );
  assign n5659 = n351 & n2530 ;
  assign n5660 = ( ~n309 & n5658 ) | ( ~n309 & n5659 ) | ( n5658 & n5659 );
  assign n5661 = n310 | n5660 ;
  assign n5662 = n323 | n5661 ;
  assign n5663 = n334 | n5662 ;
  assign n5664 = n5641 & n5663 ;
  assign n5665 = n5643 & n5663 ;
  assign n5666 = ( n5425 & n5664 ) | ( n5425 & n5665 ) | ( n5664 & n5665 );
  assign n5667 = ( n5421 & n5664 ) | ( n5421 & n5665 ) | ( n5664 & n5665 );
  assign n5668 = ( n5142 & n5666 ) | ( n5142 & n5667 ) | ( n5666 & n5667 );
  assign n5669 = n5641 | n5663 ;
  assign n5670 = n5643 | n5663 ;
  assign n5671 = ( n5425 & n5669 ) | ( n5425 & n5670 ) | ( n5669 & n5670 );
  assign n5672 = ( n5421 & n5669 ) | ( n5421 & n5670 ) | ( n5669 & n5670 );
  assign n5673 = ( n5142 & n5671 ) | ( n5142 & n5672 ) | ( n5671 & n5672 );
  assign n5674 = ~n5668 & n5673 ;
  assign n5675 = n5368 & n5674 ;
  assign n5676 = n5223 & n5675 ;
  assign n5677 = n5637 & n5676 ;
  assign n5678 = n5368 | n5674 ;
  assign n5679 = ( n5223 & n5674 ) | ( n5223 & n5678 ) | ( n5674 & n5678 );
  assign n5680 = ( n5637 & n5674 ) | ( n5637 & n5679 ) | ( n5674 & n5679 );
  assign n5681 = ~n5677 & n5680 ;
  assign n5682 = n5610 | n5652 ;
  assign n5683 = ( n3848 & n5578 ) | ( n3848 & n5682 ) | ( n5578 & n5682 );
  assign n5684 = ~n5681 & n5683 ;
  assign n5685 = n5681 & ~n5683 ;
  assign n5686 = n5684 | n5685 ;
  assign n5687 = n5652 | n5681 ;
  assign n5688 = n5610 | n5687 ;
  assign n5689 = ( n3848 & n5578 ) | ( n3848 & n5688 ) | ( n5578 & n5688 );
  assign n5690 = n310 | n568 ;
  assign n5691 = n5642 | n5690 ;
  assign n5692 = n5595 | n5690 ;
  assign n5693 = ( n383 & n5691 ) | ( n383 & n5692 ) | ( n5691 & n5692 );
  assign n5694 = ( n5663 & n5690 ) | ( n5663 & n5693 ) | ( n5690 & n5693 );
  assign n5695 = n5640 | n5690 ;
  assign n5696 = n5596 | n5690 ;
  assign n5697 = ( n383 & n5695 ) | ( n383 & n5696 ) | ( n5695 & n5696 );
  assign n5698 = ( n5663 & n5690 ) | ( n5663 & n5697 ) | ( n5690 & n5697 );
  assign n5699 = ( n5425 & n5694 ) | ( n5425 & n5698 ) | ( n5694 & n5698 );
  assign n5700 = ( n5421 & n5694 ) | ( n5421 & n5698 ) | ( n5694 & n5698 );
  assign n5701 = ( n5142 & n5699 ) | ( n5142 & n5700 ) | ( n5699 & n5700 );
  assign n5702 = n5676 & n5701 ;
  assign n5703 = ( ~n5637 & n5676 ) | ( ~n5637 & n5702 ) | ( n5676 & n5702 );
  assign n5704 = n5642 & n5690 ;
  assign n5705 = n5595 & n5690 ;
  assign n5706 = ( n383 & n5704 ) | ( n383 & n5705 ) | ( n5704 & n5705 );
  assign n5707 = n5663 & n5706 ;
  assign n5708 = n5640 & n5690 ;
  assign n5709 = n5596 & n5690 ;
  assign n5710 = ( n383 & n5708 ) | ( n383 & n5709 ) | ( n5708 & n5709 );
  assign n5711 = n5663 & n5710 ;
  assign n5712 = ( n5425 & n5707 ) | ( n5425 & n5711 ) | ( n5707 & n5711 );
  assign n5713 = ( n5421 & n5707 ) | ( n5421 & n5711 ) | ( n5707 & n5711 );
  assign n5714 = ( n5142 & n5712 ) | ( n5142 & n5713 ) | ( n5712 & n5713 );
  assign n5715 = n5701 & ~n5714 ;
  assign n5716 = ~n5676 & n5715 ;
  assign n5717 = ( ~n5637 & n5715 ) | ( ~n5637 & n5716 ) | ( n5715 & n5716 );
  assign n5718 = ( n5676 & ~n5703 ) | ( n5676 & n5717 ) | ( ~n5703 & n5717 );
  assign n5719 = n5689 & ~n5718 ;
  assign n5720 = ~n5689 & n5718 ;
  assign n5721 = n5719 | n5720 ;
  assign n5722 = n5701 | n5714 ;
  assign n5723 = ( ~n5676 & n5701 ) | ( ~n5676 & n5714 ) | ( n5701 & n5714 );
  assign n5724 = ( ~n5637 & n5722 ) | ( ~n5637 & n5723 ) | ( n5722 & n5723 );
  assign n5725 = n5677 & n5724 ;
  assign n5726 = ( n5676 & n5714 ) | ( n5676 & n5722 ) | ( n5714 & n5722 );
  assign n5727 = n5714 & n5722 ;
  assign n5728 = ( n5637 & n5726 ) | ( n5637 & n5727 ) | ( n5726 & n5727 );
  assign n5729 = ~n5725 & n5728 ;
  assign n5730 = n5688 | n5718 ;
  assign n5731 = ( n3848 & n5578 ) | ( n3848 & n5730 ) | ( n5578 & n5730 );
  assign n5732 = n5729 & n5731 ;
  assign n5733 = n51 | n53 ;
  assign n5734 = ( ~n5731 & n5732 ) | ( ~n5731 & n5733 ) | ( n5732 & n5733 );
  assign n5735 = ( ~n5729 & n5732 ) | ( ~n5729 & n5734 ) | ( n5732 & n5734 );
  assign n5736 = ~n53 & n3848 ;
  assign n5737 = ~n51 & n5736 ;
  assign n5738 = ~n5577 & n5728 ;
  assign n5739 = ( ~n5577 & n5730 ) | ( ~n5577 & n5738 ) | ( n5730 & n5738 );
  assign n5740 = n5577 & n5725 ;
  assign n5741 = ( n5725 & n5730 ) | ( n5725 & n5740 ) | ( n5730 & n5740 );
  assign n5742 = ( n5577 & n5739 ) | ( n5577 & ~n5741 ) | ( n5739 & ~n5741 );
  assign n5743 = ( n3848 & n5737 ) | ( n3848 & n5742 ) | ( n5737 & n5742 );
  assign po0 = n3845 ;
  assign po1 = n4025 ;
  assign po2 = n4164 ;
  assign po3 = n4311 ;
  assign po4 = n4468 ;
  assign po5 = n4596 ;
  assign po6 = n4707 ;
  assign po7 = n4799 ;
  assign po8 = n4895 ;
  assign po9 = n4990 ;
  assign po10 = n5084 ;
  assign po11 = n5153 ;
  assign po12 = n5229 ;
  assign po13 = n5306 ;
  assign po14 = n5376 ;
  assign po15 = n5441 ;
  assign po16 = n5498 ;
  assign po17 = n5539 ;
  assign po18 = n5575 ;
  assign po19 = n5613 ;
  assign po20 = n5657 ;
  assign po21 = n5686 ;
  assign po22 = n5721 ;
  assign po23 = ~n5735 ;
  assign po24 = n5743 ;
endmodule
