module top(G7 , G121 , G119 , G147 , G53 , G86 , G43 , G96 , G32 , G76 , G64 , G106 , G146 , G145 , G89 , G99 , G79 , G109 , G115 , G124 , G137 , G139 , G140 , G141 , G142 , G11 , G2 , G74 , G88 , G98 , G78 , G108 , G90 , G100 , G80 , G110 , G120 , G117 , G57 , G46 , G36 , G68 , G58 , G47 , G37 , G69 , G59 , G48 , G38 , G70 , G122 , G52 , G42 , G31 , G63 , G28 , G116 , G1 , G3 , G60 , G49 , G39 , G71 , G56 , G35 , G67 , G55 , G45 , G34 , G66 , G54 , G44 , G33 , G65 , G61 , G50 , G40 , G72 , G123 , G118 , G144 , G143 , G87 , G97 , G77 , G107 , G155 , G154 , G125 , G126 , G153 , G152 , G151 , G150 , G149 , G148 , G10 , G157 , G138 , G133 , G134 , G135 , G136 , G131 , G132 , G129 , G130 , G156 , G128 , G9 , G22 , G23 , G27 , G24 , G93 , G103 , G83 , G113 , G20 , G92 , G102 , G82 , G112 , G25 , G91 , G101 , G81 , G111 , G21 , G26 , G16 , G12 , G17 , G6 , G18 , G19 , G85 , G95 , G75 , G105 , G13 , G4 , G14 , G5 , G15 , G62 , G51 , G41 , G73 , G94 , G104 , G84 , G114 , G29 , G30 , G127 , G8 , G2551 , G2552 , G2553 , G2554 , G2555 , G2556 , G2557 , G2531 , G2532 , G2533 , G2534 , G2535 , G2536 , G2537 , G2538 , G2539 , G2540 , G2541 , G2542 , G2543 , G2544 , G2545 , G2546 , G2547 , G2548 , G2549 , G2550 , G2558 , G2559 , G2560 , G2561 , G2562 , G2563 , G2564 , G2565 , G2566 , G2567 , G2568 , G2569 , G2570 , G2571 , G2572 , G2573 , G2574 , G2575 , G2576 , G2577 , G2578 , G2579 , G2580 , G2581 , G2582 , G2583 , G2584 , G2585 , G2586 , G2587 , G2588 , G2589 , G2590 , G2591 , G2592 , G2593 , G2594 );
  input G7 , G121 , G119 , G147 , G53 , G86 , G43 , G96 , G32 , G76 , G64 , G106 , G146 , G145 , G89 , G99 , G79 , G109 , G115 , G124 , G137 , G139 , G140 , G141 , G142 , G11 , G2 , G74 , G88 , G98 , G78 , G108 , G90 , G100 , G80 , G110 , G120 , G117 , G57 , G46 , G36 , G68 , G58 , G47 , G37 , G69 , G59 , G48 , G38 , G70 , G122 , G52 , G42 , G31 , G63 , G28 , G116 , G1 , G3 , G60 , G49 , G39 , G71 , G56 , G35 , G67 , G55 , G45 , G34 , G66 , G54 , G44 , G33 , G65 , G61 , G50 , G40 , G72 , G123 , G118 , G144 , G143 , G87 , G97 , G77 , G107 , G155 , G154 , G125 , G126 , G153 , G152 , G151 , G150 , G149 , G148 , G10 , G157 , G138 , G133 , G134 , G135 , G136 , G131 , G132 , G129 , G130 , G156 , G128 , G9 , G22 , G23 , G27 , G24 , G93 , G103 , G83 , G113 , G20 , G92 , G102 , G82 , G112 , G25 , G91 , G101 , G81 , G111 , G21 , G26 , G16 , G12 , G17 , G6 , G18 , G19 , G85 , G95 , G75 , G105 , G13 , G4 , G14 , G5 , G15 , G62 , G51 , G41 , G73 , G94 , G104 , G84 , G114 , G29 , G30 , G127 , G8 ;
  output G2551 , G2552 , G2553 , G2554 , G2555 , G2556 , G2557 , G2531 , G2532 , G2533 , G2534 , G2535 , G2536 , G2537 , G2538 , G2539 , G2540 , G2541 , G2542 , G2543 , G2544 , G2545 , G2546 , G2547 , G2548 , G2549 , G2550 , G2558 , G2559 , G2560 , G2561 , G2562 , G2563 , G2564 , G2565 , G2566 , G2567 , G2568 , G2569 , G2570 , G2571 , G2572 , G2573 , G2574 , G2575 , G2576 , G2577 , G2578 , G2579 , G2580 , G2581 , G2582 , G2583 , G2584 , G2585 , G2586 , G2587 , G2588 , G2589 , G2590 , G2591 , G2592 , G2593 , G2594 ;
  wire n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702;
  assign n158 = G7 & G121 ;
  assign n159 = G119 & n158 ;
  assign n160 = G147 & n158 ;
  assign n161 = G53 & G43 ;
  assign n162 = G86 & n161 ;
  assign n163 = G96 & n162 ;
  assign n164 = G32 & G64 ;
  assign n165 = G76 & n164 ;
  assign n166 = G106 & n165 ;
  assign n167 = n163 & n166 ;
  assign n168 = G147 & ~n166 ;
  assign n169 = G119 & ~n163 ;
  assign n170 = n168 | n169 ;
  assign n171 = G146 | G145 ;
  assign n172 = G89 & ~n171 ;
  assign n173 = ~G146 & G145 ;
  assign n174 = G99 & n173 ;
  assign n175 = n172 | n174 ;
  assign n176 = G146 & ~G145 ;
  assign n177 = G79 & n176 ;
  assign n178 = G146 & G145 ;
  assign n179 = G109 & n178 ;
  assign n180 = n177 | n179 ;
  assign n181 = n175 | n180 ;
  assign n182 = G139 & G141 ;
  assign n183 = G140 & n182 ;
  assign n184 = G142 & n183 ;
  assign n185 = G121 & G2 ;
  assign n186 = G11 & n185 ;
  assign n187 = ~G115 & G74 ;
  assign n188 = G88 & ~n171 ;
  assign n189 = G108 & n178 ;
  assign n190 = G98 & n173 ;
  assign n191 = G78 & n176 ;
  assign n192 = n190 | n191 ;
  assign n193 = n189 | n192 ;
  assign n194 = n188 | n193 ;
  assign n195 = G80 & n176 ;
  assign n196 = G90 & ~n171 ;
  assign n197 = n195 | n196 ;
  assign n198 = G110 & n178 ;
  assign n199 = G100 & n173 ;
  assign n200 = n198 | n199 ;
  assign n201 = n197 | n200 ;
  assign n202 = G117 | G57 ;
  assign n203 = G117 & ~G46 ;
  assign n204 = G120 | n203 ;
  assign n205 = n202 & ~n204 ;
  assign n206 = G117 | G36 ;
  assign n207 = G117 & ~G68 ;
  assign n208 = G120 & ~n207 ;
  assign n209 = n206 & n208 ;
  assign n210 = n205 | n209 ;
  assign n211 = G117 | G37 ;
  assign n212 = G117 & ~G69 ;
  assign n213 = G120 & ~n212 ;
  assign n214 = n211 & n213 ;
  assign n215 = G117 | G58 ;
  assign n216 = G117 & ~G47 ;
  assign n217 = n215 & ~n216 ;
  assign n218 = ~G120 & n217 ;
  assign n219 = n214 | n218 ;
  assign n220 = G117 | G38 ;
  assign n221 = G117 & ~G70 ;
  assign n222 = G120 & ~n221 ;
  assign n223 = n220 & n222 ;
  assign n224 = G117 | G59 ;
  assign n225 = G117 & ~G48 ;
  assign n226 = n224 & ~n225 ;
  assign n227 = ~G120 & n226 ;
  assign n228 = n223 | n227 ;
  assign n229 = G117 | G31 ;
  assign n230 = G117 & ~G63 ;
  assign n231 = G120 & ~n230 ;
  assign n232 = n229 & n231 ;
  assign n233 = G117 | G52 ;
  assign n234 = G117 & ~G42 ;
  assign n235 = n233 & ~n234 ;
  assign n236 = ~G120 & n235 ;
  assign n237 = n232 | n236 ;
  assign n238 = G122 & n237 ;
  assign n239 = G122 & ~n238 ;
  assign n240 = ~G121 & G116 ;
  assign n241 = ~n170 & n240 ;
  assign n242 = G28 & n241 ;
  assign n243 = G1 & G3 ;
  assign n244 = n170 | n243 ;
  assign n245 = n240 & ~n244 ;
  assign n246 = G117 | G39 ;
  assign n247 = G117 & ~G71 ;
  assign n248 = G120 & ~n247 ;
  assign n249 = n246 & n248 ;
  assign n250 = G117 | G60 ;
  assign n251 = G117 & ~G49 ;
  assign n252 = n250 & ~n251 ;
  assign n253 = ~G120 & n252 ;
  assign n254 = n249 | n253 ;
  assign n255 = G120 | G117 ;
  assign n256 = G56 | n255 ;
  assign n257 = ~G117 & G35 ;
  assign n258 = G117 & G67 ;
  assign n259 = G120 & ~n258 ;
  assign n260 = ~n257 & n259 ;
  assign n261 = n256 & ~n260 ;
  assign n262 = G117 | G34 ;
  assign n263 = G117 & ~G66 ;
  assign n264 = G120 & ~n263 ;
  assign n265 = n262 & n264 ;
  assign n266 = G117 | G55 ;
  assign n267 = G117 & ~G45 ;
  assign n268 = n266 & ~n267 ;
  assign n269 = ~G120 & n268 ;
  assign n270 = n265 | n269 ;
  assign n271 = G117 | G33 ;
  assign n272 = G117 & ~G65 ;
  assign n273 = G120 & ~n272 ;
  assign n274 = n271 & n273 ;
  assign n275 = G117 | G54 ;
  assign n276 = G117 & ~G44 ;
  assign n277 = n275 & ~n276 ;
  assign n278 = ~G120 & n277 ;
  assign n279 = n274 | n278 ;
  assign n280 = G123 & ~n228 ;
  assign n281 = G117 | G40 ;
  assign n282 = G117 & ~G72 ;
  assign n283 = G120 & ~n282 ;
  assign n284 = n281 & n283 ;
  assign n285 = G117 | G61 ;
  assign n286 = G117 & ~G50 ;
  assign n287 = n285 & ~n286 ;
  assign n288 = ~G120 & n287 ;
  assign n289 = n284 | n288 ;
  assign n290 = ~G123 & n289 ;
  assign n291 = n280 | n290 ;
  assign n292 = G123 & ~n219 ;
  assign n293 = ~G123 & n254 ;
  assign n294 = n292 | n293 ;
  assign n295 = ~G122 & G118 ;
  assign n296 = n289 | n295 ;
  assign n297 = G118 | n289 ;
  assign n298 = G123 & n297 ;
  assign n299 = ~G123 & n237 ;
  assign n300 = n298 | n299 ;
  assign n301 = G107 & n178 ;
  assign n302 = G87 & ~n171 ;
  assign n303 = G77 & n176 ;
  assign n304 = G97 & n173 ;
  assign n305 = n303 | n304 ;
  assign n306 = n302 | n305 ;
  assign n307 = n301 | n306 ;
  assign n308 = G143 & n307 ;
  assign n309 = G143 | n307 ;
  assign n310 = ~G144 & n309 ;
  assign n311 = ~n308 & n310 ;
  assign n312 = ~G125 & G126 ;
  assign n313 = G125 & ~G126 ;
  assign n314 = n312 | n313 ;
  assign n315 = G155 | n314 ;
  assign n316 = G155 & n314 ;
  assign n317 = n315 & ~n316 ;
  assign n318 = ~G154 & n317 ;
  assign n319 = G154 & ~n317 ;
  assign n320 = n318 | n319 ;
  assign n321 = G149 & ~G148 ;
  assign n322 = ~G149 & G148 ;
  assign n323 = n321 | n322 ;
  assign n324 = ~G153 & G151 ;
  assign n325 = G153 & ~G151 ;
  assign n326 = n324 | n325 ;
  assign n327 = ~G152 & G150 ;
  assign n328 = G152 & ~G150 ;
  assign n329 = n327 | n328 ;
  assign n330 = n326 & ~n329 ;
  assign n331 = ~n326 & n329 ;
  assign n332 = n330 | n331 ;
  assign n333 = ~n323 & n332 ;
  assign n334 = n323 & ~n332 ;
  assign n335 = n333 | n334 ;
  assign n336 = n320 & ~n335 ;
  assign n337 = ~n320 & n335 ;
  assign n338 = n336 | n337 ;
  assign n339 = G10 & n338 ;
  assign n340 = ~G139 & G142 ;
  assign n341 = G139 & ~G142 ;
  assign n342 = n340 | n341 ;
  assign n343 = ~G140 & G141 ;
  assign n344 = G140 & ~G141 ;
  assign n345 = n343 | n344 ;
  assign n346 = ~G157 & G138 ;
  assign n347 = G157 & ~G138 ;
  assign n348 = n346 | n347 ;
  assign n349 = n345 & ~n348 ;
  assign n350 = ~n345 & n348 ;
  assign n351 = n349 | n350 ;
  assign n352 = n342 & ~n351 ;
  assign n353 = ~n342 & n351 ;
  assign n354 = n352 | n353 ;
  assign n355 = G144 | n354 ;
  assign n356 = G144 & n354 ;
  assign n357 = n355 & ~n356 ;
  assign n358 = ~G143 & n357 ;
  assign n359 = G143 & ~n357 ;
  assign n360 = n358 | n359 ;
  assign n361 = ~G133 & G135 ;
  assign n362 = G133 & ~G135 ;
  assign n363 = n361 | n362 ;
  assign n364 = G136 | n363 ;
  assign n365 = G136 & n363 ;
  assign n366 = n364 & ~n365 ;
  assign n367 = ~G134 & n366 ;
  assign n368 = G134 & ~n366 ;
  assign n369 = n367 | n368 ;
  assign n370 = ~G156 & G128 ;
  assign n371 = G156 & ~G128 ;
  assign n372 = n370 | n371 ;
  assign n373 = ~G131 & G129 ;
  assign n374 = G131 & ~G129 ;
  assign n375 = n373 | n374 ;
  assign n376 = ~G132 & G130 ;
  assign n377 = G132 & ~G130 ;
  assign n378 = n376 | n377 ;
  assign n379 = n375 & ~n378 ;
  assign n380 = ~n375 & n378 ;
  assign n381 = n379 | n380 ;
  assign n382 = ~n372 & n381 ;
  assign n383 = n372 & ~n381 ;
  assign n384 = n382 | n383 ;
  assign n385 = n369 & ~n384 ;
  assign n386 = ~n369 & n384 ;
  assign n387 = n385 | n386 ;
  assign n388 = G12 & G13 ;
  assign n389 = ~G12 & n237 ;
  assign n390 = n388 | n389 ;
  assign n391 = G125 & ~n390 ;
  assign n392 = G12 & G5 ;
  assign n393 = ~G12 & n228 ;
  assign n394 = n392 | n393 ;
  assign n395 = G129 & ~n394 ;
  assign n396 = G12 & G15 ;
  assign n397 = ~G12 & n219 ;
  assign n398 = n396 | n397 ;
  assign n399 = G130 | n398 ;
  assign n400 = G130 & n398 ;
  assign n401 = n399 & ~n400 ;
  assign n402 = n395 | n401 ;
  assign n403 = n391 | n402 ;
  assign n404 = ~G129 & n394 ;
  assign n405 = G12 & ~G14 ;
  assign n406 = G12 | n254 ;
  assign n407 = ~n405 & n406 ;
  assign n408 = G128 | n407 ;
  assign n409 = G128 & n407 ;
  assign n410 = n408 & ~n409 ;
  assign n411 = n404 | n410 ;
  assign n412 = ~G125 & n390 ;
  assign n413 = G12 & G4 ;
  assign n414 = ~G12 & n289 ;
  assign n415 = n413 | n414 ;
  assign n416 = G126 | n415 ;
  assign n417 = G126 & n415 ;
  assign n418 = n416 & ~n417 ;
  assign n419 = n412 | n418 ;
  assign n420 = n411 | n419 ;
  assign n421 = n403 | n420 ;
  assign n422 = G12 & G6 ;
  assign n423 = ~G12 & n270 ;
  assign n424 = n422 | n423 ;
  assign n425 = G133 & ~n424 ;
  assign n426 = G23 & ~G27 ;
  assign n427 = G23 | n194 ;
  assign n428 = ~n426 & n427 ;
  assign n429 = G142 | n428 ;
  assign n430 = G142 & n428 ;
  assign n431 = n429 & ~n430 ;
  assign n432 = n425 | n431 ;
  assign n433 = G23 & G19 ;
  assign n434 = G105 & n178 ;
  assign n435 = G75 & n176 ;
  assign n436 = G85 & ~n171 ;
  assign n437 = G95 & n173 ;
  assign n438 = n436 | n437 ;
  assign n439 = n435 | n438 ;
  assign n440 = n434 | n439 ;
  assign n441 = ~G23 & n440 ;
  assign n442 = n433 | n441 ;
  assign n443 = ~G135 & n442 ;
  assign n444 = ~G133 & n424 ;
  assign n445 = n443 | n444 ;
  assign n446 = n432 | n445 ;
  assign n447 = G135 & ~n442 ;
  assign n448 = G23 & G26 ;
  assign n449 = ~G23 & n181 ;
  assign n450 = n448 | n449 ;
  assign n451 = ~G141 & n450 ;
  assign n452 = G23 & G21 ;
  assign n453 = ~G23 & n201 ;
  assign n454 = n452 | n453 ;
  assign n455 = G140 & ~n454 ;
  assign n456 = G22 & G23 ;
  assign n457 = ~G23 & n307 ;
  assign n458 = n456 | n457 ;
  assign n459 = ~n455 & n458 ;
  assign n460 = ~n451 & n459 ;
  assign n461 = G23 & G20 ;
  assign n462 = G92 & ~n171 ;
  assign n463 = G102 & n173 ;
  assign n464 = n462 | n463 ;
  assign n465 = G82 & n176 ;
  assign n466 = G112 & n178 ;
  assign n467 = n465 | n466 ;
  assign n468 = n464 | n467 ;
  assign n469 = ~G23 & n468 ;
  assign n470 = n461 | n469 ;
  assign n471 = ~G138 & n470 ;
  assign n472 = G12 & ~G18 ;
  assign n473 = G12 | n279 ;
  assign n474 = ~n472 & n473 ;
  assign n475 = ~G134 & n474 ;
  assign n476 = G134 & ~n474 ;
  assign n477 = n475 | n476 ;
  assign n478 = n471 | n477 ;
  assign n479 = n460 & ~n478 ;
  assign n480 = G23 & G25 ;
  assign n481 = G91 & ~n171 ;
  assign n482 = G101 & n173 ;
  assign n483 = n481 | n482 ;
  assign n484 = G81 & n176 ;
  assign n485 = G111 & n178 ;
  assign n486 = n484 | n485 ;
  assign n487 = n483 | n486 ;
  assign n488 = ~G23 & n487 ;
  assign n489 = n480 | n488 ;
  assign n490 = G139 | n489 ;
  assign n491 = G139 & n489 ;
  assign n492 = n490 & ~n491 ;
  assign n493 = ~G140 & n454 ;
  assign n494 = n492 | n493 ;
  assign n495 = G23 & G24 ;
  assign n496 = G93 & ~n171 ;
  assign n497 = G103 & n173 ;
  assign n498 = n496 | n497 ;
  assign n499 = G83 & n176 ;
  assign n500 = G113 & n178 ;
  assign n501 = n499 | n500 ;
  assign n502 = n498 | n501 ;
  assign n503 = ~G23 & n502 ;
  assign n504 = n495 | n503 ;
  assign n505 = G136 | n504 ;
  assign n506 = G136 & n504 ;
  assign n507 = n505 & ~n506 ;
  assign n508 = G141 & ~n450 ;
  assign n509 = G138 & ~n470 ;
  assign n510 = n508 | n509 ;
  assign n511 = n507 | n510 ;
  assign n512 = n494 | n511 ;
  assign n513 = n479 & ~n512 ;
  assign n514 = ~n447 & n513 ;
  assign n515 = G12 & G17 ;
  assign n516 = ~G12 & n261 ;
  assign n517 = n515 | n516 ;
  assign n518 = G132 | n517 ;
  assign n519 = G132 & n517 ;
  assign n520 = n518 & ~n519 ;
  assign n521 = G12 | n210 ;
  assign n522 = ~G16 & G12 ;
  assign n523 = n521 & ~n522 ;
  assign n524 = G131 & ~n523 ;
  assign n525 = ~G131 & n523 ;
  assign n526 = n524 | n525 ;
  assign n527 = n520 | n526 ;
  assign n528 = n514 & ~n527 ;
  assign n529 = ~n446 & n528 ;
  assign n530 = G9 & n529 ;
  assign n531 = ~n421 & n530 ;
  assign n532 = G62 & ~n255 ;
  assign n533 = ~G120 & G51 ;
  assign n534 = G117 & n533 ;
  assign n535 = G117 & ~G73 ;
  assign n536 = G117 | G41 ;
  assign n537 = ~n535 & n536 ;
  assign n538 = G120 & n537 ;
  assign n539 = n534 | n538 ;
  assign n540 = n532 | n539 ;
  assign n541 = ~n237 & n540 ;
  assign n542 = n237 & ~n540 ;
  assign n543 = n541 | n542 ;
  assign n544 = ~n289 & n295 ;
  assign n545 = n238 | n544 ;
  assign n546 = ~n543 & n545 ;
  assign n547 = n543 & ~n545 ;
  assign n548 = n546 | n547 ;
  assign n549 = ~n440 & n468 ;
  assign n550 = n440 & ~n468 ;
  assign n551 = n549 | n550 ;
  assign n552 = ~n194 & n502 ;
  assign n553 = n194 & ~n502 ;
  assign n554 = n552 | n553 ;
  assign n555 = G114 & n178 ;
  assign n556 = G84 & n176 ;
  assign n557 = G104 & n173 ;
  assign n558 = G94 & ~n171 ;
  assign n559 = n557 | n558 ;
  assign n560 = n556 | n559 ;
  assign n561 = n555 | n560 ;
  assign n562 = n181 & ~n201 ;
  assign n563 = ~n181 & n201 ;
  assign n564 = n562 | n563 ;
  assign n565 = n561 & ~n564 ;
  assign n566 = ~n561 & n564 ;
  assign n567 = n565 | n566 ;
  assign n568 = n487 & ~n567 ;
  assign n569 = ~n487 & n567 ;
  assign n570 = n568 | n569 ;
  assign n571 = n554 & ~n570 ;
  assign n572 = ~n554 & n570 ;
  assign n573 = n571 | n572 ;
  assign n574 = n551 & ~n573 ;
  assign n575 = ~n551 & n573 ;
  assign n576 = n574 | n575 ;
  assign n577 = ~n307 & n576 ;
  assign n578 = n307 & ~n576 ;
  assign n579 = n577 | n578 ;
  assign n580 = ~G29 & n579 ;
  assign n581 = G123 | n540 ;
  assign n582 = n210 & ~n270 ;
  assign n583 = ~n210 & n270 ;
  assign n584 = n582 | n583 ;
  assign n585 = n261 & ~n279 ;
  assign n586 = ~n261 & n279 ;
  assign n587 = n585 | n586 ;
  assign n588 = n584 & ~n587 ;
  assign n589 = ~n584 & n587 ;
  assign n590 = n588 | n589 ;
  assign n591 = n254 & ~n289 ;
  assign n592 = ~n254 & n289 ;
  assign n593 = n591 | n592 ;
  assign n594 = ~n543 & n593 ;
  assign n595 = n543 & ~n593 ;
  assign n596 = n594 | n595 ;
  assign n597 = n297 & n596 ;
  assign n598 = n297 | n596 ;
  assign n599 = ~n597 & n598 ;
  assign n600 = n590 & n599 ;
  assign n601 = n590 | n599 ;
  assign n602 = ~n600 & n601 ;
  assign n603 = G123 & ~n602 ;
  assign n604 = n581 & ~n603 ;
  assign n605 = n219 & ~n228 ;
  assign n606 = ~n219 & n228 ;
  assign n607 = n605 | n606 ;
  assign n608 = n596 | n607 ;
  assign n609 = n596 & n607 ;
  assign n610 = n608 & ~n609 ;
  assign n611 = n590 | n610 ;
  assign n612 = n590 & n610 ;
  assign n613 = G29 | n612 ;
  assign n614 = n611 & ~n613 ;
  assign n615 = G30 & ~n181 ;
  assign n616 = ~G127 & n201 ;
  assign n617 = n615 & ~n616 ;
  assign n618 = ~n468 & n617 ;
  assign n619 = ~G138 & n617 ;
  assign n620 = ~n618 & n619 ;
  assign n621 = G135 | n440 ;
  assign n622 = n618 & ~n619 ;
  assign n623 = n620 | n622 ;
  assign n624 = n502 & n617 ;
  assign n625 = ~G136 & n617 ;
  assign n626 = ~n624 & n625 ;
  assign n627 = n624 & ~n625 ;
  assign n628 = n626 | n627 ;
  assign n629 = n623 | n628 ;
  assign n630 = n617 & ~n629 ;
  assign n631 = ~n621 & n630 ;
  assign n632 = ~n622 & n626 ;
  assign n633 = n631 | n632 ;
  assign n634 = n620 | n633 ;
  assign n635 = n261 & n270 ;
  assign n636 = n615 & n616 ;
  assign n637 = G8 & n636 ;
  assign n638 = ~n635 & n637 ;
  assign n639 = G8 & n210 ;
  assign n640 = G131 & ~n636 ;
  assign n641 = G142 & n636 ;
  assign n642 = n640 | n641 ;
  assign n643 = n639 & ~n642 ;
  assign n644 = G8 & ~n219 ;
  assign n645 = G141 & n636 ;
  assign n646 = G130 & ~n636 ;
  assign n647 = G8 & ~n646 ;
  assign n648 = ~n645 & n647 ;
  assign n649 = ~n644 & n648 ;
  assign n650 = G129 | n636 ;
  assign n651 = ~G140 & n636 ;
  assign n652 = n650 & ~n651 ;
  assign n653 = n228 & ~n652 ;
  assign n654 = n649 | n653 ;
  assign n655 = G126 | n636 ;
  assign n656 = ~G138 & n636 ;
  assign n657 = n655 & ~n656 ;
  assign n658 = n289 | n657 ;
  assign n659 = G128 | n636 ;
  assign n660 = ~G139 & n636 ;
  assign n661 = n659 & ~n660 ;
  assign n662 = n254 & ~n661 ;
  assign n663 = n658 & ~n662 ;
  assign n664 = n289 & n657 ;
  assign n665 = G136 & n636 ;
  assign n666 = G125 & ~n636 ;
  assign n667 = n237 | n666 ;
  assign n668 = n665 | n667 ;
  assign n669 = n664 | n668 ;
  assign n670 = n663 & n669 ;
  assign n671 = ~n254 & n661 ;
  assign n672 = ~n228 & n652 ;
  assign n673 = n671 | n672 ;
  assign n674 = n670 | n673 ;
  assign n675 = ~n654 & n674 ;
  assign n676 = G8 & n642 ;
  assign n677 = ~n210 & n676 ;
  assign n678 = n644 & ~n648 ;
  assign n679 = n677 | n678 ;
  assign n680 = n675 | n679 ;
  assign n681 = ~n643 & n680 ;
  assign n682 = n638 | n681 ;
  assign n683 = G133 & G132 ;
  assign n684 = G8 & ~n683 ;
  assign n685 = ~n636 & n684 ;
  assign n686 = n682 & ~n685 ;
  assign n687 = G134 | n686 ;
  assign n688 = ~n279 & n687 ;
  assign n689 = G135 & n440 ;
  assign n690 = n621 & ~n689 ;
  assign n691 = ~n688 & n690 ;
  assign n692 = n617 & ~n691 ;
  assign n693 = ~G134 & n617 ;
  assign n694 = n686 & ~n693 ;
  assign n695 = n629 | n694 ;
  assign n696 = n692 | n695 ;
  assign n697 = ~n634 & n696 ;
  assign n698 = n339 | n614 ;
  assign n699 = n360 & n387 ;
  assign n700 = ~n170 & n699 ;
  assign n701 = ~n698 & n700 ;
  assign n702 = ~n580 & n701 ;
  assign G2551 = ~n158 ;
  assign G2552 = ~n159 ;
  assign G2553 = ~n160 ;
  assign G2554 = ~n167 ;
  assign G2555 = ~n167 ;
  assign G2556 = n170 ;
  assign G2557 = ~n181 ;
  assign G2531 = ~G115 ;
  assign G2532 = ~G115 ;
  assign G2533 = ~G115 ;
  assign G2534 = ~G124 ;
  assign G2535 = ~G124 ;
  assign G2536 = ~G137 ;
  assign G2537 = ~G137 ;
  assign G2538 = ~G137 ;
  assign G2539 = ~G32 ;
  assign G2540 = ~G106 ;
  assign G2541 = ~G64 ;
  assign G2542 = ~G76 ;
  assign G2543 = ~G53 ;
  assign G2544 = ~G96 ;
  assign G2545 = ~G43 ;
  assign G2546 = ~G86 ;
  assign G2547 = ~n184 ;
  assign G2548 = ~n186 ;
  assign G2549 = G115 ;
  assign G2550 = n187 ;
  assign G2558 = ~n194 ;
  assign G2559 = ~n201 ;
  assign G2560 = ~n210 ;
  assign G2561 = ~n219 ;
  assign G2562 = ~n228 ;
  assign G2563 = ~n239 ;
  assign G2564 = ~n242 ;
  assign G2565 = ~n245 ;
  assign G2566 = n254 ;
  assign G2567 = n228 ;
  assign G2568 = n219 ;
  assign G2569 = n210 ;
  assign G2570 = n261 ;
  assign G2571 = n270 ;
  assign G2572 = n279 ;
  assign G2573 = ~n291 ;
  assign G2574 = ~n291 ;
  assign G2575 = n294 ;
  assign G2576 = n294 ;
  assign G2577 = n296 ;
  assign G2578 = ~n300 ;
  assign G2579 = ~n300 ;
  assign G2580 = ~n311 ;
  assign G2581 = ~n339 ;
  assign G2582 = ~n360 ;
  assign G2583 = ~n387 ;
  assign G2584 = ~n531 ;
  assign G2585 = ~n531 ;
  assign G2586 = n548 ;
  assign G2587 = ~n580 ;
  assign G2588 = n604 ;
  assign G2589 = n604 ;
  assign G2590 = ~n614 ;
  assign G2591 = n697 ;
  assign G2592 = 1'b0 ;
  assign G2593 = ~n702 ;
  assign G2594 = ~n702 ;
endmodule
