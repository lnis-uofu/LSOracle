module top(G1 , G5 , G9 , G13 , G33 , G41 , G17 , G18 , G19 , G20 , G21 , G22 , G23 , G24 , G4 , G8 , G12 , G16 , G36 , G29 , G30 , G31 , G32 , G3 , G7 , G11 , G15 , G35 , G25 , G26 , G27 , G28 , G2 , G6 , G10 , G14 , G34 , G40 , G39 , G38 , G37 , G1324 , G1344 , G1325 , G1326 , G1327 , G1328 , G1329 , G1330 , G1343 , G1331 , G1332 , G1333 , G1334 , G1335 , G1336 , G1337 , G1338 , G1339 , G1340 , G1341 , G1342 , G1345 , G1346 , G1347 , G1348 , G1349 , G1350 , G1351 , G1352 , G1353 , G1354 , G1355 );
  input G1 , G5 , G9 , G13 , G33 , G41 , G17 , G18 , G19 , G20 , G21 , G22 , G23 , G24 , G4 , G8 , G12 , G16 , G36 , G29 , G30 , G31 , G32 , G3 , G7 , G11 , G15 , G35 , G25 , G26 , G27 , G28 , G2 , G6 , G10 , G14 , G34 , G40 , G39 , G38 , G37 ;
  output G1324 , G1344 , G1325 , G1326 , G1327 , G1328 , G1329 , G1330 , G1343 , G1331 , G1332 , G1333 , G1334 , G1335 , G1336 , G1337 , G1338 , G1339 , G1340 , G1341 , G1342 , G1345 , G1346 , G1347 , G1348 , G1349 , G1350 , G1351 , G1352 , G1353 , G1354 , G1355 ;
  wire n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491;
  assign n42 = G4 & ~G12 ;
  assign n43 = ( ~G4 & G12 ) | ( ~G4 & n42 ) | ( G12 & n42 );
  assign n44 = n42 | n43 ;
  assign n45 = ( G8 & ~G16 ) | ( G8 & n42 ) | ( ~G16 & n42 );
  assign n46 = ~G8 & G16 ;
  assign n47 = ( n43 & n45 ) | ( n43 & ~n46 ) | ( n45 & ~n46 );
  assign n48 = ( ~G8 & G16 ) | ( ~G8 & n42 ) | ( G16 & n42 );
  assign n49 = G8 & ~G16 ;
  assign n50 = ( n43 & n48 ) | ( n43 & ~n49 ) | ( n48 & ~n49 );
  assign n51 = ( ~n44 & n47 ) | ( ~n44 & n50 ) | ( n47 & n50 );
  assign n52 = G21 & ~G23 ;
  assign n53 = ( ~G21 & G23 ) | ( ~G21 & n52 ) | ( G23 & n52 );
  assign n54 = n52 | n53 ;
  assign n55 = ( G22 & ~G24 ) | ( G22 & n54 ) | ( ~G24 & n54 );
  assign n56 = ( ~G22 & G24 ) | ( ~G22 & n54 ) | ( G24 & n54 );
  assign n57 = ( ~n54 & n55 ) | ( ~n54 & n56 ) | ( n55 & n56 );
  assign n58 = n51 | n57 ;
  assign n59 = ( n51 & n57 ) | ( n51 & ~n58 ) | ( n57 & ~n58 );
  assign n60 = n58 & ~n59 ;
  assign n61 = G41 & G36 ;
  assign n62 = G29 & ~G31 ;
  assign n63 = ( ~G29 & G31 ) | ( ~G29 & n62 ) | ( G31 & n62 );
  assign n64 = n62 | n63 ;
  assign n65 = ( G30 & ~G32 ) | ( G30 & n64 ) | ( ~G32 & n64 );
  assign n66 = ( ~G30 & G32 ) | ( ~G30 & n64 ) | ( G32 & n64 );
  assign n67 = ( ~n64 & n65 ) | ( ~n64 & n66 ) | ( n65 & n66 );
  assign n68 = n61 & n67 ;
  assign n69 = n61 | n67 ;
  assign n70 = ( n57 & n61 ) | ( n57 & n67 ) | ( n61 & n67 );
  assign n71 = ( n51 & n69 ) | ( n51 & n70 ) | ( n69 & n70 );
  assign n72 = ( ~n59 & n68 ) | ( ~n59 & n71 ) | ( n68 & n71 );
  assign n73 = ( ~n57 & n61 ) | ( ~n57 & n67 ) | ( n61 & n67 );
  assign n74 = ( ~n51 & n68 ) | ( ~n51 & n73 ) | ( n68 & n73 );
  assign n75 = ( n59 & n69 ) | ( n59 & n74 ) | ( n69 & n74 );
  assign n76 = ( n60 & ~n72 ) | ( n60 & n75 ) | ( ~n72 & n75 );
  assign n77 = G3 & ~G11 ;
  assign n78 = ( ~G3 & G11 ) | ( ~G3 & n77 ) | ( G11 & n77 );
  assign n79 = n77 | n78 ;
  assign n80 = ( G7 & ~G15 ) | ( G7 & n77 ) | ( ~G15 & n77 );
  assign n81 = ~G7 & G15 ;
  assign n82 = ( n78 & n80 ) | ( n78 & ~n81 ) | ( n80 & ~n81 );
  assign n83 = ( ~G7 & G15 ) | ( ~G7 & n77 ) | ( G15 & n77 );
  assign n84 = G7 & ~G15 ;
  assign n85 = ( n78 & n83 ) | ( n78 & ~n84 ) | ( n83 & ~n84 );
  assign n86 = ( ~n79 & n82 ) | ( ~n79 & n85 ) | ( n82 & n85 );
  assign n87 = G17 & ~G19 ;
  assign n88 = ( ~G17 & G19 ) | ( ~G17 & n87 ) | ( G19 & n87 );
  assign n89 = n87 | n88 ;
  assign n90 = ( G18 & ~G20 ) | ( G18 & n89 ) | ( ~G20 & n89 );
  assign n91 = ( ~G18 & G20 ) | ( ~G18 & n89 ) | ( G20 & n89 );
  assign n92 = ( ~n89 & n90 ) | ( ~n89 & n91 ) | ( n90 & n91 );
  assign n93 = n86 | n92 ;
  assign n94 = ( n86 & n92 ) | ( n86 & ~n93 ) | ( n92 & ~n93 );
  assign n95 = n93 & ~n94 ;
  assign n96 = G41 & G35 ;
  assign n97 = G25 & ~G27 ;
  assign n98 = ( ~G25 & G27 ) | ( ~G25 & n97 ) | ( G27 & n97 );
  assign n99 = n97 | n98 ;
  assign n100 = ( G26 & ~G28 ) | ( G26 & n99 ) | ( ~G28 & n99 );
  assign n101 = ( ~G26 & G28 ) | ( ~G26 & n99 ) | ( G28 & n99 );
  assign n102 = ( ~n99 & n100 ) | ( ~n99 & n101 ) | ( n100 & n101 );
  assign n103 = n96 & n102 ;
  assign n104 = n96 | n102 ;
  assign n105 = ( n92 & n96 ) | ( n92 & n102 ) | ( n96 & n102 );
  assign n106 = ( n86 & n104 ) | ( n86 & n105 ) | ( n104 & n105 );
  assign n107 = ( ~n94 & n103 ) | ( ~n94 & n106 ) | ( n103 & n106 );
  assign n108 = ( ~n92 & n96 ) | ( ~n92 & n102 ) | ( n96 & n102 );
  assign n109 = ( ~n86 & n103 ) | ( ~n86 & n108 ) | ( n103 & n108 );
  assign n110 = ( n94 & n104 ) | ( n94 & n109 ) | ( n104 & n109 );
  assign n111 = ( n95 & ~n107 ) | ( n95 & n110 ) | ( ~n107 & n110 );
  assign n112 = ~n76 & n111 ;
  assign n113 = n76 | n111 ;
  assign n114 = G1 & ~G9 ;
  assign n115 = ( ~G1 & G9 ) | ( ~G1 & n114 ) | ( G9 & n114 );
  assign n116 = n114 | n115 ;
  assign n117 = ( G5 & ~G13 ) | ( G5 & n114 ) | ( ~G13 & n114 );
  assign n118 = ~G5 & G13 ;
  assign n119 = ( n115 & n117 ) | ( n115 & ~n118 ) | ( n117 & ~n118 );
  assign n120 = ( ~G5 & G13 ) | ( ~G5 & n114 ) | ( G13 & n114 );
  assign n121 = G5 & ~G13 ;
  assign n122 = ( n115 & n120 ) | ( n115 & ~n121 ) | ( n120 & ~n121 );
  assign n123 = ( ~n116 & n119 ) | ( ~n116 & n122 ) | ( n119 & n122 );
  assign n124 = n92 | n123 ;
  assign n125 = ( n92 & n123 ) | ( n92 & ~n124 ) | ( n123 & ~n124 );
  assign n126 = n124 & ~n125 ;
  assign n127 = G33 & G41 ;
  assign n128 = n57 & n127 ;
  assign n129 = n57 | n127 ;
  assign n130 = ( n57 & n92 ) | ( n57 & n127 ) | ( n92 & n127 );
  assign n131 = ( n123 & n129 ) | ( n123 & n130 ) | ( n129 & n130 );
  assign n132 = ( ~n125 & n128 ) | ( ~n125 & n131 ) | ( n128 & n131 );
  assign n133 = ( n57 & ~n92 ) | ( n57 & n127 ) | ( ~n92 & n127 );
  assign n134 = ( ~n123 & n128 ) | ( ~n123 & n133 ) | ( n128 & n133 );
  assign n135 = ( n125 & n129 ) | ( n125 & n134 ) | ( n129 & n134 );
  assign n136 = ( n126 & ~n132 ) | ( n126 & n135 ) | ( ~n132 & n135 );
  assign n137 = G2 & ~G10 ;
  assign n138 = ( ~G2 & G10 ) | ( ~G2 & n137 ) | ( G10 & n137 );
  assign n139 = n137 | n138 ;
  assign n140 = ( G6 & ~G14 ) | ( G6 & n137 ) | ( ~G14 & n137 );
  assign n141 = ~G6 & G14 ;
  assign n142 = ( n138 & n140 ) | ( n138 & ~n141 ) | ( n140 & ~n141 );
  assign n143 = ( ~G6 & G14 ) | ( ~G6 & n137 ) | ( G14 & n137 );
  assign n144 = G6 & ~G14 ;
  assign n145 = ( n138 & n143 ) | ( n138 & ~n144 ) | ( n143 & ~n144 );
  assign n146 = ( ~n139 & n142 ) | ( ~n139 & n145 ) | ( n142 & n145 );
  assign n147 = n67 | n146 ;
  assign n148 = ( n67 & n146 ) | ( n67 & ~n147 ) | ( n146 & ~n147 );
  assign n149 = n147 & ~n148 ;
  assign n150 = G41 & G34 ;
  assign n151 = n102 & n150 ;
  assign n152 = n102 | n150 ;
  assign n153 = ( n67 & n102 ) | ( n67 & n150 ) | ( n102 & n150 );
  assign n154 = ( n146 & n152 ) | ( n146 & n153 ) | ( n152 & n153 );
  assign n155 = ( ~n148 & n151 ) | ( ~n148 & n154 ) | ( n151 & n154 );
  assign n156 = ( ~n67 & n102 ) | ( ~n67 & n150 ) | ( n102 & n150 );
  assign n157 = ( ~n146 & n151 ) | ( ~n146 & n156 ) | ( n151 & n156 );
  assign n158 = ( n148 & n152 ) | ( n148 & n157 ) | ( n152 & n157 );
  assign n159 = ( n149 & ~n155 ) | ( n149 & n158 ) | ( ~n155 & n158 );
  assign n160 = ( n113 & n136 ) | ( n113 & n159 ) | ( n136 & n159 );
  assign n161 = n136 | n159 ;
  assign n162 = ( n76 & ~n111 ) | ( n76 & n161 ) | ( ~n111 & n161 );
  assign n163 = ( n112 & ~n160 ) | ( n112 & n162 ) | ( ~n160 & n162 );
  assign n164 = G13 & ~G15 ;
  assign n165 = ( ~G13 & G15 ) | ( ~G13 & n164 ) | ( G15 & n164 );
  assign n166 = n164 | n165 ;
  assign n167 = ( G16 & ~G14 ) | ( G16 & n164 ) | ( ~G14 & n164 );
  assign n168 = ~G16 & G14 ;
  assign n169 = ( n165 & n167 ) | ( n165 & ~n168 ) | ( n167 & ~n168 );
  assign n170 = ( ~G16 & G14 ) | ( ~G16 & n164 ) | ( G14 & n164 );
  assign n171 = G16 & ~G14 ;
  assign n172 = ( n165 & n170 ) | ( n165 & ~n171 ) | ( n170 & ~n171 );
  assign n173 = ( ~n166 & n169 ) | ( ~n166 & n172 ) | ( n169 & n172 );
  assign n174 = G41 & G40 ;
  assign n175 = G5 & ~G7 ;
  assign n176 = ( ~G5 & G7 ) | ( ~G5 & n175 ) | ( G7 & n175 );
  assign n177 = n175 | n176 ;
  assign n178 = ( G8 & ~G6 ) | ( G8 & n177 ) | ( ~G6 & n177 );
  assign n179 = ( ~G8 & G6 ) | ( ~G8 & n177 ) | ( G6 & n177 );
  assign n180 = ( ~n177 & n178 ) | ( ~n177 & n179 ) | ( n178 & n179 );
  assign n181 = ( n173 & n174 ) | ( n173 & ~n180 ) | ( n174 & ~n180 );
  assign n182 = ( ~n174 & n180 ) | ( ~n174 & n181 ) | ( n180 & n181 );
  assign n183 = ( ~n173 & n181 ) | ( ~n173 & n182 ) | ( n181 & n182 );
  assign n184 = G20 & ~G32 ;
  assign n185 = ( ~G20 & G32 ) | ( ~G20 & n184 ) | ( G32 & n184 );
  assign n186 = n184 | n185 ;
  assign n187 = ( G24 & ~G28 ) | ( G24 & n184 ) | ( ~G28 & n184 );
  assign n188 = ~G24 & G28 ;
  assign n189 = ( n185 & n187 ) | ( n185 & ~n188 ) | ( n187 & ~n188 );
  assign n190 = ( ~G24 & G28 ) | ( ~G24 & n184 ) | ( G28 & n184 );
  assign n191 = G24 & ~G28 ;
  assign n192 = ( n185 & n190 ) | ( n185 & ~n191 ) | ( n190 & ~n191 );
  assign n193 = ( ~n186 & n189 ) | ( ~n186 & n192 ) | ( n189 & n192 );
  assign n194 = n183 & ~n193 ;
  assign n195 = ~n183 & n193 ;
  assign n196 = n194 | n195 ;
  assign n197 = n136 & ~n196 ;
  assign n198 = G41 & G38 ;
  assign n199 = G9 & ~G11 ;
  assign n200 = ( ~G9 & G11 ) | ( ~G9 & n199 ) | ( G11 & n199 );
  assign n201 = n199 | n200 ;
  assign n202 = ( G12 & ~G10 ) | ( G12 & n199 ) | ( ~G10 & n199 );
  assign n203 = ~G12 & G10 ;
  assign n204 = ( n200 & n202 ) | ( n200 & ~n203 ) | ( n202 & ~n203 );
  assign n205 = ( ~G12 & G10 ) | ( ~G12 & n199 ) | ( G10 & n199 );
  assign n206 = G12 & ~G10 ;
  assign n207 = ( n200 & n205 ) | ( n200 & ~n206 ) | ( n205 & ~n206 );
  assign n208 = ( ~n201 & n204 ) | ( ~n201 & n207 ) | ( n204 & n207 );
  assign n209 = ~n173 & n208 ;
  assign n210 = n173 | n209 ;
  assign n211 = ~n198 & n209 ;
  assign n212 = n198 | n208 ;
  assign n213 = ( n210 & n211 ) | ( n210 & ~n212 ) | ( n211 & ~n212 );
  assign n214 = ( ~n208 & n209 ) | ( ~n208 & n210 ) | ( n209 & n210 );
  assign n215 = G18 & ~G30 ;
  assign n216 = ( ~G18 & G30 ) | ( ~G18 & n215 ) | ( G30 & n215 );
  assign n217 = n215 | n216 ;
  assign n218 = ( G22 & ~G26 ) | ( G22 & n217 ) | ( ~G26 & n217 );
  assign n219 = ( ~G22 & G26 ) | ( ~G22 & n217 ) | ( G26 & n217 );
  assign n220 = ( ~n217 & n218 ) | ( ~n217 & n219 ) | ( n218 & n219 );
  assign n221 = ( ~n213 & n214 ) | ( ~n213 & n220 ) | ( n214 & n220 );
  assign n222 = ( n198 & n213 ) | ( n198 & ~n221 ) | ( n213 & ~n221 );
  assign n223 = ( ~n198 & n209 ) | ( ~n198 & n220 ) | ( n209 & n220 );
  assign n224 = ( n198 & n208 ) | ( n198 & ~n220 ) | ( n208 & ~n220 );
  assign n225 = ( n210 & n223 ) | ( n210 & ~n224 ) | ( n223 & ~n224 );
  assign n226 = ~n213 & n225 ;
  assign n227 = G41 & G37 ;
  assign n228 = G1 & ~G3 ;
  assign n229 = ( ~G1 & G3 ) | ( ~G1 & n228 ) | ( G3 & n228 );
  assign n230 = n228 | n229 ;
  assign n231 = ( G4 & ~G2 ) | ( G4 & n230 ) | ( ~G2 & n230 );
  assign n232 = ( ~G4 & G2 ) | ( ~G4 & n230 ) | ( G2 & n230 );
  assign n233 = ( ~n230 & n231 ) | ( ~n230 & n232 ) | ( n231 & n232 );
  assign n234 = ( n180 & n227 ) | ( n180 & ~n233 ) | ( n227 & ~n233 );
  assign n235 = ( ~n180 & n233 ) | ( ~n180 & n234 ) | ( n233 & n234 );
  assign n236 = ( ~n227 & n234 ) | ( ~n227 & n235 ) | ( n234 & n235 );
  assign n237 = G17 & ~G29 ;
  assign n238 = ( ~G17 & G29 ) | ( ~G17 & n237 ) | ( G29 & n237 );
  assign n239 = n237 | n238 ;
  assign n240 = ( G21 & ~G25 ) | ( G21 & n237 ) | ( ~G25 & n237 );
  assign n241 = ~G21 & G25 ;
  assign n242 = ( n238 & n240 ) | ( n238 & ~n241 ) | ( n240 & ~n241 );
  assign n243 = ( ~G21 & G25 ) | ( ~G21 & n237 ) | ( G25 & n237 );
  assign n244 = G21 & ~G25 ;
  assign n245 = ( n238 & n243 ) | ( n238 & ~n244 ) | ( n243 & ~n244 );
  assign n246 = ( ~n239 & n242 ) | ( ~n239 & n245 ) | ( n242 & n245 );
  assign n247 = n236 & ~n246 ;
  assign n248 = ~n236 & n246 ;
  assign n249 = n247 | n248 ;
  assign n250 = ~n226 & n249 ;
  assign n251 = ~n222 & n250 ;
  assign n252 = G41 & G39 ;
  assign n253 = ( n208 & ~n233 ) | ( n208 & n252 ) | ( ~n233 & n252 );
  assign n254 = ( n233 & ~n252 ) | ( n233 & n253 ) | ( ~n252 & n253 );
  assign n255 = ( ~n208 & n253 ) | ( ~n208 & n254 ) | ( n253 & n254 );
  assign n256 = G19 & ~G31 ;
  assign n257 = ( ~G19 & G31 ) | ( ~G19 & n256 ) | ( G31 & n256 );
  assign n258 = n256 | n257 ;
  assign n259 = ( G23 & ~G27 ) | ( G23 & n256 ) | ( ~G27 & n256 );
  assign n260 = ~G23 & G27 ;
  assign n261 = ( n257 & n259 ) | ( n257 & ~n260 ) | ( n259 & ~n260 );
  assign n262 = ( ~G23 & G27 ) | ( ~G23 & n256 ) | ( G27 & n256 );
  assign n263 = G23 & ~G27 ;
  assign n264 = ( n257 & n262 ) | ( n257 & ~n263 ) | ( n262 & ~n263 );
  assign n265 = ( ~n258 & n261 ) | ( ~n258 & n264 ) | ( n261 & n264 );
  assign n266 = n255 & ~n265 ;
  assign n267 = ~n255 & n265 ;
  assign n268 = n266 | n267 ;
  assign n269 = n251 & n268 ;
  assign n270 = n197 & n269 ;
  assign n271 = n163 & n270 ;
  assign n272 = G1 & ~n271 ;
  assign n273 = ~G1 & n271 ;
  assign n274 = n272 | n273 ;
  assign n275 = n136 & ~n159 ;
  assign n276 = ~n111 & n275 ;
  assign n277 = n76 & n276 ;
  assign n278 = ( n196 & n213 ) | ( n196 & n268 ) | ( n213 & n268 );
  assign n279 = ( n196 & n198 ) | ( n196 & n268 ) | ( n198 & n268 );
  assign n280 = ( ~n221 & n278 ) | ( ~n221 & n279 ) | ( n278 & n279 );
  assign n281 = ( n196 & ~n249 ) | ( n196 & n268 ) | ( ~n249 & n268 );
  assign n282 = n196 & n268 ;
  assign n283 = ( ~n226 & n281 ) | ( ~n226 & n282 ) | ( n281 & n282 );
  assign n284 = ~n280 & n283 ;
  assign n285 = n196 | n268 ;
  assign n286 = ( ~n198 & n209 ) | ( ~n198 & n249 ) | ( n209 & n249 );
  assign n287 = ( n198 & n208 ) | ( n198 & ~n249 ) | ( n208 & ~n249 );
  assign n288 = ( n210 & n286 ) | ( n210 & ~n287 ) | ( n286 & ~n287 );
  assign n289 = n225 & ~n288 ;
  assign n290 = ( n222 & ~n249 ) | ( n222 & n289 ) | ( ~n249 & n289 );
  assign n291 = ( n251 & ~n285 ) | ( n251 & n290 ) | ( ~n285 & n290 );
  assign n292 = n284 | n291 ;
  assign n293 = n277 & n292 ;
  assign n294 = n249 & n293 ;
  assign n295 = G21 & n293 ;
  assign n296 = n249 & n295 ;
  assign n297 = G21 & ~n295 ;
  assign n298 = ( G21 & ~n249 ) | ( G21 & n297 ) | ( ~n249 & n297 );
  assign n299 = ( n294 & ~n296 ) | ( n294 & n298 ) | ( ~n296 & n298 );
  assign n300 = n163 & ~n196 ;
  assign n301 = n159 & n269 ;
  assign n302 = n300 & n301 ;
  assign n303 = ~G2 & n302 ;
  assign n304 = G2 | n302 ;
  assign n305 = ( ~n302 & n303 ) | ( ~n302 & n304 ) | ( n303 & n304 );
  assign n306 = n111 & n269 ;
  assign n307 = n300 & n306 ;
  assign n308 = ~G3 & n307 ;
  assign n309 = G3 | n307 ;
  assign n310 = ( ~n307 & n308 ) | ( ~n307 & n309 ) | ( n308 & n309 );
  assign n311 = n76 & n269 ;
  assign n312 = n300 & n311 ;
  assign n313 = ~G4 & n312 ;
  assign n314 = G4 | n312 ;
  assign n315 = ( ~n312 & n313 ) | ( ~n312 & n314 ) | ( n313 & n314 );
  assign n316 = n163 & n196 ;
  assign n317 = n213 | n268 ;
  assign n318 = n198 | n268 ;
  assign n319 = ( ~n221 & n317 ) | ( ~n221 & n318 ) | ( n317 & n318 );
  assign n320 = ( n196 & ~n250 ) | ( n196 & n319 ) | ( ~n250 & n319 );
  assign n321 = ~n250 & n319 ;
  assign n322 = ( n163 & n320 ) | ( n163 & n321 ) | ( n320 & n321 );
  assign n323 = n316 & ~n322 ;
  assign n324 = n136 & n323 ;
  assign n325 = ~G5 & n136 ;
  assign n326 = n323 & n325 ;
  assign n327 = G5 | n325 ;
  assign n328 = ( G5 & n323 ) | ( G5 & n327 ) | ( n323 & n327 );
  assign n329 = ( ~n324 & n326 ) | ( ~n324 & n328 ) | ( n326 & n328 );
  assign n330 = n159 & n323 ;
  assign n331 = ~G6 & n159 ;
  assign n332 = n323 & n331 ;
  assign n333 = G6 | n331 ;
  assign n334 = ( G6 & n323 ) | ( G6 & n333 ) | ( n323 & n333 );
  assign n335 = ( ~n330 & n332 ) | ( ~n330 & n334 ) | ( n332 & n334 );
  assign n336 = n111 & n323 ;
  assign n337 = ~G7 & n111 ;
  assign n338 = n323 & n337 ;
  assign n339 = G7 | n337 ;
  assign n340 = ( G7 & n323 ) | ( G7 & n339 ) | ( n323 & n339 );
  assign n341 = ( ~n336 & n338 ) | ( ~n336 & n340 ) | ( n338 & n340 );
  assign n342 = n111 & n275 ;
  assign n343 = ~n76 & n284 ;
  assign n344 = ( ~n76 & n291 ) | ( ~n76 & n343 ) | ( n291 & n343 );
  assign n345 = n342 & n344 ;
  assign n346 = n196 & n345 ;
  assign n347 = G20 & n345 ;
  assign n348 = n196 & n347 ;
  assign n349 = G20 & ~n347 ;
  assign n350 = ( G20 & ~n196 ) | ( G20 & n349 ) | ( ~n196 & n349 );
  assign n351 = ( n346 & ~n348 ) | ( n346 & n350 ) | ( ~n348 & n350 );
  assign n352 = n76 & n323 ;
  assign n353 = ~G8 & n76 ;
  assign n354 = n323 & n353 ;
  assign n355 = G8 | n353 ;
  assign n356 = ( G8 & n323 ) | ( G8 & n355 ) | ( n323 & n355 );
  assign n357 = ( ~n352 & n354 ) | ( ~n352 & n356 ) | ( n354 & n356 );
  assign n358 = n268 & n289 ;
  assign n359 = ~n249 & n268 ;
  assign n360 = ( n222 & n358 ) | ( n222 & n359 ) | ( n358 & n359 );
  assign n361 = n197 & n360 ;
  assign n362 = n163 & n361 ;
  assign n363 = G9 & ~n362 ;
  assign n364 = ~G9 & n362 ;
  assign n365 = n363 | n364 ;
  assign n366 = n159 & n360 ;
  assign n367 = n300 & n366 ;
  assign n368 = ~G10 & n366 ;
  assign n369 = n300 & n368 ;
  assign n370 = G10 | n369 ;
  assign n371 = ( ~n367 & n369 ) | ( ~n367 & n370 ) | ( n369 & n370 );
  assign n372 = n111 & n360 ;
  assign n373 = n300 & n372 ;
  assign n374 = ~G11 & n372 ;
  assign n375 = n300 & n374 ;
  assign n376 = G11 | n375 ;
  assign n377 = ( ~n373 & n375 ) | ( ~n373 & n376 ) | ( n375 & n376 );
  assign n378 = n76 & n360 ;
  assign n379 = n300 & n378 ;
  assign n380 = ~G12 & n378 ;
  assign n381 = n300 & n380 ;
  assign n382 = G12 | n381 ;
  assign n383 = ( ~n379 & n381 ) | ( ~n379 & n382 ) | ( n381 & n382 );
  assign n384 = ~n268 & n289 ;
  assign n385 = n249 | n268 ;
  assign n386 = ( n222 & n384 ) | ( n222 & ~n385 ) | ( n384 & ~n385 );
  assign n387 = n136 & n386 ;
  assign n388 = n316 & n387 ;
  assign n389 = ~G13 & n387 ;
  assign n390 = n316 & n389 ;
  assign n391 = G13 | n390 ;
  assign n392 = ( ~n388 & n390 ) | ( ~n388 & n391 ) | ( n390 & n391 );
  assign n393 = n159 & n386 ;
  assign n394 = n316 & n393 ;
  assign n395 = ~G14 & n393 ;
  assign n396 = n316 & n395 ;
  assign n397 = G14 | n396 ;
  assign n398 = ( ~n394 & n396 ) | ( ~n394 & n397 ) | ( n396 & n397 );
  assign n399 = n111 & n386 ;
  assign n400 = n316 & n399 ;
  assign n401 = ~G15 & n399 ;
  assign n402 = n316 & n401 ;
  assign n403 = G15 | n402 ;
  assign n404 = ( ~n400 & n402 ) | ( ~n400 & n403 ) | ( n402 & n403 );
  assign n405 = n76 & n386 ;
  assign n406 = n316 & n405 ;
  assign n407 = ~G16 & n405 ;
  assign n408 = n316 & n407 ;
  assign n409 = G16 | n408 ;
  assign n410 = ( ~n406 & n408 ) | ( ~n406 & n409 ) | ( n408 & n409 );
  assign n411 = n249 & n345 ;
  assign n412 = G17 & ~n411 ;
  assign n413 = ~G17 & n411 ;
  assign n414 = n412 | n413 ;
  assign n415 = n222 | n226 ;
  assign n416 = n345 & n415 ;
  assign n417 = G18 & n416 ;
  assign n418 = G18 & ~n417 ;
  assign n419 = ( n416 & ~n417 ) | ( n416 & n418 ) | ( ~n417 & n418 );
  assign n420 = n268 & n345 ;
  assign n421 = G19 & n345 ;
  assign n422 = n268 & n421 ;
  assign n423 = G19 & ~n421 ;
  assign n424 = ( G19 & ~n268 ) | ( G19 & n423 ) | ( ~n268 & n423 );
  assign n425 = ( n420 & ~n422 ) | ( n420 & n424 ) | ( ~n422 & n424 );
  assign n426 = n293 & n415 ;
  assign n427 = G22 & n426 ;
  assign n428 = G22 & ~n427 ;
  assign n429 = ( n426 & ~n427 ) | ( n426 & n428 ) | ( ~n427 & n428 );
  assign n430 = n268 & n293 ;
  assign n431 = G23 & n293 ;
  assign n432 = n268 & n431 ;
  assign n433 = G23 & ~n431 ;
  assign n434 = ( G23 & ~n268 ) | ( G23 & n433 ) | ( ~n268 & n433 );
  assign n435 = ( n430 & ~n432 ) | ( n430 & n434 ) | ( ~n432 & n434 );
  assign n436 = n196 & n293 ;
  assign n437 = G24 & n293 ;
  assign n438 = n196 & n437 ;
  assign n439 = G24 & ~n437 ;
  assign n440 = ( G24 & ~n196 ) | ( G24 & n439 ) | ( ~n196 & n439 );
  assign n441 = ( n436 & ~n438 ) | ( n436 & n440 ) | ( ~n438 & n440 );
  assign n442 = ~n136 & n159 ;
  assign n443 = n111 & n442 ;
  assign n444 = n344 & n443 ;
  assign n445 = n249 & n444 ;
  assign n446 = G25 & n444 ;
  assign n447 = n249 & n446 ;
  assign n448 = G25 & ~n446 ;
  assign n449 = ( G25 & ~n249 ) | ( G25 & n448 ) | ( ~n249 & n448 );
  assign n450 = ( n445 & ~n447 ) | ( n445 & n449 ) | ( ~n447 & n449 );
  assign n451 = n415 & n444 ;
  assign n452 = G26 & n451 ;
  assign n453 = G26 & ~n452 ;
  assign n454 = ( n451 & ~n452 ) | ( n451 & n453 ) | ( ~n452 & n453 );
  assign n455 = n268 & n444 ;
  assign n456 = G27 & n444 ;
  assign n457 = n268 & n456 ;
  assign n458 = G27 & ~n456 ;
  assign n459 = ( G27 & ~n268 ) | ( G27 & n458 ) | ( ~n268 & n458 );
  assign n460 = ( n455 & ~n457 ) | ( n455 & n459 ) | ( ~n457 & n459 );
  assign n461 = n196 & n444 ;
  assign n462 = G28 & n444 ;
  assign n463 = n196 & n462 ;
  assign n464 = G28 & ~n462 ;
  assign n465 = ( G28 & ~n196 ) | ( G28 & n464 ) | ( ~n196 & n464 );
  assign n466 = ( n461 & ~n463 ) | ( n461 & n465 ) | ( ~n463 & n465 );
  assign n467 = n76 & n292 ;
  assign n468 = ~n111 & n442 ;
  assign n469 = n467 & n468 ;
  assign n470 = n249 & n469 ;
  assign n471 = G29 & n469 ;
  assign n472 = n249 & n471 ;
  assign n473 = G29 & ~n471 ;
  assign n474 = ( G29 & ~n249 ) | ( G29 & n473 ) | ( ~n249 & n473 );
  assign n475 = ( n470 & ~n472 ) | ( n470 & n474 ) | ( ~n472 & n474 );
  assign n476 = n415 & n469 ;
  assign n477 = G30 & n476 ;
  assign n478 = G30 & ~n477 ;
  assign n479 = ( n476 & ~n477 ) | ( n476 & n478 ) | ( ~n477 & n478 );
  assign n480 = n268 & n469 ;
  assign n481 = G31 & n469 ;
  assign n482 = n268 & n481 ;
  assign n483 = G31 & ~n481 ;
  assign n484 = ( G31 & ~n268 ) | ( G31 & n483 ) | ( ~n268 & n483 );
  assign n485 = ( n480 & ~n482 ) | ( n480 & n484 ) | ( ~n482 & n484 );
  assign n486 = n196 & n469 ;
  assign n487 = G32 & n469 ;
  assign n488 = n196 & n487 ;
  assign n489 = G32 & ~n487 ;
  assign n490 = ( G32 & ~n196 ) | ( G32 & n489 ) | ( ~n196 & n489 );
  assign n491 = ( n486 & ~n488 ) | ( n486 & n490 ) | ( ~n488 & n490 );
  assign G1324 = ~n274 ;
  assign G1344 = ~n299 ;
  assign G1325 = ~n305 ;
  assign G1326 = ~n310 ;
  assign G1327 = ~n315 ;
  assign G1328 = ~n329 ;
  assign G1329 = ~n335 ;
  assign G1330 = ~n341 ;
  assign G1343 = ~n351 ;
  assign G1331 = ~n357 ;
  assign G1332 = ~n365 ;
  assign G1333 = ~n371 ;
  assign G1334 = ~n377 ;
  assign G1335 = ~n383 ;
  assign G1336 = ~n392 ;
  assign G1337 = ~n398 ;
  assign G1338 = ~n404 ;
  assign G1339 = ~n410 ;
  assign G1340 = ~n414 ;
  assign G1341 = ~n419 ;
  assign G1342 = ~n425 ;
  assign G1345 = ~n429 ;
  assign G1346 = ~n435 ;
  assign G1347 = ~n441 ;
  assign G1348 = ~n450 ;
  assign G1349 = ~n454 ;
  assign G1350 = ~n460 ;
  assign G1351 = ~n466 ;
  assign G1352 = ~n475 ;
  assign G1353 = ~n479 ;
  assign G1354 = ~n485 ;
  assign G1355 = ~n491 ;
endmodule
