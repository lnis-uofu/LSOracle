module top(pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 , pi8 , pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 , pi16 , pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 , po0 , po1 , po2 , po3 , po4 , po5 , po6 , po7 , po8 , po9 , po10 , po11 , po12 , po13 , po14 , po15 , po16 , po17 , po18 , po19 , po20 , po21 , po22 , po23 , po24 );
  input pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 , pi8 , pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 , pi16 , pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 ;
  output po0 , po1 , po2 , po3 , po4 , po5 , po6 , po7 , po8 , po9 , po10 , po11 , po12 , po13 , po14 , po15 , po16 , po17 , po18 , po19 , po20 , po21 , po22 , po23 , po24 ;
  wire n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500;
  assign n25 = pi2 & pi22 ;
  assign n26 = pi0 & ~pi22 ;
  assign n27 = pi1 | pi2 ;
  assign n28 = ( ~pi22 & n26 ) | ( ~pi22 & n27 ) | ( n26 & n27 );
  assign n29 = pi0 | pi1 ;
  assign n30 = pi2 & n29 ;
  assign n31 = n28 & ~n30 ;
  assign n32 = n25 | n31 ;
  assign n33 = pi5 | pi8 ;
  assign n34 = pi7 | pi10 ;
  assign n35 = pi4 | pi6 ;
  assign n36 = n34 | n35 ;
  assign n37 = n33 | n36 ;
  assign n38 = pi0 | n27 ;
  assign n39 = pi3 | n38 ;
  assign n40 = pi9 | n39 ;
  assign n41 = pi11 | pi12 ;
  assign n42 = n40 | n41 ;
  assign n43 = n37 | n42 ;
  assign n44 = ~pi22 & n43 ;
  assign n45 = pi13 & ~n44 ;
  assign n46 = ~pi13 & n44 ;
  assign n47 = n45 | n46 ;
  assign n48 = pi13 | n43 ;
  assign n49 = pi14 | n48 ;
  assign n50 = ~pi22 & n49 ;
  assign n51 = ~pi15 & n50 ;
  assign n52 = pi15 & ~n50 ;
  assign n53 = n51 | n52 ;
  assign n54 = pi17 | n49 ;
  assign n55 = pi16 | n54 ;
  assign n56 = pi15 | pi18 ;
  assign n57 = pi19 | n56 ;
  assign n58 = n55 | n57 ;
  assign n59 = ~pi22 & n58 ;
  assign n60 = ~pi20 & n59 ;
  assign n61 = pi20 & ~n59 ;
  assign n62 = n60 | n61 ;
  assign n63 = pi16 | pi20 ;
  assign n64 = n54 | n63 ;
  assign n65 = n57 | n64 ;
  assign n66 = ~pi22 & n65 ;
  assign n67 = ~pi21 & n66 ;
  assign n68 = pi21 & ~n66 ;
  assign n69 = n67 | n68 ;
  assign n70 = n62 & n69 ;
  assign n71 = n53 & n70 ;
  assign n72 = ~n53 & n70 ;
  assign n73 = n71 | n72 ;
  assign n74 = pi16 | n49 ;
  assign n75 = pi15 | pi17 ;
  assign n76 = n74 | n75 ;
  assign n77 = ~pi22 & n76 ;
  assign n78 = ~pi18 & n77 ;
  assign n79 = pi18 & ~n77 ;
  assign n80 = n78 | n79 ;
  assign n81 = pi18 | n76 ;
  assign n82 = ~pi22 & n81 ;
  assign n83 = pi19 & ~n82 ;
  assign n84 = pi19 | pi22 ;
  assign n85 = n81 & ~n84 ;
  assign n86 = n83 | n85 ;
  assign n87 = n80 & n86 ;
  assign n88 = pi15 | n49 ;
  assign n89 = ~pi22 & n88 ;
  assign n90 = pi16 & ~n89 ;
  assign n91 = ~pi16 & n89 ;
  assign n92 = n90 | n91 ;
  assign n93 = pi16 | n88 ;
  assign n94 = ~pi22 & n93 ;
  assign n95 = pi17 & ~n94 ;
  assign n96 = ~pi17 & n94 ;
  assign n97 = n95 | n96 ;
  assign n98 = n92 & n97 ;
  assign n99 = n87 & n98 ;
  assign n100 = ~n92 & n97 ;
  assign n101 = n80 | n86 ;
  assign n102 = n100 & ~n101 ;
  assign n103 = n99 | n102 ;
  assign n104 = n73 & n103 ;
  assign n105 = n87 & n100 ;
  assign n106 = n72 & n105 ;
  assign n107 = n80 & ~n86 ;
  assign n108 = n98 & n107 ;
  assign n109 = n71 & n108 ;
  assign n110 = n92 | n97 ;
  assign n111 = ~n80 & n86 ;
  assign n112 = ~n110 & n111 ;
  assign n113 = ~n62 & n69 ;
  assign n114 = ~n53 & n113 ;
  assign n115 = n112 & n114 ;
  assign n116 = n53 & n113 ;
  assign n117 = n112 & n116 ;
  assign n118 = n115 | n117 ;
  assign n119 = n109 | n118 ;
  assign n120 = n107 & ~n110 ;
  assign n121 = n71 & n120 ;
  assign n122 = n72 & n108 ;
  assign n123 = n100 & n107 ;
  assign n124 = n71 & n123 ;
  assign n125 = n122 | n124 ;
  assign n126 = n92 & ~n97 ;
  assign n127 = n111 & n126 ;
  assign n128 = n114 & n127 ;
  assign n129 = n72 & n120 ;
  assign n130 = n128 | n129 ;
  assign n131 = n125 | n130 ;
  assign n132 = n121 | n131 ;
  assign n133 = n119 | n132 ;
  assign n134 = n106 | n133 ;
  assign n135 = n99 & n116 ;
  assign n136 = n101 | n110 ;
  assign n137 = n72 & ~n136 ;
  assign n138 = n135 | n137 ;
  assign n139 = n98 & ~n101 ;
  assign n140 = n71 & n139 ;
  assign n141 = n87 & n126 ;
  assign n142 = n116 & n141 ;
  assign n143 = n140 | n142 ;
  assign n144 = n100 & n111 ;
  assign n145 = n71 & n144 ;
  assign n146 = n72 & n144 ;
  assign n147 = n98 & n111 ;
  assign n148 = n72 & n147 ;
  assign n149 = n146 | n148 ;
  assign n150 = n87 & ~n110 ;
  assign n151 = n116 & n150 ;
  assign n152 = n72 & n139 ;
  assign n153 = n151 | n152 ;
  assign n154 = n149 | n153 ;
  assign n155 = n145 | n154 ;
  assign n156 = n143 | n155 ;
  assign n157 = n114 & n150 ;
  assign n158 = n114 & n141 ;
  assign n159 = n157 | n158 ;
  assign n160 = n156 | n159 ;
  assign n161 = n138 | n160 ;
  assign n162 = n134 | n161 ;
  assign n163 = n72 & n141 ;
  assign n164 = n116 & n127 ;
  assign n165 = n71 & n127 ;
  assign n166 = n164 | n165 ;
  assign n167 = n71 & ~n136 ;
  assign n168 = n71 & n141 ;
  assign n169 = ~n101 & n126 ;
  assign n170 = n72 & n169 ;
  assign n171 = n168 | n170 ;
  assign n172 = n167 | n171 ;
  assign n173 = n166 | n172 ;
  assign n174 = n163 | n173 ;
  assign n175 = n162 | n174 ;
  assign n176 = n71 & n105 ;
  assign n177 = n71 & n169 ;
  assign n178 = n176 | n177 ;
  assign n179 = n71 & n147 ;
  assign n180 = n105 & n116 ;
  assign n181 = n72 & n150 ;
  assign n182 = n180 | n181 ;
  assign n183 = n179 | n182 ;
  assign n184 = n99 & n114 ;
  assign n185 = n71 & n150 ;
  assign n186 = n105 & n114 ;
  assign n187 = n185 | n186 ;
  assign n188 = n184 | n187 ;
  assign n189 = n183 | n188 ;
  assign n190 = n116 & n147 ;
  assign n191 = n116 & n144 ;
  assign n192 = n114 & n144 ;
  assign n193 = n191 | n192 ;
  assign n194 = n71 & n112 ;
  assign n195 = n114 & n147 ;
  assign n196 = n72 & n112 ;
  assign n197 = n195 | n196 ;
  assign n198 = n194 | n197 ;
  assign n199 = n193 | n198 ;
  assign n200 = n116 & n123 ;
  assign n201 = n108 & n114 ;
  assign n202 = n200 | n201 ;
  assign n203 = n107 & n126 ;
  assign n204 = n71 & n203 ;
  assign n205 = n108 & n116 ;
  assign n206 = n204 | n205 ;
  assign n207 = n72 & n203 ;
  assign n208 = n72 & n127 ;
  assign n209 = n72 & n123 ;
  assign n210 = n208 | n209 ;
  assign n211 = n207 | n210 ;
  assign n212 = n206 | n211 ;
  assign n213 = n202 | n212 ;
  assign n214 = n199 | n213 ;
  assign n215 = n190 | n214 ;
  assign n216 = n189 | n215 ;
  assign n217 = n178 | n216 ;
  assign n218 = n175 | n217 ;
  assign n219 = n104 | n218 ;
  assign n220 = n47 & n219 ;
  assign n221 = ~pi22 & n48 ;
  assign n222 = ~pi14 & n221 ;
  assign n223 = pi14 & ~n221 ;
  assign n224 = n222 | n223 ;
  assign n225 = n62 | n69 ;
  assign n226 = n53 & ~n225 ;
  assign n227 = n127 & n226 ;
  assign n228 = n53 | n225 ;
  assign n229 = n147 & ~n228 ;
  assign n230 = n144 & n226 ;
  assign n231 = n229 | n230 ;
  assign n232 = n144 & ~n228 ;
  assign n233 = n147 & n226 ;
  assign n234 = n127 & ~n228 ;
  assign n235 = n233 | n234 ;
  assign n236 = n232 | n235 ;
  assign n237 = n231 | n236 ;
  assign n238 = n150 & ~n228 ;
  assign n239 = n99 & n226 ;
  assign n240 = n105 & n226 ;
  assign n241 = n62 & ~n69 ;
  assign n242 = ~n53 & n241 ;
  assign n243 = ~n136 & n242 ;
  assign n244 = n240 | n243 ;
  assign n245 = n53 & n241 ;
  assign n246 = ~n136 & n245 ;
  assign n247 = n116 & n120 ;
  assign n248 = n116 & n203 ;
  assign n249 = n247 | n248 ;
  assign n250 = n246 | n249 ;
  assign n251 = n150 & n226 ;
  assign n252 = n141 & n226 ;
  assign n253 = n251 | n252 ;
  assign n254 = n250 | n253 ;
  assign n255 = n105 & ~n228 ;
  assign n256 = n114 & n120 ;
  assign n257 = n114 & n203 ;
  assign n258 = n256 | n257 ;
  assign n259 = n255 | n258 ;
  assign n260 = n254 | n259 ;
  assign n261 = n244 | n260 ;
  assign n262 = n239 | n261 ;
  assign n263 = n99 & ~n228 ;
  assign n264 = n141 & ~n228 ;
  assign n265 = n263 | n264 ;
  assign n266 = n262 | n265 ;
  assign n267 = n238 | n266 ;
  assign n268 = n112 & n226 ;
  assign n269 = n150 & n242 ;
  assign n270 = n147 & n245 ;
  assign n271 = n147 & n242 ;
  assign n272 = n270 | n271 ;
  assign n273 = n105 & n245 ;
  assign n274 = n141 & n242 ;
  assign n275 = n150 & n245 ;
  assign n276 = n141 & n245 ;
  assign n277 = n275 | n276 ;
  assign n278 = n274 | n277 ;
  assign n279 = n273 | n278 ;
  assign n280 = n272 | n279 ;
  assign n281 = n144 & n245 ;
  assign n282 = n114 & n169 ;
  assign n283 = n281 | n282 ;
  assign n284 = n99 & n245 ;
  assign n285 = n105 & n242 ;
  assign n286 = n114 & n139 ;
  assign n287 = n285 | n286 ;
  assign n288 = n284 | n287 ;
  assign n289 = n283 | n288 ;
  assign n290 = n102 & n116 ;
  assign n291 = n116 & n169 ;
  assign n292 = n290 | n291 ;
  assign n293 = n99 & n242 ;
  assign n294 = n114 & n123 ;
  assign n295 = n293 | n294 ;
  assign n296 = n102 & n114 ;
  assign n297 = n116 & n139 ;
  assign n298 = n296 | n297 ;
  assign n299 = n295 | n298 ;
  assign n300 = n292 | n299 ;
  assign n301 = n289 | n300 ;
  assign n302 = n280 | n301 ;
  assign n303 = n269 | n302 ;
  assign n304 = n114 & ~n136 ;
  assign n305 = n116 & ~n136 ;
  assign n306 = n304 | n305 ;
  assign n307 = n303 | n306 ;
  assign n308 = n268 | n307 ;
  assign n309 = n267 | n308 ;
  assign n310 = n237 | n309 ;
  assign n311 = n227 | n310 ;
  assign n312 = n203 & n242 ;
  assign n313 = n139 & n245 ;
  assign n314 = n120 & n242 ;
  assign n315 = n313 | n314 ;
  assign n316 = n102 & n245 ;
  assign n317 = n169 & n245 ;
  assign n318 = n102 & n242 ;
  assign n319 = n139 & n242 ;
  assign n320 = n120 & n245 ;
  assign n321 = n169 & n242 ;
  assign n322 = n320 | n321 ;
  assign n323 = n319 | n322 ;
  assign n324 = n318 | n323 ;
  assign n325 = n317 | n324 ;
  assign n326 = n316 | n325 ;
  assign n327 = n315 | n326 ;
  assign n328 = n112 & n245 ;
  assign n329 = n203 & n245 ;
  assign n330 = n108 & n242 ;
  assign n331 = n123 & n242 ;
  assign n332 = n330 | n331 ;
  assign n333 = n329 | n332 ;
  assign n334 = n123 & n245 ;
  assign n335 = n108 & n245 ;
  assign n336 = n144 & n242 ;
  assign n337 = n335 | n336 ;
  assign n338 = n334 | n337 ;
  assign n339 = n333 | n338 ;
  assign n340 = n328 | n339 ;
  assign n341 = n127 & n245 ;
  assign n342 = n112 & n242 ;
  assign n343 = n127 & n242 ;
  assign n344 = n342 | n343 ;
  assign n345 = n341 | n344 ;
  assign n346 = n340 | n345 ;
  assign n347 = n249 | n346 ;
  assign n348 = n307 | n347 ;
  assign n349 = n258 | n348 ;
  assign n350 = n327 | n349 ;
  assign n351 = n312 | n350 ;
  assign n352 = n311 & n351 ;
  assign n353 = n219 & ~n352 ;
  assign n354 = n224 | n353 ;
  assign n355 = ~n311 & n351 ;
  assign n356 = n311 & ~n351 ;
  assign n357 = n355 | n356 ;
  assign n358 = ~n353 & n357 ;
  assign n359 = n311 | n351 ;
  assign n360 = ~n219 & n359 ;
  assign n361 = n357 | n360 ;
  assign n362 = n224 & ~n361 ;
  assign n363 = n358 | n362 ;
  assign n364 = n354 & ~n363 ;
  assign n365 = ~n220 & n364 ;
  assign n366 = pi8 | pi10 ;
  assign n367 = pi4 | pi5 ;
  assign n368 = n366 | n367 ;
  assign n369 = pi6 | pi7 ;
  assign n370 = n40 | n369 ;
  assign n371 = n368 | n370 ;
  assign n372 = ~pi22 & n371 ;
  assign n373 = pi11 & ~n372 ;
  assign n374 = ~pi11 & n372 ;
  assign n375 = n373 | n374 ;
  assign n376 = n219 & n375 ;
  assign n377 = n108 & ~n228 ;
  assign n378 = n297 | n329 ;
  assign n379 = n377 | n378 ;
  assign n380 = n181 | n256 ;
  assign n381 = n264 | n304 ;
  assign n382 = n203 & n226 ;
  assign n383 = n120 & ~n228 ;
  assign n384 = n305 | n383 ;
  assign n385 = n247 | n384 ;
  assign n386 = n167 | n207 ;
  assign n387 = n109 | n341 ;
  assign n388 = n386 | n387 ;
  assign n389 = n123 & ~n228 ;
  assign n390 = n328 | n389 ;
  assign n391 = n246 | n331 ;
  assign n392 = n120 & n226 ;
  assign n393 = n255 | n392 ;
  assign n394 = n210 | n393 ;
  assign n395 = n124 | n165 ;
  assign n396 = n394 | n395 ;
  assign n397 = n391 | n396 ;
  assign n398 = n390 | n397 ;
  assign n399 = n71 & n99 ;
  assign n400 = n112 & ~n228 ;
  assign n401 = n203 & ~n228 ;
  assign n402 = n149 | n337 ;
  assign n403 = n108 & n226 ;
  assign n404 = n244 | n257 ;
  assign n405 = n71 & n102 ;
  assign n406 = n121 | n405 ;
  assign n407 = n179 | n406 ;
  assign n408 = n404 | n407 ;
  assign n409 = n403 | n408 ;
  assign n410 = n294 | n409 ;
  assign n411 = n402 | n410 ;
  assign n412 = n248 | n411 ;
  assign n413 = n106 | n152 ;
  assign n414 = n129 | n413 ;
  assign n415 = n178 | n330 ;
  assign n416 = n414 | n415 ;
  assign n417 = n412 | n416 ;
  assign n418 = n401 | n417 ;
  assign n419 = n400 | n418 ;
  assign n420 = n399 | n419 ;
  assign n421 = n398 | n420 ;
  assign n422 = n251 | n286 ;
  assign n423 = n196 | n342 ;
  assign n424 = n170 | n423 ;
  assign n425 = n422 | n424 ;
  assign n426 = n421 | n425 ;
  assign n427 = n388 | n426 ;
  assign n428 = n385 | n427 ;
  assign n429 = n382 | n428 ;
  assign n430 = n381 | n429 ;
  assign n431 = n380 | n430 ;
  assign n432 = n185 | n290 ;
  assign n433 = n72 & n99 ;
  assign n434 = n137 | n184 ;
  assign n435 = n168 | n343 ;
  assign n436 = n434 | n435 ;
  assign n437 = n433 | n436 ;
  assign n438 = n334 | n437 ;
  assign n439 = n432 | n438 ;
  assign n440 = n140 | n291 ;
  assign n441 = n122 | n194 ;
  assign n442 = n252 | n441 ;
  assign n443 = n440 | n442 ;
  assign n444 = n135 | n282 ;
  assign n445 = n163 | n444 ;
  assign n446 = n239 | n445 ;
  assign n447 = n123 & n226 ;
  assign n448 = n72 & n102 ;
  assign n449 = n145 | n296 ;
  assign n450 = n448 | n449 ;
  assign n451 = n447 | n450 ;
  assign n452 = n204 | n451 ;
  assign n453 = n446 | n452 ;
  assign n454 = n443 | n453 ;
  assign n455 = n439 | n454 ;
  assign n456 = n431 | n455 ;
  assign n457 = n379 | n456 ;
  assign n458 = n263 | n457 ;
  assign n459 = n186 | n248 ;
  assign n460 = n191 | n400 ;
  assign n461 = n336 | n460 ;
  assign n462 = n459 | n461 ;
  assign n463 = n257 | n286 ;
  assign n464 = n157 | n276 ;
  assign n465 = n463 | n464 ;
  assign n466 = n273 | n312 ;
  assign n467 = n165 | n466 ;
  assign n468 = n210 | n447 ;
  assign n469 = n467 | n468 ;
  assign n470 = n149 | n163 ;
  assign n471 = n122 | n176 ;
  assign n472 = n470 | n471 ;
  assign n473 = n180 | n285 ;
  assign n474 = n109 | n403 ;
  assign n475 = n473 | n474 ;
  assign n476 = n472 | n475 ;
  assign n477 = n469 | n476 ;
  assign n478 = n314 | n477 ;
  assign n479 = n194 | n478 ;
  assign n480 = n293 | n328 ;
  assign n481 = n243 | n480 ;
  assign n482 = n479 | n481 ;
  assign n483 = n139 & ~n228 ;
  assign n484 = n151 | n483 ;
  assign n485 = n482 | n484 ;
  assign n486 = n320 | n433 ;
  assign n487 = n344 | n486 ;
  assign n488 = n230 | n487 ;
  assign n489 = n284 | n297 ;
  assign n490 = n124 | n190 ;
  assign n491 = n247 | n490 ;
  assign n492 = n196 | n491 ;
  assign n493 = n238 | n492 ;
  assign n494 = n489 | n493 ;
  assign n495 = n488 | n494 ;
  assign n496 = n485 | n495 ;
  assign n497 = n465 | n496 ;
  assign n498 = n462 | n497 ;
  assign n499 = n102 & ~n228 ;
  assign n500 = n142 | n233 ;
  assign n501 = n158 | n500 ;
  assign n502 = n204 | n263 ;
  assign n503 = n102 & n226 ;
  assign n504 = n389 | n503 ;
  assign n505 = n207 | n504 ;
  assign n506 = n502 | n505 ;
  assign n507 = n246 | n341 ;
  assign n508 = n168 | n185 ;
  assign n509 = n195 | n508 ;
  assign n510 = n380 | n509 ;
  assign n511 = n229 | n510 ;
  assign n512 = n507 | n511 ;
  assign n513 = n139 & n226 ;
  assign n514 = n239 | n313 ;
  assign n515 = n513 | n514 ;
  assign n516 = n145 | n399 ;
  assign n517 = n179 | n516 ;
  assign n518 = n515 | n517 ;
  assign n519 = n512 | n518 ;
  assign n520 = n506 | n519 ;
  assign n521 = n501 | n520 ;
  assign n522 = n499 | n521 ;
  assign n523 = n106 | n294 ;
  assign n524 = n522 | n523 ;
  assign n525 = n377 | n524 ;
  assign n526 = n498 | n525 ;
  assign n527 = n458 & n526 ;
  assign n528 = n311 & ~n527 ;
  assign n529 = n376 & ~n528 ;
  assign n530 = ~n376 & n528 ;
  assign n531 = n529 | n530 ;
  assign n532 = pi11 & ~pi22 ;
  assign n533 = n372 | n532 ;
  assign n534 = pi12 & n533 ;
  assign n535 = pi12 | n532 ;
  assign n536 = n372 | n535 ;
  assign n537 = ~n534 & n536 ;
  assign n538 = n219 & n537 ;
  assign n539 = ~n531 & n538 ;
  assign n540 = n529 | n539 ;
  assign n541 = n220 & ~n364 ;
  assign n542 = n365 | n541 ;
  assign n543 = n540 & ~n542 ;
  assign n544 = n365 | n543 ;
  assign n545 = n458 | n526 ;
  assign n546 = ~n311 & n545 ;
  assign n547 = n458 & ~n526 ;
  assign n548 = ~n458 & n526 ;
  assign n549 = n547 | n548 ;
  assign n550 = n546 | n549 ;
  assign n551 = n224 & ~n550 ;
  assign n552 = n528 | n549 ;
  assign n553 = n224 & ~n552 ;
  assign n554 = ( n528 & ~n551 ) | ( n528 & n553 ) | ( ~n551 & n553 );
  assign n555 = ~n376 & n554 ;
  assign n556 = n376 & ~n554 ;
  assign n557 = n555 | n556 ;
  assign n558 = n353 | n357 ;
  assign n559 = n537 | n558 ;
  assign n560 = ~n361 & n536 ;
  assign n561 = ~n534 & n560 ;
  assign n562 = n559 & ~n561 ;
  assign n563 = n357 & ~n360 ;
  assign n564 = n47 & n563 ;
  assign n565 = ~n47 & n358 ;
  assign n566 = n564 | n565 ;
  assign n567 = n562 & ~n566 ;
  assign n568 = ~n557 & n567 ;
  assign n569 = n555 | n568 ;
  assign n570 = n224 & n563 ;
  assign n571 = ~n223 & n358 ;
  assign n572 = ~n222 & n571 ;
  assign n573 = n47 & ~n361 ;
  assign n574 = n47 | n558 ;
  assign n575 = ~n573 & n574 ;
  assign n576 = ~n572 & n575 ;
  assign n577 = ~n570 & n576 ;
  assign n578 = n569 & n577 ;
  assign n579 = n569 | n577 ;
  assign n580 = ~n578 & n579 ;
  assign n581 = n531 & ~n538 ;
  assign n582 = n539 | n581 ;
  assign n583 = n580 & ~n582 ;
  assign n584 = n578 | n583 ;
  assign n585 = ~n540 & n542 ;
  assign n586 = n543 | n585 ;
  assign n587 = n584 & ~n586 ;
  assign n588 = n169 & n226 ;
  assign n589 = n233 | n588 ;
  assign n590 = n145 | n181 ;
  assign n591 = n168 | n238 ;
  assign n592 = n269 | n591 ;
  assign n593 = n590 | n592 ;
  assign n594 = n140 | n255 ;
  assign n595 = n151 | n594 ;
  assign n596 = n165 | n595 ;
  assign n597 = n593 | n596 ;
  assign n598 = n227 | n341 ;
  assign n599 = n158 | n598 ;
  assign n600 = n448 | n599 ;
  assign n601 = n284 | n293 ;
  assign n602 = n192 | n601 ;
  assign n603 = n296 | n602 ;
  assign n604 = n600 | n603 ;
  assign n605 = n597 | n604 ;
  assign n606 = n180 | n319 ;
  assign n607 = n605 | n606 ;
  assign n608 = n164 | n185 ;
  assign n609 = n607 | n608 ;
  assign n610 = n318 | n320 ;
  assign n611 = n433 | n610 ;
  assign n612 = n609 | n611 ;
  assign n613 = n274 | n513 ;
  assign n614 = n186 | n613 ;
  assign n615 = n252 | n614 ;
  assign n616 = n246 | n615 ;
  assign n617 = n117 | n163 ;
  assign n618 = n128 | n142 ;
  assign n619 = n617 | n618 ;
  assign n620 = n232 | n466 ;
  assign n621 = n290 | n382 ;
  assign n622 = n169 & ~n228 ;
  assign n623 = n291 | n483 ;
  assign n624 = n622 | n623 ;
  assign n625 = n621 | n624 ;
  assign n626 = n620 | n625 ;
  assign n627 = n316 | n626 ;
  assign n628 = n275 | n627 ;
  assign n629 = n420 | n628 ;
  assign n630 = n619 | n629 ;
  assign n631 = n616 | n630 ;
  assign n632 = n612 | n631 ;
  assign n633 = n589 | n632 ;
  assign n634 = n208 | n275 ;
  assign n635 = n335 | n634 ;
  assign n636 = n164 | n588 ;
  assign n637 = n190 | n636 ;
  assign n638 = n336 | n637 ;
  assign n639 = n250 | n638 ;
  assign n640 = n255 | n639 ;
  assign n641 = n240 | n640 ;
  assign n642 = n635 | n641 ;
  assign n643 = n196 | n317 ;
  assign n644 = n331 | n343 ;
  assign n645 = n643 | n644 ;
  assign n646 = n400 | n645 ;
  assign n647 = n316 | n503 ;
  assign n648 = n646 | n647 ;
  assign n649 = n642 | n648 ;
  assign n650 = n186 | n649 ;
  assign n651 = n142 | n290 ;
  assign n652 = n282 | n651 ;
  assign n653 = n650 | n652 ;
  assign n654 = ~n136 & n226 ;
  assign n655 = n140 | n314 ;
  assign n656 = n274 | n655 ;
  assign n657 = n137 | n170 ;
  assign n658 = n656 | n657 ;
  assign n659 = n232 | n658 ;
  assign n660 = n654 | n659 ;
  assign n661 = n238 | n660 ;
  assign n662 = n129 | n661 ;
  assign n663 = n264 | n284 ;
  assign n664 = n234 | n663 ;
  assign n665 = n312 | n328 ;
  assign n666 = n115 | n192 ;
  assign n667 = n665 | n666 ;
  assign n668 = n664 | n667 ;
  assign n669 = n377 | n668 ;
  assign n670 = n662 | n669 ;
  assign n671 = n382 | n392 ;
  assign n672 = n256 | n671 ;
  assign n673 = n152 | n672 ;
  assign n674 = n157 | n294 ;
  assign n675 = n441 | n674 ;
  assign n676 = n447 | n675 ;
  assign n677 = n673 | n676 ;
  assign n678 = n670 | n677 ;
  assign n679 = n109 | n229 ;
  assign n680 = n270 | n319 ;
  assign n681 = n205 | n680 ;
  assign n682 = n679 | n681 ;
  assign n683 = n239 | n682 ;
  assign n684 = n121 | n167 ;
  assign n685 = n334 | n684 ;
  assign n686 = n683 | n685 ;
  assign n687 = n473 | n686 ;
  assign n688 = n678 | n687 ;
  assign n689 = n653 | n688 ;
  assign n690 = n513 | n689 ;
  assign n691 = n633 & n690 ;
  assign n692 = n526 & ~n691 ;
  assign n693 = pi4 | n39 ;
  assign n694 = pi5 | n693 ;
  assign n695 = n369 | n694 ;
  assign n696 = pi8 | n695 ;
  assign n697 = ~pi22 & n696 ;
  assign n698 = pi9 & ~n697 ;
  assign n699 = ~pi9 & n697 ;
  assign n700 = n698 | n699 ;
  assign n701 = n219 & n700 ;
  assign n702 = ~n692 & n701 ;
  assign n703 = n692 & ~n701 ;
  assign n704 = n702 | n703 ;
  assign n705 = pi9 | n696 ;
  assign n706 = ~pi22 & n705 ;
  assign n707 = ~pi10 & n706 ;
  assign n708 = pi10 & ~n706 ;
  assign n709 = n707 | n708 ;
  assign n710 = n219 & n709 ;
  assign n711 = ~n704 & n710 ;
  assign n712 = n702 | n711 ;
  assign n713 = ~n528 & n549 ;
  assign n714 = ~n224 & n713 ;
  assign n715 = ( n47 & n552 ) | ( n47 & ~n714 ) | ( n552 & ~n714 );
  assign n716 = ( n47 & ~n550 ) | ( n47 & n714 ) | ( ~n550 & n714 );
  assign n717 = n715 & ~n716 ;
  assign n718 = n358 & ~n537 ;
  assign n719 = n375 | n558 ;
  assign n720 = n537 & n563 ;
  assign n721 = ~n361 & n375 ;
  assign n722 = n720 | n721 ;
  assign n723 = n719 & ~n722 ;
  assign n724 = ~n718 & n723 ;
  assign n725 = ~n546 & n549 ;
  assign n726 = ~n224 & n724 ;
  assign n727 = ( n724 & ~n725 ) | ( n724 & n726 ) | ( ~n725 & n726 );
  assign n728 = n717 & n727 ;
  assign n729 = n633 | n690 ;
  assign n730 = ~n526 & n729 ;
  assign n731 = n633 & ~n690 ;
  assign n732 = ~n633 & n690 ;
  assign n733 = n731 | n732 ;
  assign n734 = n730 | n733 ;
  assign n735 = n224 & ~n734 ;
  assign n736 = n692 | n733 ;
  assign n737 = n224 & ~n736 ;
  assign n738 = ( n692 & ~n735 ) | ( n692 & n737 ) | ( ~n735 & n737 );
  assign n739 = ~n701 & n738 ;
  assign n740 = n47 & n725 ;
  assign n741 = ~n47 & n713 ;
  assign n742 = ( n537 & n552 ) | ( n537 & ~n741 ) | ( n552 & ~n741 );
  assign n743 = ( n537 & ~n550 ) | ( n537 & n741 ) | ( ~n550 & n741 );
  assign n744 = n742 & ~n743 ;
  assign n745 = ~n740 & n744 ;
  assign n746 = n701 & ~n738 ;
  assign n747 = n739 | n746 ;
  assign n748 = n745 & ~n747 ;
  assign n749 = n739 | n748 ;
  assign n750 = n224 & ~n724 ;
  assign n751 = n725 & n750 ;
  assign n752 = ( n717 & n724 ) | ( n717 & ~n751 ) | ( n724 & ~n751 );
  assign n753 = ~n728 & n752 ;
  assign n754 = n749 & n753 ;
  assign n755 = n728 | n754 ;
  assign n756 = n712 & n755 ;
  assign n757 = n557 & ~n567 ;
  assign n758 = n568 | n757 ;
  assign n759 = n712 | n755 ;
  assign n760 = ~n756 & n759 ;
  assign n761 = ~n758 & n760 ;
  assign n762 = n756 | n761 ;
  assign n763 = ~n580 & n582 ;
  assign n764 = n583 | n763 ;
  assign n765 = n762 & ~n764 ;
  assign n766 = ~n762 & n764 ;
  assign n767 = n765 | n766 ;
  assign n768 = n758 & ~n760 ;
  assign n769 = n761 | n768 ;
  assign n770 = n375 & n563 ;
  assign n771 = n358 & ~n375 ;
  assign n772 = n558 | n709 ;
  assign n773 = ~n361 & n709 ;
  assign n774 = n772 & ~n773 ;
  assign n775 = ~n771 & n774 ;
  assign n776 = ~n770 & n775 ;
  assign n777 = ~pi22 & n694 ;
  assign n778 = pi6 & ~pi22 ;
  assign n779 = n777 | n778 ;
  assign n780 = ~pi7 & n779 ;
  assign n781 = pi7 & ~n779 ;
  assign n782 = n780 | n781 ;
  assign n783 = n219 & n782 ;
  assign n784 = n128 | n140 ;
  assign n785 = n263 | n483 ;
  assign n786 = n119 | n145 ;
  assign n787 = n336 | n786 ;
  assign n788 = n268 | n296 ;
  assign n789 = n234 | n293 ;
  assign n790 = n788 | n789 ;
  assign n791 = n787 | n790 ;
  assign n792 = n785 | n791 ;
  assign n793 = n201 | n208 ;
  assign n794 = n435 | n793 ;
  assign n795 = n515 | n794 ;
  assign n796 = n792 | n795 ;
  assign n797 = n312 | n796 ;
  assign n798 = n784 | n797 ;
  assign n799 = n499 | n622 ;
  assign n800 = n192 | n654 ;
  assign n801 = n195 | n238 ;
  assign n802 = n170 | n801 ;
  assign n803 = n800 | n802 ;
  assign n804 = n319 | n342 ;
  assign n805 = n106 | n405 ;
  assign n806 = n200 | n805 ;
  assign n807 = n184 | n806 ;
  assign n808 = n284 | n807 ;
  assign n809 = n206 | n808 ;
  assign n810 = n804 | n809 ;
  assign n811 = n377 | n503 ;
  assign n812 = n274 | n305 ;
  assign n813 = n163 | n285 ;
  assign n814 = n812 | n813 ;
  assign n815 = n233 | n814 ;
  assign n816 = n269 | n334 ;
  assign n817 = n815 | n816 ;
  assign n818 = n811 | n817 ;
  assign n819 = n810 | n818 ;
  assign n820 = n803 | n819 ;
  assign n821 = n403 | n820 ;
  assign n822 = n151 | n433 ;
  assign n823 = n335 | n822 ;
  assign n824 = n821 | n823 ;
  assign n825 = n148 | n824 ;
  assign n826 = n317 | n825 ;
  assign n827 = n136 | n228 ;
  assign n828 = ~n164 & n827 ;
  assign n829 = n271 | n399 ;
  assign n830 = n240 | n829 ;
  assign n831 = n322 | n491 ;
  assign n832 = n176 | n400 ;
  assign n833 = n121 | n832 ;
  assign n834 = n831 | n833 ;
  assign n835 = n830 | n834 ;
  assign n836 = n828 & ~n835 ;
  assign n837 = ~n290 & n836 ;
  assign n838 = n167 | n256 ;
  assign n839 = n157 | n838 ;
  assign n840 = n180 | n191 ;
  assign n841 = n588 | n840 ;
  assign n842 = n839 | n841 ;
  assign n843 = n251 | n842 ;
  assign n844 = n837 & ~n843 ;
  assign n845 = ~n826 & n844 ;
  assign n846 = ~n799 & n845 ;
  assign n847 = ~n798 & n846 ;
  assign n848 = ~n135 & n847 ;
  assign n849 = n297 | n341 ;
  assign n850 = n270 | n849 ;
  assign n851 = n314 | n330 ;
  assign n852 = n157 | n176 ;
  assign n853 = n192 | n313 ;
  assign n854 = n852 | n853 ;
  assign n855 = n851 | n854 ;
  assign n856 = n850 | n855 ;
  assign n857 = n343 | n410 ;
  assign n858 = n271 | n334 ;
  assign n859 = n195 | n858 ;
  assign n860 = n229 | n859 ;
  assign n861 = n247 | n860 ;
  assign n862 = n129 | n170 ;
  assign n863 = n399 | n862 ;
  assign n864 = n158 | n194 ;
  assign n865 = n863 | n864 ;
  assign n866 = n246 | n865 ;
  assign n867 = n861 | n866 ;
  assign n868 = n106 | n433 ;
  assign n869 = n181 | n276 ;
  assign n870 = n868 | n869 ;
  assign n871 = n196 | n870 ;
  assign n872 = n186 | n377 ;
  assign n873 = n871 | n872 ;
  assign n874 = n867 | n873 ;
  assign n875 = n185 | n448 ;
  assign n876 = n210 | n875 ;
  assign n877 = n400 | n444 ;
  assign n878 = n124 | n168 ;
  assign n879 = n227 | n274 ;
  assign n880 = n878 | n879 ;
  assign n881 = n790 | n880 ;
  assign n882 = n877 | n881 ;
  assign n883 = n876 | n882 ;
  assign n884 = n874 | n883 ;
  assign n885 = n230 | n239 ;
  assign n886 = n115 | n180 ;
  assign n887 = n232 | n886 ;
  assign n888 = n305 | n887 ;
  assign n889 = n163 | n201 ;
  assign n890 = n888 | n889 ;
  assign n891 = n885 | n890 ;
  assign n892 = n319 | n891 ;
  assign n893 = n884 | n892 ;
  assign n894 = n857 | n893 ;
  assign n895 = n128 | n263 ;
  assign n896 = n894 | n895 ;
  assign n897 = n856 | n896 ;
  assign n898 = ~n848 & n897 ;
  assign n899 = n690 & ~n898 ;
  assign n900 = n783 & ~n899 ;
  assign n901 = ~n783 & n899 ;
  assign n902 = n900 | n901 ;
  assign n903 = ~pi22 & n695 ;
  assign n904 = ~pi8 & n903 ;
  assign n905 = pi8 & ~n903 ;
  assign n906 = n904 | n905 ;
  assign n907 = n219 & n906 ;
  assign n908 = ~n902 & n907 ;
  assign n909 = n900 | n908 ;
  assign n910 = n776 & n909 ;
  assign n911 = ~n730 & n733 ;
  assign n912 = n224 & n911 ;
  assign n913 = ~n692 & n733 ;
  assign n914 = ~n224 & n913 ;
  assign n915 = n47 | n736 ;
  assign n916 = n47 & ~n734 ;
  assign n917 = n915 & ~n916 ;
  assign n918 = ~n914 & n917 ;
  assign n919 = ~n912 & n918 ;
  assign n920 = n537 & n725 ;
  assign n921 = ~n537 & n713 ;
  assign n922 = ( n375 & n552 ) | ( n375 & ~n921 ) | ( n552 & ~n921 );
  assign n923 = ( n375 & ~n550 ) | ( n375 & n921 ) | ( ~n550 & n921 );
  assign n924 = n922 & ~n923 ;
  assign n925 = ~n920 & n924 ;
  assign n926 = n919 & n925 ;
  assign n927 = n563 & n709 ;
  assign n928 = n358 & ~n709 ;
  assign n929 = n558 | n700 ;
  assign n930 = ~n361 & n700 ;
  assign n931 = n929 & ~n930 ;
  assign n932 = ~n928 & n931 ;
  assign n933 = ~n927 & n932 ;
  assign n934 = n919 & ~n925 ;
  assign n935 = ~n919 & n925 ;
  assign n936 = n934 | n935 ;
  assign n937 = n933 & n936 ;
  assign n938 = n926 | n937 ;
  assign n939 = n776 | n909 ;
  assign n940 = ~n910 & n939 ;
  assign n941 = n938 & n940 ;
  assign n942 = n910 | n941 ;
  assign n943 = n704 & ~n710 ;
  assign n944 = n711 | n943 ;
  assign n945 = n942 & ~n944 ;
  assign n946 = n749 | n753 ;
  assign n947 = ~n754 & n946 ;
  assign n948 = ~n942 & n944 ;
  assign n949 = n945 | n948 ;
  assign n950 = ~n945 & n949 ;
  assign n951 = ( n945 & n947 ) | ( n945 & ~n950 ) | ( n947 & ~n950 );
  assign n952 = ~n769 & n951 ;
  assign n953 = n769 & ~n951 ;
  assign n954 = n952 | n953 ;
  assign n955 = n563 & n700 ;
  assign n956 = n358 & ~n700 ;
  assign n957 = n558 | n906 ;
  assign n958 = ~n361 & n906 ;
  assign n959 = n957 & ~n958 ;
  assign n960 = ~n956 & n959 ;
  assign n961 = ~n955 & n960 ;
  assign n962 = n375 & n725 ;
  assign n963 = ~n375 & n713 ;
  assign n964 = ( n552 & n709 ) | ( n552 & ~n963 ) | ( n709 & ~n963 );
  assign n965 = ( ~n550 & n709 ) | ( ~n550 & n963 ) | ( n709 & n963 );
  assign n966 = n964 & ~n965 ;
  assign n967 = ~n962 & n966 ;
  assign n968 = n961 & n967 ;
  assign n969 = n186 | n499 ;
  assign n970 = n305 | n969 ;
  assign n971 = n294 | n317 ;
  assign n972 = n321 | n971 ;
  assign n973 = n185 | n286 ;
  assign n974 = n264 | n973 ;
  assign n975 = n343 | n974 ;
  assign n976 = n972 | n975 ;
  assign n977 = n970 | n976 ;
  assign n978 = n865 | n977 ;
  assign n979 = n466 | n978 ;
  assign n980 = n433 | n979 ;
  assign n981 = n284 | n980 ;
  assign n982 = n201 | n981 ;
  assign n983 = n230 | n982 ;
  assign n984 = n275 | n328 ;
  assign n985 = n380 | n621 ;
  assign n986 = n816 | n985 ;
  assign n987 = n128 | n247 ;
  assign n988 = n109 | n987 ;
  assign n989 = n986 | n988 ;
  assign n990 = n984 | n989 ;
  assign n991 = n233 | n990 ;
  assign n992 = n157 | n168 ;
  assign n993 = n991 | n992 ;
  assign n994 = n240 | n271 ;
  assign n995 = n296 | n994 ;
  assign n996 = n281 | n335 ;
  assign n997 = n192 | n270 ;
  assign n998 = n996 | n997 ;
  assign n999 = n995 | n998 ;
  assign n1000 = n191 | n320 ;
  assign n1001 = n318 | n389 ;
  assign n1002 = n1000 | n1001 ;
  assign n1003 = n207 | n263 ;
  assign n1004 = n204 | n503 ;
  assign n1005 = n1003 | n1004 ;
  assign n1006 = n1002 | n1005 ;
  assign n1007 = n999 | n1006 ;
  assign n1008 = n993 | n1007 ;
  assign n1009 = n227 | n383 ;
  assign n1010 = n117 | n209 ;
  assign n1011 = n1009 | n1010 ;
  assign n1012 = n406 | n1011 ;
  assign n1013 = n828 & ~n1012 ;
  assign n1014 = n167 | n297 ;
  assign n1015 = n654 | n1014 ;
  assign n1016 = n268 | n1015 ;
  assign n1017 = n1013 & ~n1016 ;
  assign n1018 = ~n1008 & n1017 ;
  assign n1019 = ~n152 & n1018 ;
  assign n1020 = ~n983 & n1019 ;
  assign n1021 = ~n180 & n1020 ;
  assign n1022 = ~n274 & n1021 ;
  assign n1023 = ~n316 & n1022 ;
  assign n1024 = ~n377 & n1023 ;
  assign n1025 = n378 | n851 ;
  assign n1026 = n243 | n318 ;
  assign n1027 = n1025 | n1026 ;
  assign n1028 = n304 | n341 ;
  assign n1029 = n146 | n399 ;
  assign n1030 = n124 | n1009 ;
  assign n1031 = n608 | n1030 ;
  assign n1032 = n292 | n1031 ;
  assign n1033 = n1029 | n1032 ;
  assign n1034 = n240 | n320 ;
  assign n1035 = n193 | n1034 ;
  assign n1036 = n272 | n281 ;
  assign n1037 = n1035 | n1036 ;
  assign n1038 = n442 | n833 ;
  assign n1039 = n1037 | n1038 ;
  assign n1040 = n206 | n1039 ;
  assign n1041 = n1033 | n1040 ;
  assign n1042 = n868 | n1041 ;
  assign n1043 = n1028 | n1042 ;
  assign n1044 = n140 | n321 ;
  assign n1045 = n319 | n401 ;
  assign n1046 = n129 | n285 ;
  assign n1047 = n207 | n1046 ;
  assign n1048 = n269 | n1047 ;
  assign n1049 = n337 | n1048 ;
  assign n1050 = n278 | n1049 ;
  assign n1051 = n663 | n1050 ;
  assign n1052 = n1045 | n1051 ;
  assign n1053 = n294 | n434 ;
  assign n1054 = n167 | n1053 ;
  assign n1055 = n801 | n1054 ;
  assign n1056 = n128 | n377 ;
  assign n1057 = n177 | n1056 ;
  assign n1058 = n588 | n1057 ;
  assign n1059 = n1055 | n1058 ;
  assign n1060 = ~n501 & n827 ;
  assign n1061 = ~n887 & n1060 ;
  assign n1062 = ~n249 & n1061 ;
  assign n1063 = ~n1059 & n1062 ;
  assign n1064 = ~n190 & n1063 ;
  assign n1065 = ~n117 & n1064 ;
  assign n1066 = n403 | n622 ;
  assign n1067 = n654 | n1066 ;
  assign n1068 = n392 | n1067 ;
  assign n1069 = n1065 & ~n1068 ;
  assign n1070 = ~n148 & n1069 ;
  assign n1071 = ~n210 & n1070 ;
  assign n1072 = ~n1052 & n1071 ;
  assign n1073 = ~n1044 & n1072 ;
  assign n1074 = ~n1043 & n1073 ;
  assign n1075 = ~n1027 & n1074 ;
  assign n1076 = n1024 | n1075 ;
  assign n1077 = ~n848 & n1076 ;
  assign n1078 = n1024 & ~n1077 ;
  assign n1079 = ~pi6 & n777 ;
  assign n1080 = pi6 & ~n777 ;
  assign n1081 = n1079 | n1080 ;
  assign n1082 = n219 & n1081 ;
  assign n1083 = ~n1024 & n1077 ;
  assign n1084 = n1078 | n1083 ;
  assign n1085 = n1082 & ~n1084 ;
  assign n1086 = n1078 | n1085 ;
  assign n1087 = n961 | n967 ;
  assign n1088 = ~n968 & n1087 ;
  assign n1089 = n1086 & n1088 ;
  assign n1090 = n968 | n1089 ;
  assign n1091 = n224 | n899 ;
  assign n1092 = n848 & ~n897 ;
  assign n1093 = n690 | n1092 ;
  assign n1094 = n848 & n897 ;
  assign n1095 = n848 | n897 ;
  assign n1096 = ~n1094 & n1095 ;
  assign n1097 = n1093 & n1096 ;
  assign n1098 = n224 & n1097 ;
  assign n1099 = n899 | n1096 ;
  assign n1100 = ~n1098 & n1099 ;
  assign n1101 = n1091 & n1100 ;
  assign n1102 = ~n783 & n1101 ;
  assign n1103 = n783 & ~n1101 ;
  assign n1104 = n1102 | n1103 ;
  assign n1105 = n47 & n911 ;
  assign n1106 = ~n47 & n913 ;
  assign n1107 = ( n537 & n736 ) | ( n537 & ~n1106 ) | ( n736 & ~n1106 );
  assign n1108 = ( n537 & ~n734 ) | ( n537 & n1106 ) | ( ~n734 & n1106 );
  assign n1109 = n1107 & ~n1108 ;
  assign n1110 = ~n1105 & n1109 ;
  assign n1111 = ~n1104 & n1110 ;
  assign n1112 = n1102 | n1111 ;
  assign n1113 = n1090 & n1112 ;
  assign n1114 = n1090 | n1112 ;
  assign n1115 = ~n1113 & n1114 ;
  assign n1116 = n902 & ~n907 ;
  assign n1117 = n908 | n1116 ;
  assign n1118 = n1115 & ~n1117 ;
  assign n1119 = n1113 | n1118 ;
  assign n1120 = ~n745 & n747 ;
  assign n1121 = n748 | n1120 ;
  assign n1122 = n1119 & ~n1121 ;
  assign n1123 = ~n1119 & n1121 ;
  assign n1124 = n1122 | n1123 ;
  assign n1125 = n938 | n940 ;
  assign n1126 = ~n941 & n1125 ;
  assign n1127 = ~n1124 & n1126 ;
  assign n1128 = n1122 | n1127 ;
  assign n1129 = n947 & ~n949 ;
  assign n1130 = ~n947 & n949 ;
  assign n1131 = n1129 | n1130 ;
  assign n1132 = n1128 & ~n1131 ;
  assign n1133 = n933 | n936 ;
  assign n1134 = ~n937 & n1133 ;
  assign n1135 = n1104 & ~n1110 ;
  assign n1136 = n1111 | n1135 ;
  assign n1137 = n563 & n906 ;
  assign n1138 = n358 & ~n906 ;
  assign n1139 = n558 | n782 ;
  assign n1140 = ~n361 & n782 ;
  assign n1141 = n1139 & ~n1140 ;
  assign n1142 = ~n1138 & n1141 ;
  assign n1143 = ~n1137 & n1142 ;
  assign n1144 = n552 | n700 ;
  assign n1145 = ~n550 & n700 ;
  assign n1146 = n1144 & ~n1145 ;
  assign n1147 = ( n709 & n725 ) | ( n709 & ~n1146 ) | ( n725 & ~n1146 );
  assign n1148 = ( n709 & ~n713 ) | ( n709 & n1146 ) | ( ~n713 & n1146 );
  assign n1149 = ~n1147 & n1148 ;
  assign n1150 = n1093 & ~n1096 ;
  assign n1151 = ~n899 & n1096 ;
  assign n1152 = ~n47 & n1151 ;
  assign n1153 = n47 & n1097 ;
  assign n1154 = n1152 | n1153 ;
  assign n1155 = ( n224 & n1150 ) | ( n224 & n1154 ) | ( n1150 & n1154 );
  assign n1156 = ( n224 & n1099 ) | ( n224 & ~n1154 ) | ( n1099 & ~n1154 );
  assign n1157 = ~n1155 & n1156 ;
  assign n1158 = ( n1143 & n1149 ) | ( n1143 & n1157 ) | ( n1149 & n1157 );
  assign n1159 = ~n1136 & n1158 ;
  assign n1160 = n1086 | n1088 ;
  assign n1161 = ~n1089 & n1160 ;
  assign n1162 = n1136 | n1158 ;
  assign n1163 = ( ~n1158 & n1159 ) | ( ~n1158 & n1162 ) | ( n1159 & n1162 );
  assign n1164 = n1161 & ~n1163 ;
  assign n1165 = n1159 | n1164 ;
  assign n1166 = n1134 & n1165 ;
  assign n1167 = n1134 | n1165 ;
  assign n1168 = ~n1166 & n1167 ;
  assign n1169 = ~n1115 & n1117 ;
  assign n1170 = n1118 | n1169 ;
  assign n1171 = n1168 & ~n1170 ;
  assign n1172 = n1166 | n1171 ;
  assign n1173 = n1124 & ~n1126 ;
  assign n1174 = n1127 | n1173 ;
  assign n1175 = n1172 & ~n1174 ;
  assign n1176 = ~n1082 & n1084 ;
  assign n1177 = n1085 | n1176 ;
  assign n1178 = n537 & n911 ;
  assign n1179 = ~n537 & n913 ;
  assign n1180 = ( n375 & n736 ) | ( n375 & ~n1179 ) | ( n736 & ~n1179 );
  assign n1181 = ( n375 & ~n734 ) | ( n375 & n1179 ) | ( ~n734 & n1179 );
  assign n1182 = n1180 & ~n1181 ;
  assign n1183 = ~n1178 & n1182 ;
  assign n1184 = ~n1177 & n1183 ;
  assign n1185 = n1177 & ~n1183 ;
  assign n1186 = n1184 | n1185 ;
  assign n1187 = ~pi22 & n693 ;
  assign n1188 = pi5 & ~n1187 ;
  assign n1189 = ~pi5 & n1187 ;
  assign n1190 = n1188 | n1189 ;
  assign n1191 = n219 & n1190 ;
  assign n1192 = n1024 & ~n1191 ;
  assign n1193 = n1024 & ~n1075 ;
  assign n1194 = ~n1024 & n1075 ;
  assign n1195 = n1193 | n1194 ;
  assign n1196 = n224 & ~n1195 ;
  assign n1197 = n1077 | n1196 ;
  assign n1198 = n1024 & n1075 ;
  assign n1199 = n848 & ~n1198 ;
  assign n1200 = n1196 & ~n1199 ;
  assign n1201 = n1197 & ~n1200 ;
  assign n1202 = ~n1192 & n1201 ;
  assign n1203 = ~n1024 & n1191 ;
  assign n1204 = n1202 | n1203 ;
  assign n1205 = ~n1186 & n1204 ;
  assign n1206 = n1184 | n1205 ;
  assign n1207 = n47 & n1150 ;
  assign n1208 = n47 | n1099 ;
  assign n1209 = ( n537 & ~n1151 ) | ( n537 & n1208 ) | ( ~n1151 & n1208 );
  assign n1210 = ( n537 & n1097 ) | ( n537 & ~n1208 ) | ( n1097 & ~n1208 );
  assign n1211 = n1209 & ~n1210 ;
  assign n1212 = ~n1207 & n1211 ;
  assign n1213 = n375 & n911 ;
  assign n1214 = ~n375 & n913 ;
  assign n1215 = ( n709 & n736 ) | ( n709 & ~n1214 ) | ( n736 & ~n1214 );
  assign n1216 = ( n709 & ~n734 ) | ( n709 & n1214 ) | ( ~n734 & n1214 );
  assign n1217 = n1215 & ~n1216 ;
  assign n1218 = ~n1213 & n1217 ;
  assign n1219 = n700 & n725 ;
  assign n1220 = ~n700 & n713 ;
  assign n1221 = ( n552 & n906 ) | ( n552 & ~n1220 ) | ( n906 & ~n1220 );
  assign n1222 = ( ~n550 & n906 ) | ( ~n550 & n1220 ) | ( n906 & n1220 );
  assign n1223 = n1221 & ~n1222 ;
  assign n1224 = ~n1219 & n1223 ;
  assign n1225 = ( n1212 & n1218 ) | ( n1212 & n1224 ) | ( n1218 & n1224 );
  assign n1226 = ( n1143 & ~n1149 ) | ( n1143 & n1157 ) | ( ~n1149 & n1157 );
  assign n1227 = ( ~n1143 & n1149 ) | ( ~n1143 & n1226 ) | ( n1149 & n1226 );
  assign n1228 = ( ~n1157 & n1226 ) | ( ~n1157 & n1227 ) | ( n1226 & n1227 );
  assign n1229 = n1225 & n1228 ;
  assign n1230 = ~pi22 & n39 ;
  assign n1231 = ~pi4 & n1230 ;
  assign n1232 = pi4 & ~n1230 ;
  assign n1233 = n1231 | n1232 ;
  assign n1234 = n219 & n1233 ;
  assign n1235 = ~n1024 & n1234 ;
  assign n1236 = n1024 & ~n1234 ;
  assign n1237 = n1195 & ~n1199 ;
  assign n1238 = n224 & n1237 ;
  assign n1239 = n1195 | n1199 ;
  assign n1240 = n47 & ~n1239 ;
  assign n1241 = n1077 | n1195 ;
  assign n1242 = n47 | n1241 ;
  assign n1243 = ~n1077 & n1195 ;
  assign n1244 = ~n224 & n1243 ;
  assign n1245 = n1242 & ~n1244 ;
  assign n1246 = ~n1240 & n1245 ;
  assign n1247 = ~n1238 & n1246 ;
  assign n1248 = ~n1236 & n1247 ;
  assign n1249 = ~n1235 & n1248 ;
  assign n1250 = n1235 | n1249 ;
  assign n1251 = n563 & n782 ;
  assign n1252 = n358 & ~n782 ;
  assign n1253 = n558 | n1081 ;
  assign n1254 = ~n361 & n1081 ;
  assign n1255 = n1253 & ~n1254 ;
  assign n1256 = ~n1252 & n1255 ;
  assign n1257 = ~n1251 & n1256 ;
  assign n1258 = n1250 & n1257 ;
  assign n1259 = n1250 | n1257 ;
  assign n1260 = ~n1258 & n1259 ;
  assign n1261 = n709 & n911 ;
  assign n1262 = ~n709 & n913 ;
  assign n1263 = ( n700 & n736 ) | ( n700 & ~n1262 ) | ( n736 & ~n1262 );
  assign n1264 = ( n700 & ~n734 ) | ( n700 & n1262 ) | ( ~n734 & n1262 );
  assign n1265 = n1263 & ~n1264 ;
  assign n1266 = ~n1261 & n1265 ;
  assign n1267 = n537 & n1150 ;
  assign n1268 = n537 | n1099 ;
  assign n1269 = ( n375 & ~n1151 ) | ( n375 & n1268 ) | ( ~n1151 & n1268 );
  assign n1270 = ( n375 & n1097 ) | ( n375 & ~n1268 ) | ( n1097 & ~n1268 );
  assign n1271 = n1269 & ~n1270 ;
  assign n1272 = ~n1267 & n1271 ;
  assign n1273 = n725 & n906 ;
  assign n1274 = n713 & ~n906 ;
  assign n1275 = ( n552 & n782 ) | ( n552 & ~n1274 ) | ( n782 & ~n1274 );
  assign n1276 = ( ~n550 & n782 ) | ( ~n550 & n1274 ) | ( n782 & n1274 );
  assign n1277 = n1275 & ~n1276 ;
  assign n1278 = ~n1273 & n1277 ;
  assign n1279 = ( n1266 & n1272 ) | ( n1266 & n1278 ) | ( n1272 & n1278 );
  assign n1280 = n1260 & n1279 ;
  assign n1281 = n1258 | n1280 ;
  assign n1282 = n1225 | n1228 ;
  assign n1283 = ~n1229 & n1282 ;
  assign n1284 = n1281 & n1283 ;
  assign n1285 = n1229 | n1284 ;
  assign n1286 = n1206 & n1285 ;
  assign n1287 = n1206 | n1285 ;
  assign n1288 = ~n1286 & n1287 ;
  assign n1289 = ~n1161 & n1163 ;
  assign n1290 = n1164 | n1289 ;
  assign n1291 = n1288 & ~n1290 ;
  assign n1292 = n1286 | n1291 ;
  assign n1293 = ~n1168 & n1170 ;
  assign n1294 = n1171 | n1293 ;
  assign n1295 = n1292 & ~n1294 ;
  assign n1296 = n1192 | n1203 ;
  assign n1297 = n1201 | n1296 ;
  assign n1298 = n1201 & n1296 ;
  assign n1299 = n1297 & ~n1298 ;
  assign n1300 = ( n1212 & n1224 ) | ( n1212 & ~n1225 ) | ( n1224 & ~n1225 );
  assign n1301 = ( n1218 & ~n1225 ) | ( n1218 & n1300 ) | ( ~n1225 & n1300 );
  assign n1302 = ~n1299 & n1301 ;
  assign n1303 = n1299 & ~n1301 ;
  assign n1304 = n1302 | n1303 ;
  assign n1305 = n563 & n1081 ;
  assign n1306 = n358 & ~n1081 ;
  assign n1307 = n558 | n1190 ;
  assign n1308 = ~n361 & n1190 ;
  assign n1309 = n1307 & ~n1308 ;
  assign n1310 = ~n1306 & n1309 ;
  assign n1311 = ~n1305 & n1310 ;
  assign n1312 = pi3 & ~n28 ;
  assign n1313 = ~pi3 & n28 ;
  assign n1314 = n1312 | n1313 ;
  assign n1315 = n219 & n1314 ;
  assign n1316 = n181 | n320 ;
  assign n1317 = n207 | n377 ;
  assign n1318 = n1316 | n1317 ;
  assign n1319 = n383 | n499 ;
  assign n1320 = n329 | n622 ;
  assign n1321 = n124 | n319 ;
  assign n1322 = n192 | n1321 ;
  assign n1323 = n178 | n1322 ;
  assign n1324 = n465 | n1323 ;
  assign n1325 = n381 | n886 ;
  assign n1326 = n1324 | n1325 ;
  assign n1327 = n196 | n1326 ;
  assign n1328 = n167 | n1327 ;
  assign n1329 = n263 | n313 ;
  assign n1330 = n1328 | n1329 ;
  assign n1331 = n158 | n1330 ;
  assign n1332 = n297 | n343 ;
  assign n1333 = ~n305 & n827 ;
  assign n1334 = n243 | n336 ;
  assign n1335 = n246 | n1334 ;
  assign n1336 = n1333 & ~n1335 ;
  assign n1337 = ~n1332 & n1336 ;
  assign n1338 = ~n251 & n1337 ;
  assign n1339 = ~n403 & n1338 ;
  assign n1340 = ~n393 & n1339 ;
  assign n1341 = ~n1331 & n1340 ;
  assign n1342 = ~n156 & n1341 ;
  assign n1343 = n204 | n623 ;
  assign n1344 = n195 | n1343 ;
  assign n1345 = n601 | n1344 ;
  assign n1346 = n290 | n1345 ;
  assign n1347 = n164 | n1346 ;
  assign n1348 = n1342 & ~n1347 ;
  assign n1349 = ~n1320 & n1348 ;
  assign n1350 = ~n1319 & n1349 ;
  assign n1351 = ~n1318 & n1350 ;
  assign n1352 = ~n382 & n1351 ;
  assign n1353 = n224 & n1352 ;
  assign n1354 = n1024 | n1353 ;
  assign n1355 = n1315 & ~n1354 ;
  assign n1356 = ~n1315 & n1354 ;
  assign n1357 = n1355 | n1356 ;
  assign n1358 = n47 & n1237 ;
  assign n1359 = n537 & ~n1239 ;
  assign n1360 = n537 | n1241 ;
  assign n1361 = ~n47 & n1243 ;
  assign n1362 = n1360 & ~n1361 ;
  assign n1363 = ~n1359 & n1362 ;
  assign n1364 = ~n1358 & n1363 ;
  assign n1365 = ~n1357 & n1364 ;
  assign n1366 = n1355 | n1365 ;
  assign n1367 = n1311 & n1366 ;
  assign n1368 = n1311 | n1366 ;
  assign n1369 = ~n1367 & n1368 ;
  assign n1370 = n700 & n911 ;
  assign n1371 = ~n700 & n913 ;
  assign n1372 = ( n736 & n906 ) | ( n736 & ~n1371 ) | ( n906 & ~n1371 );
  assign n1373 = ( ~n734 & n906 ) | ( ~n734 & n1371 ) | ( n906 & n1371 );
  assign n1374 = n1372 & ~n1373 ;
  assign n1375 = ~n1370 & n1374 ;
  assign n1376 = n375 & n1150 ;
  assign n1377 = n375 | n1099 ;
  assign n1378 = ( n709 & ~n1151 ) | ( n709 & n1377 ) | ( ~n1151 & n1377 );
  assign n1379 = ( n709 & n1097 ) | ( n709 & ~n1377 ) | ( n1097 & ~n1377 );
  assign n1380 = n1378 & ~n1379 ;
  assign n1381 = ~n1376 & n1380 ;
  assign n1382 = n725 & n782 ;
  assign n1383 = n713 & ~n782 ;
  assign n1384 = ( n552 & n1081 ) | ( n552 & ~n1383 ) | ( n1081 & ~n1383 );
  assign n1385 = ( ~n550 & n1081 ) | ( ~n550 & n1383 ) | ( n1081 & n1383 );
  assign n1386 = n1384 & ~n1385 ;
  assign n1387 = ~n1382 & n1386 ;
  assign n1388 = ( n1375 & n1381 ) | ( n1375 & n1387 ) | ( n1381 & n1387 );
  assign n1389 = n1369 & n1388 ;
  assign n1390 = n1367 | n1389 ;
  assign n1391 = ~n1304 & n1390 ;
  assign n1392 = n1302 | n1391 ;
  assign n1393 = n1186 & ~n1204 ;
  assign n1394 = n1205 | n1393 ;
  assign n1395 = n1392 & ~n1394 ;
  assign n1396 = n1281 | n1283 ;
  assign n1397 = ~n1284 & n1396 ;
  assign n1398 = ~n1302 & n1394 ;
  assign n1399 = ~n1391 & n1398 ;
  assign n1400 = n1397 & ~n1399 ;
  assign n1401 = ~n1395 & n1400 ;
  assign n1402 = n1395 | n1401 ;
  assign n1403 = ~n1288 & n1290 ;
  assign n1404 = n1291 | n1403 ;
  assign n1405 = n1402 & ~n1404 ;
  assign n1406 = n1395 | n1399 ;
  assign n1407 = ~n1397 & n1406 ;
  assign n1408 = n1260 | n1279 ;
  assign n1409 = ~n1280 & n1408 ;
  assign n1410 = n563 & n1314 ;
  assign n1411 = n353 & n558 ;
  assign n1412 = ~n1410 & n1411 ;
  assign n1413 = n224 & ~n1352 ;
  assign n1414 = n1024 & ~n1413 ;
  assign n1415 = ~n1024 & n1413 ;
  assign n1416 = n47 & n1352 ;
  assign n1417 = n1415 | n1416 ;
  assign n1418 = n1414 | n1417 ;
  assign n1419 = n1412 & ~n1418 ;
  assign n1420 = n563 & n1190 ;
  assign n1421 = n358 & ~n1190 ;
  assign n1422 = n558 | n1233 ;
  assign n1423 = ~n361 & n1233 ;
  assign n1424 = n1422 & ~n1423 ;
  assign n1425 = ~n1421 & n1424 ;
  assign n1426 = ~n1420 & n1425 ;
  assign n1427 = n1419 & n1426 ;
  assign n1428 = n1419 | n1426 ;
  assign n1429 = ~n1427 & n1428 ;
  assign n1430 = n709 & n1150 ;
  assign n1431 = n709 | n1099 ;
  assign n1432 = ( n700 & ~n1151 ) | ( n700 & n1431 ) | ( ~n1151 & n1431 );
  assign n1433 = ( n700 & n1097 ) | ( n700 & ~n1431 ) | ( n1097 & ~n1431 );
  assign n1434 = n1432 & ~n1433 ;
  assign n1435 = ~n1430 & n1434 ;
  assign n1436 = n906 & n911 ;
  assign n1437 = ~n906 & n913 ;
  assign n1438 = ( n736 & n782 ) | ( n736 & ~n1437 ) | ( n782 & ~n1437 );
  assign n1439 = ( ~n734 & n782 ) | ( ~n734 & n1437 ) | ( n782 & n1437 );
  assign n1440 = n1438 & ~n1439 ;
  assign n1441 = ~n1436 & n1440 ;
  assign n1442 = n725 & n1081 ;
  assign n1443 = n713 & ~n1081 ;
  assign n1444 = ( n552 & n1190 ) | ( n552 & ~n1443 ) | ( n1190 & ~n1443 );
  assign n1445 = ( ~n550 & n1190 ) | ( ~n550 & n1443 ) | ( n1190 & n1443 );
  assign n1446 = n1444 & ~n1445 ;
  assign n1447 = ~n1442 & n1446 ;
  assign n1448 = ( n1435 & n1441 ) | ( n1435 & n1447 ) | ( n1441 & n1447 );
  assign n1449 = n1429 & n1448 ;
  assign n1450 = n1427 | n1449 ;
  assign n1451 = n1236 | n1250 ;
  assign n1452 = n1247 & ~n1249 ;
  assign n1453 = n1451 & ~n1452 ;
  assign n1454 = n1450 | n1453 ;
  assign n1455 = n1450 & n1453 ;
  assign n1456 = n1454 & ~n1455 ;
  assign n1457 = ( n1266 & n1278 ) | ( n1266 & ~n1279 ) | ( n1278 & ~n1279 );
  assign n1458 = ( n1272 & ~n1279 ) | ( n1272 & n1457 ) | ( ~n1279 & n1457 );
  assign n1459 = ~n1456 & n1458 ;
  assign n1460 = n1450 & ~n1453 ;
  assign n1461 = n1459 | n1460 ;
  assign n1462 = n1409 & n1461 ;
  assign n1463 = n1409 | n1461 ;
  assign n1464 = ~n1462 & n1463 ;
  assign n1465 = n1304 & ~n1390 ;
  assign n1466 = n1391 | n1465 ;
  assign n1467 = n1464 & ~n1466 ;
  assign n1468 = n1462 | n1467 ;
  assign n1469 = ~n1401 & n1468 ;
  assign n1470 = ~n1407 & n1469 ;
  assign n1471 = ~n1464 & n1466 ;
  assign n1472 = n1467 | n1471 ;
  assign n1473 = n563 & n1233 ;
  assign n1474 = n358 & ~n1233 ;
  assign n1475 = n1473 | n1474 ;
  assign n1476 = n558 | n1314 ;
  assign n1477 = ~n361 & n1314 ;
  assign n1478 = n1476 & ~n1477 ;
  assign n1479 = ~n1475 & n1478 ;
  assign n1480 = n537 & n1237 ;
  assign n1481 = n375 & ~n1239 ;
  assign n1482 = n375 | n1241 ;
  assign n1483 = ~n537 & n1243 ;
  assign n1484 = n1482 & ~n1483 ;
  assign n1485 = ~n1481 & n1484 ;
  assign n1486 = ~n1480 & n1485 ;
  assign n1487 = n1479 & n1486 ;
  assign n1488 = n1479 | n1486 ;
  assign n1489 = ~n1412 & n1418 ;
  assign n1490 = n1419 | n1489 ;
  assign n1491 = n1488 & ~n1490 ;
  assign n1492 = n1487 | n1491 ;
  assign n1493 = n1357 & ~n1364 ;
  assign n1494 = n1365 | n1493 ;
  assign n1495 = n1492 & ~n1494 ;
  assign n1496 = ~n1492 & n1494 ;
  assign n1497 = n1495 | n1496 ;
  assign n1498 = ( n1375 & n1387 ) | ( n1375 & ~n1388 ) | ( n1387 & ~n1388 );
  assign n1499 = ( n1381 & ~n1388 ) | ( n1381 & n1498 ) | ( ~n1388 & n1498 );
  assign n1500 = ~n1497 & n1499 ;
  assign n1501 = n1495 | n1500 ;
  assign n1502 = n1369 | n1388 ;
  assign n1503 = ~n1389 & n1502 ;
  assign n1504 = n1501 & n1503 ;
  assign n1505 = n1501 | n1503 ;
  assign n1506 = ~n1504 & n1505 ;
  assign n1507 = n1456 & ~n1458 ;
  assign n1508 = n1459 | n1507 ;
  assign n1509 = n1506 & ~n1508 ;
  assign n1510 = n1504 | n1509 ;
  assign n1511 = ~n1472 & n1510 ;
  assign n1512 = n1472 & ~n1510 ;
  assign n1513 = n1511 | n1512 ;
  assign n1514 = n375 & n1237 ;
  assign n1515 = n709 & ~n1239 ;
  assign n1516 = n709 | n1241 ;
  assign n1517 = ~n375 & n1243 ;
  assign n1518 = n1516 & ~n1517 ;
  assign n1519 = ~n1515 & n1518 ;
  assign n1520 = ~n1514 & n1519 ;
  assign n1521 = n47 & ~n1352 ;
  assign n1522 = n1024 & ~n1521 ;
  assign n1523 = n537 & n1352 ;
  assign n1524 = ~n1024 & n1521 ;
  assign n1525 = n1523 | n1524 ;
  assign n1526 = n1522 | n1525 ;
  assign n1527 = n1520 & ~n1526 ;
  assign n1528 = ~n1520 & n1526 ;
  assign n1529 = n1527 | n1528 ;
  assign n1530 = n725 & n1190 ;
  assign n1531 = n713 & ~n1190 ;
  assign n1532 = ( n552 & n1233 ) | ( n552 & ~n1531 ) | ( n1233 & ~n1531 );
  assign n1533 = ( ~n550 & n1233 ) | ( ~n550 & n1531 ) | ( n1233 & n1531 );
  assign n1534 = n1532 & ~n1533 ;
  assign n1535 = ~n1530 & n1534 ;
  assign n1536 = ~n1529 & n1535 ;
  assign n1537 = n1527 | n1536 ;
  assign n1538 = n700 & n1150 ;
  assign n1539 = n700 | n1099 ;
  assign n1540 = ( n906 & ~n1151 ) | ( n906 & n1539 ) | ( ~n1151 & n1539 );
  assign n1541 = ( n906 & n1097 ) | ( n906 & ~n1539 ) | ( n1097 & ~n1539 );
  assign n1542 = n1540 & ~n1541 ;
  assign n1543 = ~n1538 & n1542 ;
  assign n1544 = n782 & n911 ;
  assign n1545 = ~n782 & n913 ;
  assign n1546 = ( n736 & n1081 ) | ( n736 & ~n1545 ) | ( n1081 & ~n1545 );
  assign n1547 = ( ~n734 & n1081 ) | ( ~n734 & n1545 ) | ( n1081 & n1545 );
  assign n1548 = n1546 & ~n1547 ;
  assign n1549 = ~n1544 & n1548 ;
  assign n1550 = n375 & n1352 ;
  assign n1551 = n537 & ~n1352 ;
  assign n1552 = ~n1024 & n1551 ;
  assign n1553 = n1024 & ~n1551 ;
  assign n1554 = n1552 | n1553 ;
  assign n1555 = n1550 | n1554 ;
  assign n1556 = n725 & n1314 ;
  assign n1557 = n528 & ~n1556 ;
  assign n1558 = ~n1555 & n1557 ;
  assign n1559 = ( n1543 & n1549 ) | ( n1543 & n1558 ) | ( n1549 & n1558 );
  assign n1560 = n1537 & n1559 ;
  assign n1561 = n1537 | n1559 ;
  assign n1562 = ~n1560 & n1561 ;
  assign n1563 = ( n1435 & n1447 ) | ( n1435 & ~n1448 ) | ( n1447 & ~n1448 );
  assign n1564 = ( n1441 & ~n1448 ) | ( n1441 & n1563 ) | ( ~n1448 & n1563 );
  assign n1565 = n1562 & n1564 ;
  assign n1566 = n1560 | n1565 ;
  assign n1567 = n1429 | n1448 ;
  assign n1568 = ~n1449 & n1567 ;
  assign n1569 = n1566 & n1568 ;
  assign n1570 = n1566 | n1568 ;
  assign n1571 = ~n1569 & n1570 ;
  assign n1572 = n1497 & ~n1499 ;
  assign n1573 = n1500 | n1572 ;
  assign n1574 = n1571 & ~n1573 ;
  assign n1575 = n1569 | n1574 ;
  assign n1576 = ~n1506 & n1508 ;
  assign n1577 = n1509 | n1576 ;
  assign n1578 = n1575 & ~n1577 ;
  assign n1579 = ~n1571 & n1573 ;
  assign n1580 = n1574 | n1579 ;
  assign n1581 = n558 & n1314 ;
  assign n1582 = ~n563 & n1581 ;
  assign n1583 = n353 | n1582 ;
  assign n1584 = ~n709 & n1243 ;
  assign n1585 = n700 | n1241 ;
  assign n1586 = n709 & n1237 ;
  assign n1587 = n700 & ~n1239 ;
  assign n1588 = n1586 | n1587 ;
  assign n1589 = n1585 & ~n1588 ;
  assign n1590 = ~n1584 & n1589 ;
  assign n1591 = n911 & n1081 ;
  assign n1592 = n913 & ~n1081 ;
  assign n1593 = n736 | n1190 ;
  assign n1594 = ~n734 & n1190 ;
  assign n1595 = n1593 & ~n1594 ;
  assign n1596 = ~n1592 & n1595 ;
  assign n1597 = ~n1591 & n1596 ;
  assign n1598 = n1590 & n1597 ;
  assign n1599 = n1590 | n1597 ;
  assign n1600 = ~n1598 & n1599 ;
  assign n1601 = n906 & n1150 ;
  assign n1602 = n906 | n1099 ;
  assign n1603 = ~n782 & n1151 ;
  assign n1604 = n782 & n1097 ;
  assign n1605 = n1603 | n1604 ;
  assign n1606 = n1602 & ~n1605 ;
  assign n1607 = ~n1601 & n1606 ;
  assign n1608 = n1600 & n1607 ;
  assign n1609 = n1598 | n1608 ;
  assign n1610 = ~n1412 & n1609 ;
  assign n1611 = n1583 & n1610 ;
  assign n1612 = ~n1412 & n1583 ;
  assign n1613 = n1609 | n1612 ;
  assign n1614 = ( n1543 & n1558 ) | ( n1543 & ~n1559 ) | ( n1558 & ~n1559 );
  assign n1615 = ( n1549 & ~n1559 ) | ( n1549 & n1614 ) | ( ~n1559 & n1614 );
  assign n1616 = ~n1611 & n1615 ;
  assign n1617 = n1613 & n1616 ;
  assign n1618 = n1611 | n1617 ;
  assign n1619 = ~n1487 & n1488 ;
  assign n1620 = n1490 | n1619 ;
  assign n1621 = n1490 & n1619 ;
  assign n1622 = n1620 & ~n1621 ;
  assign n1623 = n1618 & ~n1622 ;
  assign n1624 = n1562 | n1564 ;
  assign n1625 = ~n1565 & n1624 ;
  assign n1626 = ~n1618 & n1622 ;
  assign n1627 = n1623 | n1626 ;
  assign n1628 = n1625 & ~n1627 ;
  assign n1629 = n1623 | n1628 ;
  assign n1630 = ~n1580 & n1629 ;
  assign n1631 = n1580 & ~n1629 ;
  assign n1632 = n1630 | n1631 ;
  assign n1633 = n1529 & ~n1535 ;
  assign n1634 = n1536 | n1633 ;
  assign n1635 = n1555 & ~n1557 ;
  assign n1636 = n1558 | n1635 ;
  assign n1637 = n725 & n1233 ;
  assign n1638 = n713 & ~n1233 ;
  assign n1639 = ( n552 & n1314 ) | ( n552 & ~n1638 ) | ( n1314 & ~n1638 );
  assign n1640 = ( ~n550 & n1314 ) | ( ~n550 & n1638 ) | ( n1314 & n1638 );
  assign n1641 = n1639 & ~n1640 ;
  assign n1642 = ~n1637 & n1641 ;
  assign n1643 = ~n1636 & n1642 ;
  assign n1644 = ~n700 & n1243 ;
  assign n1645 = n906 | n1241 ;
  assign n1646 = n700 & n1237 ;
  assign n1647 = n906 & ~n1239 ;
  assign n1648 = n1646 | n1647 ;
  assign n1649 = n1645 & ~n1648 ;
  assign n1650 = ~n1644 & n1649 ;
  assign n1651 = n375 & ~n1352 ;
  assign n1652 = ~n1024 & n1651 ;
  assign n1653 = n1024 & ~n1651 ;
  assign n1654 = n709 & n1352 ;
  assign n1655 = n1653 | n1654 ;
  assign n1656 = n1652 | n1655 ;
  assign n1657 = n1650 & ~n1656 ;
  assign n1658 = ~n1650 & n1656 ;
  assign n1659 = n1657 | n1658 ;
  assign n1660 = n782 & n1150 ;
  assign n1661 = n782 | n1099 ;
  assign n1662 = ~n1081 & n1151 ;
  assign n1663 = n1081 & n1097 ;
  assign n1664 = n1662 | n1663 ;
  assign n1665 = n1661 & ~n1664 ;
  assign n1666 = ~n1660 & n1665 ;
  assign n1667 = ~n1659 & n1666 ;
  assign n1668 = n1657 | n1667 ;
  assign n1669 = n1642 & ~n1643 ;
  assign n1670 = ( n1636 & n1643 ) | ( n1636 & ~n1669 ) | ( n1643 & ~n1669 );
  assign n1671 = n1668 & ~n1670 ;
  assign n1672 = n1643 | n1671 ;
  assign n1673 = ~n1634 & n1672 ;
  assign n1674 = ~n1611 & n1613 ;
  assign n1675 = n1615 | n1674 ;
  assign n1676 = n1634 & ~n1672 ;
  assign n1677 = n1673 | n1676 ;
  assign n1678 = n1617 | n1677 ;
  assign n1679 = n1675 & ~n1678 ;
  assign n1680 = n1673 | n1679 ;
  assign n1681 = ~n1625 & n1627 ;
  assign n1682 = n1628 | n1681 ;
  assign n1683 = n1680 & ~n1682 ;
  assign n1684 = ~n1680 & n1682 ;
  assign n1685 = ~n906 & n1243 ;
  assign n1686 = n782 | n1241 ;
  assign n1687 = n906 & n1237 ;
  assign n1688 = n782 & ~n1239 ;
  assign n1689 = n1687 | n1688 ;
  assign n1690 = n1686 & ~n1689 ;
  assign n1691 = ~n1685 & n1690 ;
  assign n1692 = n1081 & n1150 ;
  assign n1693 = n1081 | n1099 ;
  assign n1694 = n1151 & ~n1190 ;
  assign n1695 = n1097 & n1190 ;
  assign n1696 = n1694 | n1695 ;
  assign n1697 = n1693 & ~n1696 ;
  assign n1698 = ~n1692 & n1697 ;
  assign n1699 = n1691 & n1698 ;
  assign n1700 = n1691 | n1698 ;
  assign n1701 = ~n1699 & n1700 ;
  assign n1702 = n911 & n1233 ;
  assign n1703 = n913 & ~n1233 ;
  assign n1704 = n736 | n1314 ;
  assign n1705 = ~n734 & n1314 ;
  assign n1706 = n1704 & ~n1705 ;
  assign n1707 = ~n1703 & n1706 ;
  assign n1708 = ~n1702 & n1707 ;
  assign n1709 = n1701 & n1708 ;
  assign n1710 = n1699 | n1709 ;
  assign n1711 = n1659 & ~n1666 ;
  assign n1712 = n1667 | n1711 ;
  assign n1713 = n1710 & ~n1712 ;
  assign n1714 = n549 & n1314 ;
  assign n1715 = n692 | n1314 ;
  assign n1716 = n911 & n1314 ;
  assign n1717 = n736 & ~n1716 ;
  assign n1718 = n1715 & n1717 ;
  assign n1719 = n692 & n1718 ;
  assign n1720 = n709 & ~n1352 ;
  assign n1721 = ~n1024 & n1720 ;
  assign n1722 = n700 | n1024 ;
  assign n1723 = n1352 & n1722 ;
  assign n1724 = ~n709 & n1024 ;
  assign n1725 = n1723 | n1724 ;
  assign n1726 = n1721 | n1725 ;
  assign n1727 = n1719 & ~n1726 ;
  assign n1728 = n911 & n1190 ;
  assign n1729 = n913 & ~n1190 ;
  assign n1730 = n736 | n1233 ;
  assign n1731 = ~n734 & n1233 ;
  assign n1732 = n1730 & ~n1731 ;
  assign n1733 = ~n1729 & n1732 ;
  assign n1734 = ~n1728 & n1733 ;
  assign n1735 = n1727 & n1734 ;
  assign n1736 = n1727 | n1734 ;
  assign n1737 = ~n1735 & n1736 ;
  assign n1738 = n1714 & n1737 ;
  assign n1739 = n1714 | n1737 ;
  assign n1740 = ~n1738 & n1739 ;
  assign n1741 = ~n1710 & n1712 ;
  assign n1742 = n1713 | n1741 ;
  assign n1743 = n1740 & ~n1742 ;
  assign n1744 = n1713 | n1743 ;
  assign n1745 = n1735 | n1738 ;
  assign n1746 = n1600 | n1607 ;
  assign n1747 = ~n1608 & n1746 ;
  assign n1748 = n1745 & n1747 ;
  assign n1749 = n1745 | n1747 ;
  assign n1750 = ~n1748 & n1749 ;
  assign n1751 = ~n1668 & n1670 ;
  assign n1752 = n1671 | n1751 ;
  assign n1753 = ~n1750 & n1752 ;
  assign n1754 = n1750 & ~n1752 ;
  assign n1755 = n1753 | n1754 ;
  assign n1756 = ~n1744 & n1755 ;
  assign n1757 = n906 & n1352 ;
  assign n1758 = n700 & ~n1352 ;
  assign n1759 = ~n1024 & n1758 ;
  assign n1760 = n1024 & ~n1758 ;
  assign n1761 = n1759 | n1760 ;
  assign n1762 = n1757 | n1761 ;
  assign n1763 = n782 & n1237 ;
  assign n1764 = ~n782 & n1243 ;
  assign n1765 = n1081 | n1241 ;
  assign n1766 = n1081 & ~n1239 ;
  assign n1767 = n1765 & ~n1766 ;
  assign n1768 = ~n1764 & n1767 ;
  assign n1769 = ~n1763 & n1768 ;
  assign n1770 = ~n1762 & n1769 ;
  assign n1771 = n1762 & ~n1769 ;
  assign n1772 = n1770 | n1771 ;
  assign n1773 = n1150 & n1190 ;
  assign n1774 = n1099 | n1190 ;
  assign n1775 = n1151 & ~n1233 ;
  assign n1776 = n1097 & n1233 ;
  assign n1777 = n1775 | n1776 ;
  assign n1778 = n1774 & ~n1777 ;
  assign n1779 = ~n1773 & n1778 ;
  assign n1780 = ~n1772 & n1779 ;
  assign n1781 = n1770 | n1780 ;
  assign n1782 = ~n1719 & n1726 ;
  assign n1783 = n1727 | n1782 ;
  assign n1784 = n1781 & ~n1783 ;
  assign n1785 = ~n1781 & n1783 ;
  assign n1786 = n1784 | n1785 ;
  assign n1787 = n1701 | n1708 ;
  assign n1788 = ~n1709 & n1787 ;
  assign n1789 = ~n1786 & n1788 ;
  assign n1790 = n1784 | n1789 ;
  assign n1791 = ~n1740 & n1742 ;
  assign n1792 = n1743 | n1791 ;
  assign n1793 = ~n1790 & n1792 ;
  assign n1794 = n692 | n1718 ;
  assign n1795 = ~n1719 & n1794 ;
  assign n1796 = n782 | n1024 ;
  assign n1797 = n1352 & n1796 ;
  assign n1798 = n906 & n1024 ;
  assign n1799 = n906 | n1024 ;
  assign n1800 = ~n1352 & n1799 ;
  assign n1801 = ~n1798 & n1800 ;
  assign n1802 = n1797 | n1801 ;
  assign n1803 = n1150 & n1314 ;
  assign n1804 = n899 & ~n1803 ;
  assign n1805 = ~n1151 & n1804 ;
  assign n1806 = ~n1802 & n1805 ;
  assign n1807 = n1795 & n1806 ;
  assign n1808 = n1795 | n1806 ;
  assign n1809 = ~n1807 & n1808 ;
  assign n1810 = n1150 & n1233 ;
  assign n1811 = n1099 | n1233 ;
  assign n1812 = n1151 & ~n1314 ;
  assign n1813 = n1097 & n1314 ;
  assign n1814 = n1812 | n1813 ;
  assign n1815 = n1811 & ~n1814 ;
  assign n1816 = ~n1810 & n1815 ;
  assign n1817 = n1190 | n1241 ;
  assign n1818 = ~n1081 & n1243 ;
  assign n1819 = n1817 & ~n1818 ;
  assign n1820 = n1081 & n1237 ;
  assign n1821 = n1190 & ~n1239 ;
  assign n1822 = n1820 | n1821 ;
  assign n1823 = n1819 & ~n1822 ;
  assign n1824 = n1816 & n1823 ;
  assign n1825 = n1816 | n1823 ;
  assign n1826 = n1802 & ~n1805 ;
  assign n1827 = n1806 | n1826 ;
  assign n1828 = n1825 & ~n1827 ;
  assign n1829 = n1824 | n1828 ;
  assign n1830 = n1809 & n1829 ;
  assign n1831 = n1807 | n1830 ;
  assign n1832 = n1786 & ~n1788 ;
  assign n1833 = n1789 | n1832 ;
  assign n1834 = ~n1831 & n1833 ;
  assign n1835 = n1793 | n1834 ;
  assign n1836 = n1809 | n1829 ;
  assign n1837 = ~n1830 & n1836 ;
  assign n1838 = ~n1824 & n1825 ;
  assign n1839 = n1827 & n1838 ;
  assign n1840 = n1827 | n1838 ;
  assign n1841 = ~n1839 & n1840 ;
  assign n1842 = n1024 | n1081 ;
  assign n1843 = n1352 & n1842 ;
  assign n1844 = n782 & n1024 ;
  assign n1845 = n1796 & ~n1844 ;
  assign n1846 = ~n1352 & n1845 ;
  assign n1847 = n1843 | n1846 ;
  assign n1848 = n1233 | n1241 ;
  assign n1849 = n1233 & ~n1239 ;
  assign n1850 = n1848 & ~n1849 ;
  assign n1851 = n1190 & n1237 ;
  assign n1852 = ~n1190 & n1243 ;
  assign n1853 = n1851 | n1852 ;
  assign n1854 = n1850 & ~n1853 ;
  assign n1855 = ~n1847 & n1854 ;
  assign n1856 = n1195 & n1314 ;
  assign n1857 = n1077 & ~n1856 ;
  assign n1858 = n1024 | n1190 ;
  assign n1859 = n1352 & n1858 ;
  assign n1860 = n1024 & n1081 ;
  assign n1861 = n1352 | n1860 ;
  assign n1862 = n1842 & ~n1861 ;
  assign n1863 = n1859 | n1862 ;
  assign n1864 = n1857 & ~n1863 ;
  assign n1865 = n1847 & ~n1854 ;
  assign n1866 = n1855 | n1865 ;
  assign n1867 = n1864 & ~n1866 ;
  assign n1868 = n1855 | n1867 ;
  assign n1869 = n1841 & ~n1868 ;
  assign n1870 = ~n1841 & n1868 ;
  assign n1871 = ~n1857 & n1863 ;
  assign n1872 = n1864 | n1871 ;
  assign n1873 = n1190 & ~n1352 ;
  assign n1874 = n1024 & n1873 ;
  assign n1875 = n1233 & n1352 ;
  assign n1876 = n1024 | n1875 ;
  assign n1877 = n1873 | n1876 ;
  assign n1878 = ~n1874 & n1877 ;
  assign n1879 = n1233 & ~n1352 ;
  assign n1880 = n1314 | n1879 ;
  assign n1881 = n1873 | n1880 ;
  assign n1882 = ~n1856 & n1881 ;
  assign n1883 = n1878 | n1882 ;
  assign n1884 = n1872 & n1883 ;
  assign n1885 = n1872 | n1883 ;
  assign n1886 = n1241 | n1314 ;
  assign n1887 = ~n1233 & n1243 ;
  assign n1888 = n1233 & n1237 ;
  assign n1889 = ~n1239 & n1314 ;
  assign n1890 = n1888 | n1889 ;
  assign n1891 = n1887 | n1890 ;
  assign n1892 = n1886 & ~n1891 ;
  assign n1893 = n1885 & ~n1892 ;
  assign n1894 = n1884 | n1893 ;
  assign n1895 = ~n1096 & n1314 ;
  assign n1896 = ~n1894 & n1895 ;
  assign n1897 = n1870 | n1896 ;
  assign n1898 = n1894 & ~n1895 ;
  assign n1899 = ~n1864 & n1866 ;
  assign n1900 = n1867 | n1899 ;
  assign n1901 = n1898 | n1900 ;
  assign n1902 = ~n1897 & n1901 ;
  assign n1903 = n1869 | n1902 ;
  assign n1904 = n1837 & ~n1903 ;
  assign n1905 = n1831 & ~n1833 ;
  assign n1906 = ~n1837 & n1903 ;
  assign n1907 = n1772 & ~n1779 ;
  assign n1908 = n1780 | n1907 ;
  assign n1909 = n1906 | n1908 ;
  assign n1910 = ~n1905 & n1909 ;
  assign n1911 = ~n1904 & n1910 ;
  assign n1912 = n1835 | n1911 ;
  assign n1913 = n1744 & ~n1755 ;
  assign n1914 = n1790 & ~n1792 ;
  assign n1915 = n1913 | n1914 ;
  assign n1916 = n1912 & ~n1915 ;
  assign n1917 = n1756 | n1916 ;
  assign n1918 = n1748 | n1754 ;
  assign n1919 = n1917 & ~n1918 ;
  assign n1920 = ~n1917 & n1918 ;
  assign n1921 = ~n1617 & n1675 ;
  assign n1922 = n1677 & ~n1921 ;
  assign n1923 = n1679 | n1922 ;
  assign n1924 = ~n1920 & n1923 ;
  assign n1925 = n1919 | n1924 ;
  assign n1926 = n1684 | n1925 ;
  assign n1927 = ~n1683 & n1926 ;
  assign n1928 = n1632 | n1927 ;
  assign n1929 = ~n1630 & n1928 ;
  assign n1930 = ~n1575 & n1577 ;
  assign n1931 = n1578 | n1930 ;
  assign n1932 = n1929 | n1931 ;
  assign n1933 = ~n1578 & n1932 ;
  assign n1934 = n1513 | n1933 ;
  assign n1935 = ~n1511 & n1934 ;
  assign n1936 = n1401 | n1407 ;
  assign n1937 = ~n1468 & n1936 ;
  assign n1938 = n1470 | n1937 ;
  assign n1939 = n1935 | n1938 ;
  assign n1940 = ~n1470 & n1939 ;
  assign n1941 = ~n1402 & n1404 ;
  assign n1942 = n1405 | n1941 ;
  assign n1943 = n1940 | n1942 ;
  assign n1944 = ~n1405 & n1943 ;
  assign n1945 = ~n1292 & n1294 ;
  assign n1946 = n1295 | n1945 ;
  assign n1947 = n1944 | n1946 ;
  assign n1948 = ~n1295 & n1947 ;
  assign n1949 = ~n1172 & n1174 ;
  assign n1950 = n1175 | n1949 ;
  assign n1951 = n1948 | n1950 ;
  assign n1952 = ~n1175 & n1951 ;
  assign n1953 = ~n1128 & n1131 ;
  assign n1954 = n1132 | n1953 ;
  assign n1955 = n1952 | n1954 ;
  assign n1956 = ~n1132 & n1955 ;
  assign n1957 = n954 | n1956 ;
  assign n1958 = ~n952 & n1957 ;
  assign n1959 = n767 | n1958 ;
  assign n1960 = ~n765 & n1959 ;
  assign n1961 = ~n584 & n586 ;
  assign n1962 = n587 | n1961 ;
  assign n1963 = n1960 | n1962 ;
  assign n1964 = ~n587 & n1963 ;
  assign n1965 = n47 | n224 ;
  assign n1966 = n47 & n224 ;
  assign n1967 = n1965 & ~n1966 ;
  assign n1968 = n352 & ~n1967 ;
  assign n1969 = ~n352 & n1967 ;
  assign n1970 = n1968 | n1969 ;
  assign n1971 = n219 & ~n1970 ;
  assign n1972 = ~n1964 & n1971 ;
  assign n1973 = n587 | n1971 ;
  assign n1974 = n1963 & ~n1973 ;
  assign n1975 = n1972 | n1974 ;
  assign n1976 = ~n544 & n1975 ;
  assign n1977 = n544 & ~n1974 ;
  assign n1978 = ~n1972 & n1977 ;
  assign n1979 = n1976 | n1978 ;
  assign n1980 = n115 | n622 ;
  assign n1981 = n145 | n232 ;
  assign n1982 = n263 | n1981 ;
  assign n1983 = n393 | n1027 ;
  assign n1984 = n1982 | n1983 ;
  assign n1985 = n273 | n462 ;
  assign n1986 = n180 | n1985 ;
  assign n1987 = n195 | n1986 ;
  assign n1988 = n296 | n1987 ;
  assign n1989 = n1984 | n1988 ;
  assign n1990 = n227 | n1989 ;
  assign n1991 = n176 | n403 ;
  assign n1992 = n1990 | n1991 ;
  assign n1993 = n192 | n1992 ;
  assign n1994 = n295 | n1993 ;
  assign n1995 = n146 | n654 ;
  assign n1996 = n1994 | n1995 ;
  assign n1997 = n1980 | n1996 ;
  assign n1998 = n422 | n1997 ;
  assign n1999 = n201 | n401 ;
  assign n2000 = n135 | n257 ;
  assign n2001 = n448 | n2000 ;
  assign n2002 = n229 | n2001 ;
  assign n2003 = n1999 | n2002 ;
  assign n2004 = n185 | n196 ;
  assign n2005 = n152 | n2004 ;
  assign n2006 = n321 | n2005 ;
  assign n2007 = n117 | n2006 ;
  assign n2008 = n2003 | n2007 ;
  assign n2009 = n1998 | n2008 ;
  assign n2010 = ~n810 & n828 ;
  assign n2011 = n165 | n207 ;
  assign n2012 = n2010 & ~n2011 ;
  assign n2013 = ~n2009 & n2012 ;
  assign n2014 = ~n991 & n2013 ;
  assign n2015 = n1979 & n2014 ;
  assign n2016 = n1960 & n1962 ;
  assign n2017 = n1963 & ~n2016 ;
  assign n2018 = n165 | n268 ;
  assign n2019 = n140 | n2018 ;
  assign n2020 = n194 | n335 ;
  assign n2021 = n2019 | n2020 ;
  assign n2022 = n256 | n448 ;
  assign n2023 = n157 | n186 ;
  assign n2024 = n282 | n401 ;
  assign n2025 = n251 | n318 ;
  assign n2026 = n257 | n2025 ;
  assign n2027 = n2024 | n2026 ;
  assign n2028 = n190 | n2027 ;
  assign n2029 = n2023 | n2028 ;
  assign n2030 = n316 | n483 ;
  assign n2031 = n271 | n663 ;
  assign n2032 = n2030 | n2031 ;
  assign n2033 = n2029 | n2032 ;
  assign n2034 = n588 | n2033 ;
  assign n2035 = n328 | n447 ;
  assign n2036 = n403 | n2035 ;
  assign n2037 = n137 | n386 ;
  assign n2038 = n243 | n2037 ;
  assign n2039 = n275 | n2038 ;
  assign n2040 = n250 | n504 ;
  assign n2041 = n115 | n329 ;
  assign n2042 = n473 | n2041 ;
  assign n2043 = n870 | n972 ;
  assign n2044 = n2042 | n2043 ;
  assign n2045 = n2040 | n2044 ;
  assign n2046 = n2039 | n2045 ;
  assign n2047 = n2036 | n2046 ;
  assign n2048 = n2034 | n2047 ;
  assign n2049 = n312 | n330 ;
  assign n2050 = n128 | n291 ;
  assign n2051 = n2049 | n2050 ;
  assign n2052 = n209 | n598 ;
  assign n2053 = n293 | n2052 ;
  assign n2054 = n151 | n2053 ;
  assign n2055 = n2051 | n2054 ;
  assign n2056 = n499 | n2055 ;
  assign n2057 = n149 | n617 ;
  assign n2058 = n202 | n2057 ;
  assign n2059 = n2056 | n2058 ;
  assign n2060 = n683 | n2059 ;
  assign n2061 = n2048 | n2060 ;
  assign n2062 = n2022 | n2061 ;
  assign n2063 = n2021 | n2062 ;
  assign n2064 = n263 | n392 ;
  assign n2065 = n2063 | n2064 ;
  assign n2066 = ~n2017 & n2065 ;
  assign n2067 = n767 & n1958 ;
  assign n2068 = n1959 & ~n2067 ;
  assign n2069 = n513 | n983 ;
  assign n2070 = n275 | n318 ;
  assign n2071 = n2069 | n2070 ;
  assign n2072 = n434 | n638 ;
  assign n2073 = n592 | n813 ;
  assign n2074 = n806 | n2073 ;
  assign n2075 = n244 | n2074 ;
  assign n2076 = n2072 | n2075 ;
  assign n2077 = n856 | n2076 ;
  assign n2078 = n398 | n2077 ;
  assign n2079 = n229 | n2078 ;
  assign n2080 = n291 | n2079 ;
  assign n2081 = n2071 | n2080 ;
  assign n2082 = ~n2068 & n2081 ;
  assign n2083 = n954 & n1956 ;
  assign n2084 = n1957 & ~n2083 ;
  assign n2085 = n204 | n316 ;
  assign n2086 = n240 | n313 ;
  assign n2087 = n621 | n2086 ;
  assign n2088 = n142 | n399 ;
  assign n2089 = n462 | n2088 ;
  assign n2090 = n2087 | n2089 ;
  assign n2091 = n434 | n2019 ;
  assign n2092 = n2001 | n2042 ;
  assign n2093 = n2091 | n2092 ;
  assign n2094 = n2090 | n2093 ;
  assign n2095 = n2085 | n2094 ;
  assign n2096 = n239 | n331 ;
  assign n2097 = n181 | n2096 ;
  assign n2098 = n381 | n2097 ;
  assign n2099 = n253 | n1991 ;
  assign n2100 = n2098 | n2099 ;
  assign n2101 = n282 | n812 ;
  assign n2102 = n270 | n312 ;
  assign n2103 = n2101 | n2102 ;
  assign n2104 = n503 | n2103 ;
  assign n2105 = n269 | n2104 ;
  assign n2106 = n488 | n636 ;
  assign n2107 = n2105 | n2106 ;
  assign n2108 = n158 | n179 ;
  assign n2109 = n388 | n2108 ;
  assign n2110 = n2107 | n2109 ;
  assign n2111 = n117 | n389 ;
  assign n2112 = n405 | n2111 ;
  assign n2113 = n2110 | n2112 ;
  assign n2114 = n205 | n234 ;
  assign n2115 = n334 | n2114 ;
  assign n2116 = n494 | n2115 ;
  assign n2117 = n2113 | n2116 ;
  assign n2118 = n2100 | n2117 ;
  assign n2119 = n2095 | n2118 ;
  assign n2120 = ~n2084 & n2119 ;
  assign n2121 = n2084 & ~n2119 ;
  assign n2122 = n2120 | n2121 ;
  assign n2123 = n113 & n139 ;
  assign n2124 = n190 | n205 ;
  assign n2125 = n168 | n862 ;
  assign n2126 = n270 | n513 ;
  assign n2127 = n377 | n2126 ;
  assign n2128 = n2125 | n2127 ;
  assign n2129 = n197 | n278 ;
  assign n2130 = n2097 | n2129 ;
  assign n2131 = n413 | n2130 ;
  assign n2132 = n208 | n2131 ;
  assign n2133 = n314 | n321 ;
  assign n2134 = n263 | n2133 ;
  assign n2135 = n2132 | n2134 ;
  assign n2136 = n383 | n2135 ;
  assign n2137 = n2056 | n2136 ;
  assign n2138 = n233 | n392 ;
  assign n2139 = n148 | n2138 ;
  assign n2140 = n2095 | n2139 ;
  assign n2141 = n828 & ~n2140 ;
  assign n2142 = ~n1322 & n2141 ;
  assign n2143 = ~n2137 & n2142 ;
  assign n2144 = ~n2128 & n2143 ;
  assign n2145 = ~n2124 & n2144 ;
  assign n2146 = ~n2123 & n2145 ;
  assign n2147 = ~n1175 & n1954 ;
  assign n2148 = n1951 & n2147 ;
  assign n2149 = n1955 & ~n2148 ;
  assign n2150 = n2146 | n2149 ;
  assign n2151 = n177 | n277 ;
  assign n2152 = n234 | n2151 ;
  assign n2153 = n140 | n448 ;
  assign n2154 = n179 | n313 ;
  assign n2155 = n122 | n2154 ;
  assign n2156 = n164 | n330 ;
  assign n2157 = n2155 | n2156 ;
  assign n2158 = n246 | n2157 ;
  assign n2159 = n229 | n336 ;
  assign n2160 = n2158 | n2159 ;
  assign n2161 = n194 | n230 ;
  assign n2162 = n273 | n382 ;
  assign n2163 = n248 | n2162 ;
  assign n2164 = n2161 | n2163 ;
  assign n2165 = n255 | n826 ;
  assign n2166 = n401 | n2165 ;
  assign n2167 = n196 | n1981 ;
  assign n2168 = n210 | n381 ;
  assign n2169 = n1009 | n2168 ;
  assign n2170 = n2167 | n2169 ;
  assign n2171 = n843 | n2170 ;
  assign n2172 = n291 | n2171 ;
  assign n2173 = n270 | n293 ;
  assign n2174 = n2172 | n2173 ;
  assign n2175 = n2166 | n2174 ;
  assign n2176 = n2164 | n2175 ;
  assign n2177 = n2160 | n2176 ;
  assign n2178 = n129 | n2177 ;
  assign n2179 = n2153 | n2178 ;
  assign n2180 = n328 | n2179 ;
  assign n2181 = n2152 | n2180 ;
  assign n2182 = n1948 & n1950 ;
  assign n2183 = n1951 & ~n2182 ;
  assign n2184 = n2181 & ~n2183 ;
  assign n2185 = n148 | n168 ;
  assign n2186 = n186 | n654 ;
  assign n2187 = n2185 | n2186 ;
  assign n2188 = n342 | n401 ;
  assign n2189 = n230 | n341 ;
  assign n2190 = n793 | n816 ;
  assign n2191 = n672 | n2190 ;
  assign n2192 = n2189 | n2191 ;
  assign n2193 = n2188 | n2192 ;
  assign n2194 = n122 | n273 ;
  assign n2195 = n255 | n294 ;
  assign n2196 = n503 | n2195 ;
  assign n2197 = n178 | n2196 ;
  assign n2198 = n2194 | n2197 ;
  assign n2199 = n206 | n422 ;
  assign n2200 = n2198 | n2199 ;
  assign n2201 = n1035 | n2200 ;
  assign n2202 = n2193 | n2201 ;
  assign n2203 = n263 | n2202 ;
  assign n2204 = n246 | n790 ;
  assign n2205 = n2203 | n2204 ;
  assign n2206 = n2187 | n2205 ;
  assign n2207 = n304 | n588 ;
  assign n2208 = n274 | n865 ;
  assign n2209 = n124 | n2208 ;
  assign n2210 = n2207 | n2209 ;
  assign n2211 = n444 | n786 ;
  assign n2212 = n227 | n448 ;
  assign n2213 = n2211 | n2212 ;
  assign n2214 = n333 | n336 ;
  assign n2215 = n483 | n870 ;
  assign n2216 = n2214 | n2215 ;
  assign n2217 = n2213 | n2216 ;
  assign n2218 = n2210 | n2217 ;
  assign n2219 = n2206 | n2218 ;
  assign n2220 = n248 | n2219 ;
  assign n2221 = n317 | n2220 ;
  assign n2222 = n1944 & n1946 ;
  assign n2223 = n1947 & ~n2222 ;
  assign n2224 = n2221 & ~n2223 ;
  assign n2225 = n190 | n433 ;
  assign n2226 = n293 | n2225 ;
  assign n2227 = n201 | n389 ;
  assign n2228 = n177 | n513 ;
  assign n2229 = n503 | n2228 ;
  assign n2230 = n2227 | n2229 ;
  assign n2231 = n233 | n276 ;
  assign n2232 = n135 | n2231 ;
  assign n2233 = n377 | n2232 ;
  assign n2234 = n2230 | n2233 ;
  assign n2235 = n152 | n343 ;
  assign n2236 = n247 | n294 ;
  assign n2237 = n257 | n2236 ;
  assign n2238 = n814 | n2237 ;
  assign n2239 = n2235 | n2238 ;
  assign n2240 = n272 | n2035 ;
  assign n2241 = n1993 | n2240 ;
  assign n2242 = n2239 | n2241 ;
  assign n2243 = n2234 | n2242 ;
  assign n2244 = n184 | n210 ;
  assign n2245 = n158 | n2244 ;
  assign n2246 = n205 | n281 ;
  assign n2247 = n499 | n2246 ;
  assign n2248 = n2245 | n2247 ;
  assign n2249 = n240 | n2248 ;
  assign n2250 = n204 | n399 ;
  assign n2251 = n2249 | n2250 ;
  assign n2252 = n2243 | n2251 ;
  assign n2253 = n2226 | n2252 ;
  assign n2254 = n264 | n2253 ;
  assign n2255 = n1940 & n1942 ;
  assign n2256 = n1943 & ~n2255 ;
  assign n2257 = n2254 & ~n2256 ;
  assign n2258 = n389 | n622 ;
  assign n2259 = n251 | n2258 ;
  assign n2260 = n140 | n313 ;
  assign n2261 = n870 | n2260 ;
  assign n2262 = n466 | n2261 ;
  assign n2263 = n2259 | n2262 ;
  assign n2264 = n263 | n281 ;
  assign n2265 = n138 | n258 ;
  assign n2266 = n320 | n2265 ;
  assign n2267 = n328 | n2266 ;
  assign n2268 = n2264 | n2267 ;
  assign n2269 = n484 | n2268 ;
  assign n2270 = n812 | n2115 ;
  assign n2271 = n517 | n2270 ;
  assign n2272 = n131 | n2271 ;
  assign n2273 = n297 | n2272 ;
  assign n2274 = n227 | n2273 ;
  assign n2275 = n2188 | n2274 ;
  assign n2276 = n2269 | n2275 ;
  assign n2277 = n641 | n2276 ;
  assign n2278 = n186 | n648 ;
  assign n2279 = n117 | n635 ;
  assign n2280 = n2278 | n2279 ;
  assign n2281 = n2277 | n2280 ;
  assign n2282 = n2263 | n2281 ;
  assign n2283 = n233 | n2282 ;
  assign n2284 = n194 | n2283 ;
  assign n2285 = n1935 & n1938 ;
  assign n2286 = n1939 & ~n2285 ;
  assign n2287 = n2284 & ~n2286 ;
  assign n2288 = n393 | n2127 ;
  assign n2289 = n252 | n321 ;
  assign n2290 = n269 | n1319 ;
  assign n2291 = n2289 | n2290 ;
  assign n2292 = n885 | n2291 ;
  assign n2293 = n2231 | n2292 ;
  assign n2294 = n2288 | n2293 ;
  assign n2295 = n264 | n2294 ;
  assign n2296 = n304 | n333 ;
  assign n2297 = n588 | n654 ;
  assign n2298 = n2296 | n2297 ;
  assign n2299 = n2295 | n2298 ;
  assign n2300 = n318 | n790 ;
  assign n2301 = n227 | n2300 ;
  assign n2302 = n314 | n2301 ;
  assign n2303 = n2299 | n2302 ;
  assign n2304 = n335 | n400 ;
  assign n2305 = n197 | n2304 ;
  assign n2306 = n618 | n2305 ;
  assign n2307 = n2268 | n2306 ;
  assign n2308 = n2010 & ~n2307 ;
  assign n2309 = ~n477 & n2308 ;
  assign n2310 = ~n865 & n2309 ;
  assign n2311 = ~n2303 & n2310 ;
  assign n2312 = ~n448 & n2311 ;
  assign n2313 = ~n115 & n2312 ;
  assign n2314 = ~n1014 & n2313 ;
  assign n2315 = ~n503 & n2314 ;
  assign n2316 = n1513 & n1933 ;
  assign n2317 = n1934 & ~n2316 ;
  assign n2318 = n2315 | n2317 ;
  assign n2319 = n191 | n281 ;
  assign n2320 = n234 | n2319 ;
  assign n2321 = n377 | n403 ;
  assign n2322 = n444 | n2231 ;
  assign n2323 = n244 | n2322 ;
  assign n2324 = n184 | n329 ;
  assign n2325 = n296 | n2324 ;
  assign n2326 = n168 | n2325 ;
  assign n2327 = n447 | n2326 ;
  assign n2328 = n293 | n389 ;
  assign n2329 = n2327 | n2328 ;
  assign n2330 = n2323 | n2329 ;
  assign n2331 = n148 | n179 ;
  assign n2332 = n1010 | n2331 ;
  assign n2333 = n286 | n291 ;
  assign n2334 = n314 | n2333 ;
  assign n2335 = n2193 | n2334 ;
  assign n2336 = n2332 | n2335 ;
  assign n2337 = n2330 | n2336 ;
  assign n2338 = n2321 | n2337 ;
  assign n2339 = n166 | n2338 ;
  assign n2340 = n207 | n2339 ;
  assign n2341 = n615 | n2340 ;
  assign n2342 = n330 | n2341 ;
  assign n2343 = n2320 | n2342 ;
  assign n2344 = n196 | n2343 ;
  assign n2345 = n1929 & n1931 ;
  assign n2346 = n1932 & ~n2345 ;
  assign n2347 = n2344 & ~n2346 ;
  assign n2348 = n158 | n2047 ;
  assign n2349 = n393 | n803 ;
  assign n2350 = n652 | n975 ;
  assign n2351 = n2349 | n2350 ;
  assign n2352 = n2348 | n2351 ;
  assign n2353 = n638 | n2275 ;
  assign n2354 = n271 | n318 ;
  assign n2355 = n191 | n2354 ;
  assign n2356 = n2353 | n2355 ;
  assign n2357 = n2352 | n2356 ;
  assign n2358 = n383 | n2357 ;
  assign n2359 = n1632 & n1927 ;
  assign n2360 = n1928 & ~n2359 ;
  assign n2361 = ~n2358 & n2360 ;
  assign n2362 = ~n2344 & n2346 ;
  assign n2363 = n2347 | n2362 ;
  assign n2364 = n2361 | n2363 ;
  assign n2365 = ~n2347 & n2364 ;
  assign n2366 = n2315 & n2317 ;
  assign n2367 = n2318 & ~n2366 ;
  assign n2368 = ~n2365 & n2367 ;
  assign n2369 = n2318 & ~n2368 ;
  assign n2370 = ~n2284 & n2286 ;
  assign n2371 = n2287 | n2370 ;
  assign n2372 = n2369 | n2371 ;
  assign n2373 = ~n2287 & n2372 ;
  assign n2374 = ~n2254 & n2256 ;
  assign n2375 = n2257 | n2374 ;
  assign n2376 = n2373 | n2375 ;
  assign n2377 = ~n2257 & n2376 ;
  assign n2378 = ~n2221 & n2223 ;
  assign n2379 = n2224 | n2378 ;
  assign n2380 = n2377 | n2379 ;
  assign n2381 = ~n2224 & n2380 ;
  assign n2382 = ~n2181 & n2183 ;
  assign n2383 = n2184 | n2382 ;
  assign n2384 = n2381 | n2383 ;
  assign n2385 = ~n2184 & n2384 ;
  assign n2386 = n2146 & n2149 ;
  assign n2387 = n2150 & ~n2386 ;
  assign n2388 = ~n2385 & n2387 ;
  assign n2389 = n2150 & ~n2388 ;
  assign n2390 = n2122 | n2389 ;
  assign n2391 = ~n2120 & n2390 ;
  assign n2392 = n2068 & ~n2081 ;
  assign n2393 = n2082 | n2392 ;
  assign n2394 = n2391 | n2393 ;
  assign n2395 = ~n2082 & n2394 ;
  assign n2396 = n2017 & ~n2065 ;
  assign n2397 = n2066 | n2396 ;
  assign n2398 = n2395 | n2397 ;
  assign n2399 = ~n2066 & n2398 ;
  assign n2400 = n1978 | n2014 ;
  assign n2401 = n1976 | n2400 ;
  assign n2402 = ~n2399 & n2401 ;
  assign n2403 = ~n2015 & n2402 ;
  assign n2404 = n152 | n165 ;
  assign n2405 = n179 | n195 ;
  assign n2406 = n2404 | n2405 ;
  assign n2407 = n181 | n284 ;
  assign n2408 = n129 | n2407 ;
  assign n2409 = n232 | n2408 ;
  assign n2410 = n2406 | n2409 ;
  assign n2411 = n253 | n972 ;
  assign n2412 = n2193 | n2411 ;
  assign n2413 = n2410 | n2412 ;
  assign n2414 = n1331 | n2413 ;
  assign n2415 = n466 | n2414 ;
  assign n2416 = n453 | n2415 ;
  assign n2417 = n829 | n2416 ;
  assign n2418 = n389 | n2417 ;
  assign n2419 = n1056 | n2418 ;
  assign n2420 = n227 | n2419 ;
  assign n2421 = n2401 & ~n2420 ;
  assign n2422 = ~n2403 & n2421 ;
  assign n2423 = n151 | n168 ;
  assign n2424 = n377 | n664 ;
  assign n2425 = n671 | n2424 ;
  assign n2426 = n2423 | n2425 ;
  assign n2427 = n179 | n665 ;
  assign n2428 = n115 | n2427 ;
  assign n2429 = n318 | n342 ;
  assign n2430 = n296 | n2429 ;
  assign n2431 = n290 | n401 ;
  assign n2432 = n617 | n2431 ;
  assign n2433 = n137 | n186 ;
  assign n2434 = n191 | n2019 ;
  assign n2435 = n247 | n271 ;
  assign n2436 = n177 | n433 ;
  assign n2437 = n2435 | n2436 ;
  assign n2438 = n2434 | n2437 ;
  assign n2439 = n2433 | n2438 ;
  assign n2440 = n2432 | n2439 ;
  assign n2441 = n304 | n2440 ;
  assign n2442 = n321 | n2441 ;
  assign n2443 = n270 | n2442 ;
  assign n2444 = n2430 | n2443 ;
  assign n2445 = n207 | n316 ;
  assign n2446 = n646 | n2445 ;
  assign n2447 = n2444 | n2446 ;
  assign n2448 = n2428 | n2447 ;
  assign n2449 = n135 | n389 ;
  assign n2450 = n276 | n2449 ;
  assign n2451 = n192 | n2450 ;
  assign n2452 = n256 | n447 ;
  assign n2453 = n2451 | n2452 ;
  assign n2454 = n152 | n240 ;
  assign n2455 = n157 | n285 ;
  assign n2456 = n2454 | n2455 ;
  assign n2457 = n2453 | n2456 ;
  assign n2458 = n194 | n403 ;
  assign n2459 = n122 | n294 ;
  assign n2460 = n2458 | n2459 ;
  assign n2461 = n200 | n251 ;
  assign n2462 = n176 | n255 ;
  assign n2463 = n2461 | n2462 ;
  assign n2464 = n2460 | n2463 ;
  assign n2465 = n2457 | n2464 ;
  assign n2466 = n2448 | n2465 ;
  assign n2467 = n2426 | n2466 ;
  assign n2468 = n329 | n2467 ;
  assign n2469 = n124 | n146 ;
  assign n2470 = n252 | n305 ;
  assign n2471 = n2469 | n2470 ;
  assign n2472 = n2468 | n2471 ;
  assign n2473 = n2422 & ~n2472 ;
  assign n2474 = n858 | n1319 ;
  assign n2475 = ~n623 & n827 ;
  assign n2476 = n175 | n266 ;
  assign n2477 = n2475 & ~n2476 ;
  assign n2478 = ~n2105 & n2477 ;
  assign n2479 = ~n275 & n2478 ;
  assign n2480 = ~n335 & n2479 ;
  assign n2481 = ~n2474 & n2480 ;
  assign n2482 = ~n2298 & n2481 ;
  assign n2483 = ~n284 & n2482 ;
  assign n2484 = ~n513 & n2483 ;
  assign n2485 = ~n622 & n2484 ;
  assign n2486 = n2473 & n2485 ;
  assign n2487 = n121 | n165 ;
  assign n2488 = n280 | n2487 ;
  assign n2489 = n295 | n1048 ;
  assign n2490 = n160 | n2489 ;
  assign n2491 = n2488 | n2490 ;
  assign n2492 = n189 | n202 ;
  assign n2493 = n206 | n327 ;
  assign n2494 = n266 | n2493 ;
  assign n2495 = n2492 | n2494 ;
  assign n2496 = n2491 | n2495 ;
  assign n2497 = n209 | n2496 ;
  assign n2498 = n2486 & ~n2497 ;
  assign n2499 = n152 | n312 ;
  assign n2500 = n294 | n2499 ;
  assign n2501 = n346 | n2500 ;
  assign n2502 = n140 | n281 ;
  assign n2503 = n133 | n327 ;
  assign n2504 = n164 | n215 ;
  assign n2505 = n266 | n2504 ;
  assign n2506 = n2503 | n2505 ;
  assign n2507 = n2502 | n2506 ;
  assign n2508 = n2501 | n2507 ;
  assign n2509 = ~n2498 & n2508 ;
  assign n2510 = n2498 & ~n2508 ;
  assign n2511 = n2509 | n2510 ;
  assign n2512 = pi1 & ~n26 ;
  assign n2513 = ~pi1 & n26 ;
  assign n2514 = n2512 | n2513 ;
  assign n2515 = n32 & ~n2514 ;
  assign n2516 = ~n32 & n2514 ;
  assign n2517 = n2515 | n2516 ;
  assign n2518 = pi0 & ~n2517 ;
  assign n2519 = n2511 & n2518 ;
  assign n2520 = n2473 | n2485 ;
  assign n2521 = ~n2486 & n2520 ;
  assign n2522 = ~n29 & n2517 ;
  assign n2523 = ~n2521 & n2522 ;
  assign n2524 = n2486 | n2497 ;
  assign n2525 = n2486 & n2497 ;
  assign n2526 = n2524 & ~n2525 ;
  assign n2527 = ~pi0 & n2514 ;
  assign n2528 = n2526 & n2527 ;
  assign n2529 = n2523 | n2528 ;
  assign n2530 = n2519 | n2529 ;
  assign n2531 = pi0 & n2517 ;
  assign n2532 = n2511 | n2526 ;
  assign n2533 = n2511 & n2526 ;
  assign n2534 = n2532 & ~n2533 ;
  assign n2535 = n2521 & ~n2526 ;
  assign n2536 = n2401 & ~n2403 ;
  assign n2537 = n2420 & ~n2536 ;
  assign n2538 = n2422 | n2537 ;
  assign n2539 = ~n2015 & n2401 ;
  assign n2540 = n2399 & ~n2539 ;
  assign n2541 = n2403 | n2540 ;
  assign n2542 = n2538 & ~n2541 ;
  assign n2543 = n2395 & n2397 ;
  assign n2544 = n2398 & ~n2543 ;
  assign n2545 = ~n2541 & n2544 ;
  assign n2546 = n2541 & ~n2544 ;
  assign n2547 = n2545 | n2546 ;
  assign n2548 = n2391 & n2393 ;
  assign n2549 = n2394 & ~n2548 ;
  assign n2550 = n2544 & n2549 ;
  assign n2551 = n2122 & n2389 ;
  assign n2552 = n2390 & ~n2551 ;
  assign n2553 = n2549 & n2552 ;
  assign n2554 = n2385 & ~n2387 ;
  assign n2555 = n2388 | n2554 ;
  assign n2556 = n2552 & ~n2555 ;
  assign n2557 = n2381 & n2383 ;
  assign n2558 = n2384 & ~n2557 ;
  assign n2559 = ~n2555 & n2558 ;
  assign n2560 = n2377 & n2379 ;
  assign n2561 = n2380 & ~n2560 ;
  assign n2562 = n2558 & n2561 ;
  assign n2563 = n2558 | n2561 ;
  assign n2564 = ~n2562 & n2563 ;
  assign n2565 = n2373 & n2375 ;
  assign n2566 = n2376 & ~n2565 ;
  assign n2567 = n2561 & n2566 ;
  assign n2568 = n2369 & n2371 ;
  assign n2569 = n2372 & ~n2568 ;
  assign n2570 = n2566 & n2569 ;
  assign n2571 = n2365 & ~n2367 ;
  assign n2572 = n2368 | n2571 ;
  assign n2573 = n2569 & ~n2572 ;
  assign n2574 = ~n2569 & n2572 ;
  assign n2575 = n2361 & n2363 ;
  assign n2576 = n2364 & ~n2575 ;
  assign n2577 = n2358 & ~n2360 ;
  assign n2578 = n2361 | n2577 ;
  assign n2579 = n2572 & ~n2578 ;
  assign n2580 = n2576 & ~n2579 ;
  assign n2581 = ~n2574 & n2580 ;
  assign n2582 = ~n2573 & n2581 ;
  assign n2583 = n2573 | n2582 ;
  assign n2584 = n2566 | n2569 ;
  assign n2585 = n2583 & n2584 ;
  assign n2586 = ~n2570 & n2585 ;
  assign n2587 = n2570 | n2586 ;
  assign n2588 = n2561 | n2566 ;
  assign n2589 = ~n2567 & n2588 ;
  assign n2590 = n2587 & n2589 ;
  assign n2591 = n2567 | n2590 ;
  assign n2592 = n2564 & n2591 ;
  assign n2593 = n2562 | n2592 ;
  assign n2594 = n2555 & ~n2558 ;
  assign n2595 = n2559 | n2594 ;
  assign n2596 = n2593 & ~n2595 ;
  assign n2597 = n2559 | n2596 ;
  assign n2598 = ~n2552 & n2555 ;
  assign n2599 = n2556 | n2598 ;
  assign n2600 = n2597 & ~n2599 ;
  assign n2601 = n2556 | n2600 ;
  assign n2602 = n2549 | n2552 ;
  assign n2603 = ~n2553 & n2602 ;
  assign n2604 = n2601 & n2603 ;
  assign n2605 = n2553 | n2604 ;
  assign n2606 = n2544 | n2549 ;
  assign n2607 = ~n2550 & n2606 ;
  assign n2608 = n2605 & n2607 ;
  assign n2609 = n2550 | n2608 ;
  assign n2610 = n2545 | n2609 ;
  assign n2611 = ( n2545 & ~n2547 ) | ( n2545 & n2610 ) | ( ~n2547 & n2610 );
  assign n2612 = ~n2538 & n2541 ;
  assign n2613 = n2542 | n2612 ;
  assign n2614 = ~n2542 & n2613 ;
  assign n2615 = ( n2542 & n2611 ) | ( n2542 & ~n2614 ) | ( n2611 & ~n2614 );
  assign n2616 = n2422 | n2472 ;
  assign n2617 = n2422 & n2472 ;
  assign n2618 = n2616 & ~n2617 ;
  assign n2619 = ~n2521 & n2618 ;
  assign n2620 = n2521 & ~n2618 ;
  assign n2621 = n2619 | n2620 ;
  assign n2622 = n2538 & n2618 ;
  assign n2623 = n2538 | n2618 ;
  assign n2624 = ~n2622 & n2623 ;
  assign n2625 = n2622 | n2624 ;
  assign n2626 = ~n2621 & n2625 ;
  assign n2627 = ~n2621 & n2622 ;
  assign n2628 = ( n2615 & n2626 ) | ( n2615 & n2627 ) | ( n2626 & n2627 );
  assign n2629 = ( ~n2521 & n2526 ) | ( ~n2521 & n2619 ) | ( n2526 & n2619 );
  assign n2630 = ( ~n2535 & n2628 ) | ( ~n2535 & n2629 ) | ( n2628 & n2629 );
  assign n2631 = n2534 | n2630 ;
  assign n2632 = n2534 & n2629 ;
  assign n2633 = n2534 & ~n2535 ;
  assign n2634 = ( n2628 & n2632 ) | ( n2628 & n2633 ) | ( n2632 & n2633 );
  assign n2635 = n2631 & ~n2634 ;
  assign n2636 = n2531 & n2635 ;
  assign n2637 = n2530 | n2636 ;
  assign n2638 = n32 | n2637 ;
  assign n2639 = n32 & n2637 ;
  assign n2640 = n2638 & ~n2639 ;
  assign n2641 = ~n375 & n537 ;
  assign n2642 = n375 & ~n537 ;
  assign n2643 = n2641 | n2642 ;
  assign n2644 = n2578 & n2643 ;
  assign n2645 = n224 & ~n2644 ;
  assign n2646 = ~n47 & n537 ;
  assign n2647 = n47 & ~n537 ;
  assign n2648 = n2646 | n2647 ;
  assign n2649 = ~n2643 & n2648 ;
  assign n2650 = n2578 & n2649 ;
  assign n2651 = ~n1967 & n2643 ;
  assign n2652 = n2576 & n2651 ;
  assign n2653 = n2650 | n2652 ;
  assign n2654 = ~n2576 & n2578 ;
  assign n2655 = n2576 & ~n2578 ;
  assign n2656 = n2654 | n2655 ;
  assign n2657 = n1967 & n2643 ;
  assign n2658 = n2656 & n2657 ;
  assign n2659 = n2653 | n2658 ;
  assign n2660 = n224 & ~n2659 ;
  assign n2661 = n224 & ~n2660 ;
  assign n2662 = ( n2659 & n2660 ) | ( n2659 & ~n2661 ) | ( n2660 & ~n2661 );
  assign n2663 = n2645 | n2662 ;
  assign n2664 = n224 & n2662 ;
  assign n2665 = ~n2644 & n2664 ;
  assign n2666 = n375 | n709 ;
  assign n2667 = n375 & n709 ;
  assign n2668 = n2666 & ~n2667 ;
  assign n2669 = ~n700 & n906 ;
  assign n2670 = n700 & ~n906 ;
  assign n2671 = n2669 | n2670 ;
  assign n2672 = n2668 & ~n2671 ;
  assign n2673 = ~n700 & n709 ;
  assign n2674 = n700 & ~n709 ;
  assign n2675 = n2673 | n2674 ;
  assign n2676 = n2672 & ~n2675 ;
  assign n2677 = ~n2572 & n2676 ;
  assign n2678 = ~n2671 & n2675 ;
  assign n2679 = n2569 & n2678 ;
  assign n2680 = ~n2668 & n2671 ;
  assign n2681 = n2566 & n2680 ;
  assign n2682 = n2679 | n2681 ;
  assign n2683 = n2677 | n2682 ;
  assign n2684 = n2668 & n2671 ;
  assign n2685 = n2583 & ~n2586 ;
  assign n2686 = n2584 & ~n2587 ;
  assign n2687 = n2685 | n2686 ;
  assign n2688 = n2684 & n2687 ;
  assign n2689 = n2683 | n2688 ;
  assign n2690 = n375 | n2689 ;
  assign n2691 = n375 & n2689 ;
  assign n2692 = n2690 & ~n2691 ;
  assign n2693 = ~n2665 & n2692 ;
  assign n2694 = n2663 & n2693 ;
  assign n2695 = n2578 & n2671 ;
  assign n2696 = n375 & ~n2695 ;
  assign n2697 = n2578 & n2678 ;
  assign n2698 = n2576 & n2680 ;
  assign n2699 = n2697 | n2698 ;
  assign n2700 = n2656 & n2684 ;
  assign n2701 = n2699 | n2700 ;
  assign n2702 = n375 & ~n2701 ;
  assign n2703 = ~n375 & n2701 ;
  assign n2704 = n2702 | n2703 ;
  assign n2705 = n2696 & n2704 ;
  assign n2706 = n2572 & ~n2655 ;
  assign n2707 = ~n2572 & n2655 ;
  assign n2708 = n2706 | n2707 ;
  assign n2709 = n2684 & ~n2708 ;
  assign n2710 = ~n2572 & n2680 ;
  assign n2711 = n2578 & n2676 ;
  assign n2712 = n2576 & n2678 ;
  assign n2713 = n2711 | n2712 ;
  assign n2714 = n2710 | n2713 ;
  assign n2715 = n2709 | n2714 ;
  assign n2716 = n375 | n2715 ;
  assign n2717 = n375 & n2715 ;
  assign n2718 = n2716 & ~n2717 ;
  assign n2719 = n2705 & n2718 ;
  assign n2720 = n2644 & n2719 ;
  assign n2721 = n2644 | n2719 ;
  assign n2722 = ~n2720 & n2721 ;
  assign n2723 = ~n2572 & n2678 ;
  assign n2724 = n2569 & n2680 ;
  assign n2725 = n2576 & n2676 ;
  assign n2726 = n2724 | n2725 ;
  assign n2727 = n2723 | n2726 ;
  assign n2728 = n2580 & ~n2582 ;
  assign n2729 = n2574 | n2583 ;
  assign n2730 = ~n2728 & n2729 ;
  assign n2731 = n2684 & ~n2730 ;
  assign n2732 = n2727 | n2731 ;
  assign n2733 = n375 & n2732 ;
  assign n2734 = n375 | n2732 ;
  assign n2735 = ~n2733 & n2734 ;
  assign n2736 = n2722 & n2735 ;
  assign n2737 = n2720 | n2736 ;
  assign n2738 = n2663 & ~n2665 ;
  assign n2739 = n2692 | n2738 ;
  assign n2740 = ~n2694 & n2739 ;
  assign n2741 = n2737 & n2740 ;
  assign n2742 = n2694 | n2741 ;
  assign n2743 = ~n2572 & n2651 ;
  assign n2744 = n1967 & ~n2643 ;
  assign n2745 = ~n2648 & n2744 ;
  assign n2746 = n2578 & n2745 ;
  assign n2747 = n2576 & n2649 ;
  assign n2748 = n2746 | n2747 ;
  assign n2749 = n2743 | n2748 ;
  assign n2750 = n2657 & ~n2708 ;
  assign n2751 = n2749 | n2750 ;
  assign n2752 = n224 | n2751 ;
  assign n2753 = n224 & n2751 ;
  assign n2754 = n2752 & ~n2753 ;
  assign n2755 = n2665 & n2754 ;
  assign n2756 = n2665 | n2754 ;
  assign n2757 = ~n2755 & n2756 ;
  assign n2758 = n2587 | n2589 ;
  assign n2759 = ~n2590 & n2758 ;
  assign n2760 = n2684 & n2759 ;
  assign n2761 = n2561 & n2680 ;
  assign n2762 = n2569 & n2676 ;
  assign n2763 = n2566 & n2678 ;
  assign n2764 = n2762 | n2763 ;
  assign n2765 = n2761 | n2764 ;
  assign n2766 = n2760 | n2765 ;
  assign n2767 = n375 | n2766 ;
  assign n2768 = n375 & n2766 ;
  assign n2769 = n2767 & ~n2768 ;
  assign n2770 = n2757 & n2769 ;
  assign n2771 = n2757 | n2769 ;
  assign n2772 = ~n2770 & n2771 ;
  assign n2773 = n2742 | n2772 ;
  assign n2774 = n2742 & n2772 ;
  assign n2775 = n2773 & ~n2774 ;
  assign n2776 = ~n2597 & n2599 ;
  assign n2777 = n2600 | n2776 ;
  assign n2778 = ~n782 & n906 ;
  assign n2779 = n782 & ~n906 ;
  assign n2780 = n2778 | n2779 ;
  assign n2781 = n1081 & ~n1190 ;
  assign n2782 = ~n1081 & n1190 ;
  assign n2783 = n2781 | n2782 ;
  assign n2784 = n2780 & n2783 ;
  assign n2785 = ~n2777 & n2784 ;
  assign n2786 = ~n2780 & n2783 ;
  assign n2787 = n2552 & n2786 ;
  assign n2788 = ~n782 & n1081 ;
  assign n2789 = n782 & ~n1081 ;
  assign n2790 = n2788 | n2789 ;
  assign n2791 = ~n2783 & n2790 ;
  assign n2792 = ~n2555 & n2791 ;
  assign n2793 = n2780 & ~n2783 ;
  assign n2794 = ~n2790 & n2793 ;
  assign n2795 = n2558 & n2794 ;
  assign n2796 = n2792 | n2795 ;
  assign n2797 = n2787 | n2796 ;
  assign n2798 = n2785 | n2797 ;
  assign n2799 = n906 | n2798 ;
  assign n2800 = n906 & n2798 ;
  assign n2801 = n2799 & ~n2800 ;
  assign n2802 = n2775 & n2801 ;
  assign n2803 = n2737 | n2740 ;
  assign n2804 = ~n2741 & n2803 ;
  assign n2805 = ~n2593 & n2595 ;
  assign n2806 = n2596 | n2805 ;
  assign n2807 = n2784 & ~n2806 ;
  assign n2808 = ~n2555 & n2786 ;
  assign n2809 = n2561 & n2794 ;
  assign n2810 = n2558 & n2791 ;
  assign n2811 = n2809 | n2810 ;
  assign n2812 = n2808 | n2811 ;
  assign n2813 = n2807 | n2812 ;
  assign n2814 = n906 & ~n2813 ;
  assign n2815 = ~n906 & n2813 ;
  assign n2816 = n2814 | n2815 ;
  assign n2817 = n2804 & n2816 ;
  assign n2818 = n2722 | n2735 ;
  assign n2819 = ~n2736 & n2818 ;
  assign n2820 = n2564 | n2591 ;
  assign n2821 = ~n2592 & n2820 ;
  assign n2822 = n2784 & n2821 ;
  assign n2823 = n2558 & n2786 ;
  assign n2824 = n2566 & n2794 ;
  assign n2825 = n2561 & n2791 ;
  assign n2826 = n2824 | n2825 ;
  assign n2827 = n2823 | n2826 ;
  assign n2828 = n2822 | n2827 ;
  assign n2829 = n906 | n2828 ;
  assign n2830 = n906 & n2828 ;
  assign n2831 = n2829 & ~n2830 ;
  assign n2832 = n2819 & n2831 ;
  assign n2833 = n2705 | n2718 ;
  assign n2834 = ~n2719 & n2833 ;
  assign n2835 = n2561 & n2786 ;
  assign n2836 = n2569 & n2794 ;
  assign n2837 = n2566 & n2791 ;
  assign n2838 = n2836 | n2837 ;
  assign n2839 = n2835 | n2838 ;
  assign n2840 = n2759 & n2784 ;
  assign n2841 = n2839 | n2840 ;
  assign n2842 = n906 & ~n2841 ;
  assign n2843 = ~n906 & n2841 ;
  assign n2844 = n2842 | n2843 ;
  assign n2845 = n2834 & n2844 ;
  assign n2846 = n2696 | n2704 ;
  assign n2847 = ~n2705 & n2846 ;
  assign n2848 = n2687 & n2784 ;
  assign n2849 = ~n2572 & n2794 ;
  assign n2850 = n2569 & n2791 ;
  assign n2851 = n2566 & n2786 ;
  assign n2852 = n2850 | n2851 ;
  assign n2853 = n2849 | n2852 ;
  assign n2854 = n2848 | n2853 ;
  assign n2855 = n906 | n2854 ;
  assign n2856 = n906 & n2854 ;
  assign n2857 = n2855 & ~n2856 ;
  assign n2858 = n2847 & n2857 ;
  assign n2859 = n2847 | n2857 ;
  assign n2860 = ~n2858 & n2859 ;
  assign n2861 = ~n2572 & n2786 ;
  assign n2862 = ~n2708 & n2784 ;
  assign n2863 = n2576 & n2791 ;
  assign n2864 = n2578 & n2794 ;
  assign n2865 = n2863 | n2864 ;
  assign n2866 = n2862 | n2865 ;
  assign n2867 = n2861 | n2866 ;
  assign n2868 = n906 | n2867 ;
  assign n2869 = n906 & n2867 ;
  assign n2870 = n2868 & ~n2869 ;
  assign n2871 = n2578 & n2783 ;
  assign n2872 = n906 & ~n2871 ;
  assign n2873 = n2578 & n2791 ;
  assign n2874 = n2656 & n2784 ;
  assign n2875 = n2576 & n2786 ;
  assign n2876 = n2874 | n2875 ;
  assign n2877 = n2873 | n2876 ;
  assign n2878 = n906 & ~n2877 ;
  assign n2879 = ~n906 & n2877 ;
  assign n2880 = n2878 | n2879 ;
  assign n2881 = n2872 & n2880 ;
  assign n2882 = n2870 & n2881 ;
  assign n2883 = n2695 & n2882 ;
  assign n2884 = n2695 | n2882 ;
  assign n2885 = ~n2883 & n2884 ;
  assign n2886 = ~n2730 & n2784 ;
  assign n2887 = ~n2572 & n2791 ;
  assign n2888 = n2569 & n2786 ;
  assign n2889 = n2576 & n2794 ;
  assign n2890 = n2888 | n2889 ;
  assign n2891 = n2887 | n2890 ;
  assign n2892 = n2886 | n2891 ;
  assign n2893 = n906 & ~n2892 ;
  assign n2894 = n906 & ~n2893 ;
  assign n2895 = ( n2892 & n2893 ) | ( n2892 & ~n2894 ) | ( n2893 & ~n2894 );
  assign n2896 = n2885 & n2895 ;
  assign n2897 = n2883 | n2896 ;
  assign n2898 = n2860 & n2897 ;
  assign n2899 = n2858 | n2898 ;
  assign n2900 = n2834 | n2844 ;
  assign n2901 = ~n2845 & n2900 ;
  assign n2902 = n2899 & n2901 ;
  assign n2903 = n2845 | n2902 ;
  assign n2904 = n2819 | n2831 ;
  assign n2905 = ~n2832 & n2904 ;
  assign n2906 = n2903 & n2905 ;
  assign n2907 = n2832 | n2906 ;
  assign n2908 = n2804 | n2816 ;
  assign n2909 = ~n2817 & n2908 ;
  assign n2910 = n2907 & n2909 ;
  assign n2911 = n2817 | n2910 ;
  assign n2912 = n2775 | n2801 ;
  assign n2913 = ~n2802 & n2912 ;
  assign n2914 = n2911 & n2913 ;
  assign n2915 = n2802 | n2914 ;
  assign n2916 = n2770 | n2774 ;
  assign n2917 = ~n2572 & n2649 ;
  assign n2918 = n2569 & n2651 ;
  assign n2919 = n2576 & n2745 ;
  assign n2920 = n2918 | n2919 ;
  assign n2921 = n2917 | n2920 ;
  assign n2922 = n2657 & ~n2730 ;
  assign n2923 = n2921 | n2922 ;
  assign n2924 = n224 & ~n2923 ;
  assign n2925 = ~n224 & n2923 ;
  assign n2926 = n2924 | n2925 ;
  assign n2927 = n224 & n2578 ;
  assign n2928 = n2755 | n2927 ;
  assign n2929 = n2662 & n2927 ;
  assign n2930 = n2754 & n2929 ;
  assign n2931 = ~n2644 & n2930 ;
  assign n2932 = n2928 & ~n2931 ;
  assign n2933 = n2926 & n2932 ;
  assign n2934 = n2926 | n2932 ;
  assign n2935 = ~n2933 & n2934 ;
  assign n2936 = n2558 & n2680 ;
  assign n2937 = n2566 & n2676 ;
  assign n2938 = n2561 & n2678 ;
  assign n2939 = n2937 | n2938 ;
  assign n2940 = n2936 | n2939 ;
  assign n2941 = n2684 & n2821 ;
  assign n2942 = n2940 | n2941 ;
  assign n2943 = n375 & n2942 ;
  assign n2944 = n375 | n2942 ;
  assign n2945 = ~n2943 & n2944 ;
  assign n2946 = n2935 & n2945 ;
  assign n2947 = n2935 | n2945 ;
  assign n2948 = ~n2946 & n2947 ;
  assign n2949 = n2916 & n2948 ;
  assign n2950 = n2916 | n2948 ;
  assign n2951 = ~n2949 & n2950 ;
  assign n2952 = n2601 | n2603 ;
  assign n2953 = ~n2604 & n2952 ;
  assign n2954 = n2784 & n2953 ;
  assign n2955 = n2549 & n2786 ;
  assign n2956 = n2552 & n2791 ;
  assign n2957 = ~n2555 & n2794 ;
  assign n2958 = n2956 | n2957 ;
  assign n2959 = n2955 | n2958 ;
  assign n2960 = n2954 | n2959 ;
  assign n2961 = n906 | n2960 ;
  assign n2962 = n906 & n2960 ;
  assign n2963 = n2961 & ~n2962 ;
  assign n2964 = n2951 & n2963 ;
  assign n2965 = n2951 | n2963 ;
  assign n2966 = ~n2964 & n2965 ;
  assign n2967 = n2915 & n2966 ;
  assign n2968 = n2802 | n2966 ;
  assign n2969 = n2914 | n2968 ;
  assign n2970 = ~n1190 & n1233 ;
  assign n2971 = n1190 & ~n1233 ;
  assign n2972 = n2970 | n2971 ;
  assign n2973 = n32 & ~n1314 ;
  assign n2974 = ~n32 & n1314 ;
  assign n2975 = n2973 | n2974 ;
  assign n2976 = ~n2972 & n2975 ;
  assign n2977 = n2538 & n2976 ;
  assign n2978 = n1233 & ~n1314 ;
  assign n2979 = ~n1233 & n1314 ;
  assign n2980 = n2978 | n2979 ;
  assign n2981 = n2972 & ~n2975 ;
  assign n2982 = ~n2980 & n2981 ;
  assign n2983 = n2544 & n2982 ;
  assign n2984 = ~n2975 & n2980 ;
  assign n2985 = ~n2541 & n2984 ;
  assign n2986 = n2983 | n2985 ;
  assign n2987 = n2977 | n2986 ;
  assign n2988 = n2972 & n2975 ;
  assign n2989 = n2611 & ~n2613 ;
  assign n2990 = ~n2611 & n2613 ;
  assign n2991 = n2989 | n2990 ;
  assign n2992 = n2988 & ~n2991 ;
  assign n2993 = n2987 | n2992 ;
  assign n2994 = n1190 & n2993 ;
  assign n2995 = n1190 | n2993 ;
  assign n2996 = ~n2994 & n2995 ;
  assign n2997 = n2969 & n2996 ;
  assign n2998 = ~n2967 & n2997 ;
  assign n2999 = n2817 | n2913 ;
  assign n3000 = n2910 | n2999 ;
  assign n3001 = ~n2541 & n2976 ;
  assign n3002 = n2549 & n2982 ;
  assign n3003 = n2544 & n2984 ;
  assign n3004 = n3002 | n3003 ;
  assign n3005 = n3001 | n3004 ;
  assign n3006 = ~n2547 & n2609 ;
  assign n3007 = n2547 & ~n2609 ;
  assign n3008 = n3006 | n3007 ;
  assign n3009 = n2988 & ~n3008 ;
  assign n3010 = n3005 | n3009 ;
  assign n3011 = n1190 & n3010 ;
  assign n3012 = n1190 | n3010 ;
  assign n3013 = ~n3011 & n3012 ;
  assign n3014 = n3000 & n3013 ;
  assign n3015 = ~n2914 & n3014 ;
  assign n3016 = n2832 | n2909 ;
  assign n3017 = n2906 | n3016 ;
  assign n3018 = n2544 & n2976 ;
  assign n3019 = n2605 | n2607 ;
  assign n3020 = ~n2608 & n3019 ;
  assign n3021 = n2988 & n3020 ;
  assign n3022 = n2552 & n2982 ;
  assign n3023 = n2549 & n2984 ;
  assign n3024 = n3022 | n3023 ;
  assign n3025 = n3021 | n3024 ;
  assign n3026 = n3018 | n3025 ;
  assign n3027 = n1190 | n3026 ;
  assign n3028 = n1190 & n3026 ;
  assign n3029 = n3027 & ~n3028 ;
  assign n3030 = n3017 & n3029 ;
  assign n3031 = ~n2910 & n3030 ;
  assign n3032 = n2845 | n2905 ;
  assign n3033 = n2902 | n3032 ;
  assign n3034 = n2549 & n2976 ;
  assign n3035 = n2953 & n2988 ;
  assign n3036 = ~n2555 & n2982 ;
  assign n3037 = n2552 & n2984 ;
  assign n3038 = n3036 | n3037 ;
  assign n3039 = n3035 | n3038 ;
  assign n3040 = n3034 | n3039 ;
  assign n3041 = n1190 | n3040 ;
  assign n3042 = n1190 & n3040 ;
  assign n3043 = n3041 & ~n3042 ;
  assign n3044 = n3033 & n3043 ;
  assign n3045 = ~n2906 & n3044 ;
  assign n3046 = ~n2906 & n3033 ;
  assign n3047 = n3043 | n3046 ;
  assign n3048 = n2899 | n2901 ;
  assign n3049 = ~n2902 & n3048 ;
  assign n3050 = n2552 & n2976 ;
  assign n3051 = ~n2777 & n2988 ;
  assign n3052 = n2558 & n2982 ;
  assign n3053 = ~n2555 & n2984 ;
  assign n3054 = n3052 | n3053 ;
  assign n3055 = n3051 | n3054 ;
  assign n3056 = n3050 | n3055 ;
  assign n3057 = n1190 | n3056 ;
  assign n3058 = n1190 & n3056 ;
  assign n3059 = n3057 & ~n3058 ;
  assign n3060 = n3049 & n3059 ;
  assign n3061 = n2860 | n2897 ;
  assign n3062 = ~n2898 & n3061 ;
  assign n3063 = ~n2555 & n2976 ;
  assign n3064 = ~n2806 & n2988 ;
  assign n3065 = n2561 & n2982 ;
  assign n3066 = n2558 & n2984 ;
  assign n3067 = n3065 | n3066 ;
  assign n3068 = n3064 | n3067 ;
  assign n3069 = n3063 | n3068 ;
  assign n3070 = n1190 & n3069 ;
  assign n3071 = n1190 | n3069 ;
  assign n3072 = ~n3070 & n3071 ;
  assign n3073 = n3062 & n3072 ;
  assign n3074 = n2885 | n2895 ;
  assign n3075 = ~n2896 & n3074 ;
  assign n3076 = n2821 & n2988 ;
  assign n3077 = n2558 & n2976 ;
  assign n3078 = n2566 & n2982 ;
  assign n3079 = n2561 & n2984 ;
  assign n3080 = n3078 | n3079 ;
  assign n3081 = n3077 | n3080 ;
  assign n3082 = n3076 | n3081 ;
  assign n3083 = n1190 & n3082 ;
  assign n3084 = n1190 | n3082 ;
  assign n3085 = ~n3083 & n3084 ;
  assign n3086 = n3075 & n3085 ;
  assign n3087 = n2870 | n2881 ;
  assign n3088 = ~n2882 & n3087 ;
  assign n3089 = n2561 & n2976 ;
  assign n3090 = n2569 & n2982 ;
  assign n3091 = n2566 & n2984 ;
  assign n3092 = n3090 | n3091 ;
  assign n3093 = n3089 | n3092 ;
  assign n3094 = n2759 & n2988 ;
  assign n3095 = n3093 | n3094 ;
  assign n3096 = n1190 & n3095 ;
  assign n3097 = n1190 | n3095 ;
  assign n3098 = ~n3096 & n3097 ;
  assign n3099 = n3088 & n3098 ;
  assign n3100 = ~n2572 & n2982 ;
  assign n3101 = n2569 & n2984 ;
  assign n3102 = n2566 & n2976 ;
  assign n3103 = n3101 | n3102 ;
  assign n3104 = n3100 | n3103 ;
  assign n3105 = n2687 & n2988 ;
  assign n3106 = n3104 | n3105 ;
  assign n3107 = n1190 | n3106 ;
  assign n3108 = n1190 & n3106 ;
  assign n3109 = n3107 & ~n3108 ;
  assign n3110 = n2872 | n2880 ;
  assign n3111 = ~n2881 & n3110 ;
  assign n3112 = n3109 & n3111 ;
  assign n3113 = n2578 & n2984 ;
  assign n3114 = n2656 & n2988 ;
  assign n3115 = n2576 & n2976 ;
  assign n3116 = n3114 | n3115 ;
  assign n3117 = n3113 | n3116 ;
  assign n3118 = n1190 & n3117 ;
  assign n3119 = ~n2708 & n2988 ;
  assign n3120 = n2576 & n2984 ;
  assign n3121 = n3119 | n3120 ;
  assign n3122 = n2578 & n2982 ;
  assign n3123 = ~n2572 & n2976 ;
  assign n3124 = n1190 | n3123 ;
  assign n3125 = n3122 | n3124 ;
  assign n3126 = n3121 | n3125 ;
  assign n3127 = ~n3118 & n3126 ;
  assign n3128 = n3120 | n3123 ;
  assign n3129 = n3119 | n3128 ;
  assign n3130 = n3122 | n3129 ;
  assign n3131 = n1190 & n3130 ;
  assign n3132 = n1190 | n3113 ;
  assign n3133 = n3116 | n3132 ;
  assign n3134 = n2578 & n2975 ;
  assign n3135 = n1190 & n2871 ;
  assign n3136 = ~n3134 & n3135 ;
  assign n3137 = n3133 & n3136 ;
  assign n3138 = ~n3131 & n3137 ;
  assign n3139 = n3127 & n3138 ;
  assign n3140 = n3126 & ~n3131 ;
  assign n3141 = n1190 & ~n3134 ;
  assign n3142 = n3133 & n3141 ;
  assign n3143 = ~n3118 & n3142 ;
  assign n3144 = n3140 & n3143 ;
  assign n3145 = n2871 | n3144 ;
  assign n3146 = ~n2730 & n2988 ;
  assign n3147 = ~n2572 & n2984 ;
  assign n3148 = n2569 & n2976 ;
  assign n3149 = n2576 & n2982 ;
  assign n3150 = n3148 | n3149 ;
  assign n3151 = n3147 | n3150 ;
  assign n3152 = n3146 | n3151 ;
  assign n3153 = n1190 & n3152 ;
  assign n3154 = n1190 | n3152 ;
  assign n3155 = ~n3153 & n3154 ;
  assign n3156 = ~n3139 & n3155 ;
  assign n3157 = n3145 & n3156 ;
  assign n3158 = n3139 | n3157 ;
  assign n3159 = n3109 | n3111 ;
  assign n3160 = ~n3112 & n3159 ;
  assign n3161 = n3158 & n3160 ;
  assign n3162 = n3112 | n3161 ;
  assign n3163 = n3088 | n3098 ;
  assign n3164 = ~n3099 & n3163 ;
  assign n3165 = n3162 & n3164 ;
  assign n3166 = n3099 | n3165 ;
  assign n3167 = n3075 | n3085 ;
  assign n3168 = ~n3086 & n3167 ;
  assign n3169 = n3166 & n3168 ;
  assign n3170 = n3086 | n3169 ;
  assign n3171 = n3062 | n3072 ;
  assign n3172 = ~n3073 & n3171 ;
  assign n3173 = n3170 & n3172 ;
  assign n3174 = n3073 | n3173 ;
  assign n3175 = n3049 | n3059 ;
  assign n3176 = ~n3060 & n3175 ;
  assign n3177 = n3174 & n3176 ;
  assign n3178 = n3060 | n3177 ;
  assign n3179 = ~n3045 & n3178 ;
  assign n3180 = n3047 & n3179 ;
  assign n3181 = n3045 | n3180 ;
  assign n3182 = ~n2910 & n3017 ;
  assign n3183 = n3029 | n3182 ;
  assign n3184 = ~n3031 & n3183 ;
  assign n3185 = n3181 & n3184 ;
  assign n3186 = n3031 | n3185 ;
  assign n3187 = ~n2914 & n3000 ;
  assign n3188 = n3013 | n3187 ;
  assign n3189 = ~n3015 & n3188 ;
  assign n3190 = n3186 & n3189 ;
  assign n3191 = n3015 | n3190 ;
  assign n3192 = ~n2967 & n2969 ;
  assign n3193 = n2996 | n3192 ;
  assign n3194 = ~n2998 & n3193 ;
  assign n3195 = n3191 & n3194 ;
  assign n3196 = n2998 | n3195 ;
  assign n3197 = n2964 | n2967 ;
  assign n3198 = n2946 | n2949 ;
  assign n3199 = n2931 | n2933 ;
  assign n3200 = n224 & ~n2576 ;
  assign n3201 = ~n2572 & n2745 ;
  assign n3202 = n2569 & n2649 ;
  assign n3203 = n2566 & n2651 ;
  assign n3204 = n3202 | n3203 ;
  assign n3205 = n3201 | n3204 ;
  assign n3206 = n2657 & n2687 ;
  assign n3207 = n3205 | n3206 ;
  assign n3208 = n3200 | n3207 ;
  assign n3209 = n3200 & n3207 ;
  assign n3210 = n3208 & ~n3209 ;
  assign n3211 = n3199 & n3210 ;
  assign n3212 = n3199 | n3210 ;
  assign n3213 = ~n3211 & n3212 ;
  assign n3214 = ~n2555 & n2680 ;
  assign n3215 = n2561 & n2676 ;
  assign n3216 = n2558 & n2678 ;
  assign n3217 = n3215 | n3216 ;
  assign n3218 = n3214 | n3217 ;
  assign n3219 = n2684 & ~n2806 ;
  assign n3220 = n3218 | n3219 ;
  assign n3221 = n375 & n3220 ;
  assign n3222 = n375 | n3220 ;
  assign n3223 = ~n3221 & n3222 ;
  assign n3224 = n3213 & n3223 ;
  assign n3225 = n3213 | n3223 ;
  assign n3226 = ~n3224 & n3225 ;
  assign n3227 = n3198 & n3226 ;
  assign n3228 = n3198 | n3226 ;
  assign n3229 = ~n3227 & n3228 ;
  assign n3230 = n2784 & n3020 ;
  assign n3231 = n2544 & n2786 ;
  assign n3232 = n2549 & n2791 ;
  assign n3233 = n2552 & n2794 ;
  assign n3234 = n3232 | n3233 ;
  assign n3235 = n3231 | n3234 ;
  assign n3236 = n3230 | n3235 ;
  assign n3237 = n906 | n3236 ;
  assign n3238 = n906 & n3236 ;
  assign n3239 = n3237 & ~n3238 ;
  assign n3240 = n3229 & n3239 ;
  assign n3241 = n3229 | n3239 ;
  assign n3242 = ~n3240 & n3241 ;
  assign n3243 = n3197 & n3242 ;
  assign n3244 = n2964 | n3242 ;
  assign n3245 = n2967 | n3244 ;
  assign n3246 = ~n3243 & n3245 ;
  assign n3247 = n2618 & n2976 ;
  assign n3248 = ~n2541 & n2982 ;
  assign n3249 = n2538 & n2984 ;
  assign n3250 = n3248 | n3249 ;
  assign n3251 = n3247 | n3250 ;
  assign n3252 = n2615 & n2624 ;
  assign n3253 = n2615 | n2624 ;
  assign n3254 = ~n3252 & n3253 ;
  assign n3255 = n2988 & n3254 ;
  assign n3256 = n3251 | n3255 ;
  assign n3257 = n1190 & n3256 ;
  assign n3258 = n1190 | n3256 ;
  assign n3259 = ~n3257 & n3258 ;
  assign n3260 = n3246 | n3259 ;
  assign n3261 = n3245 & n3259 ;
  assign n3262 = ~n3243 & n3261 ;
  assign n3263 = n3260 & ~n3262 ;
  assign n3264 = n3196 & n3263 ;
  assign n3265 = n3196 | n3263 ;
  assign n3266 = ~n3264 & n3265 ;
  assign n3267 = n2640 & n3266 ;
  assign n3268 = n2640 | n3266 ;
  assign n3269 = ~n3267 & n3268 ;
  assign n3270 = n2518 & n2526 ;
  assign n3271 = n2522 & n2618 ;
  assign n3272 = ~n2521 & n2527 ;
  assign n3273 = n3271 | n3272 ;
  assign n3274 = n3270 | n3273 ;
  assign n3275 = ~n2521 & n2526 ;
  assign n3276 = ( n2521 & ~n2526 ) | ( n2521 & n2619 ) | ( ~n2526 & n2619 );
  assign n3277 = ( n2628 & ~n3275 ) | ( n2628 & n3276 ) | ( ~n3275 & n3276 );
  assign n3278 = n2619 | n2628 ;
  assign n3279 = ( n2521 & ~n3277 ) | ( n2521 & n3278 ) | ( ~n3277 & n3278 );
  assign n3280 = ( n2526 & n3277 ) | ( n2526 & ~n3279 ) | ( n3277 & ~n3279 );
  assign n3281 = n2531 & ~n3280 ;
  assign n3282 = n3274 | n3281 ;
  assign n3283 = n32 | n3282 ;
  assign n3284 = n32 & n3282 ;
  assign n3285 = n3283 & ~n3284 ;
  assign n3286 = n3191 | n3194 ;
  assign n3287 = ~n3195 & n3286 ;
  assign n3288 = n3285 & n3287 ;
  assign n3289 = n2518 & ~n2521 ;
  assign n3290 = n2522 & n2538 ;
  assign n3291 = n2527 & n2618 ;
  assign n3292 = n3290 | n3291 ;
  assign n3293 = n3289 | n3292 ;
  assign n3294 = ( n2615 & n2622 ) | ( n2615 & n2625 ) | ( n2622 & n2625 );
  assign n3295 = n2621 & ~n3294 ;
  assign n3296 = n2628 | n3295 ;
  assign n3297 = n2531 & ~n3296 ;
  assign n3298 = n3293 | n3297 ;
  assign n3299 = n32 | n3298 ;
  assign n3300 = n32 & n3298 ;
  assign n3301 = n3299 & ~n3300 ;
  assign n3302 = n3186 | n3189 ;
  assign n3303 = ~n3190 & n3302 ;
  assign n3304 = n3301 & n3303 ;
  assign n3305 = n3301 | n3303 ;
  assign n3306 = ~n3304 & n3305 ;
  assign n3307 = n2518 & n2618 ;
  assign n3308 = n2522 & ~n2541 ;
  assign n3309 = n2527 & n2538 ;
  assign n3310 = n3308 | n3309 ;
  assign n3311 = n3307 | n3310 ;
  assign n3312 = n2531 & n3254 ;
  assign n3313 = n3311 | n3312 ;
  assign n3314 = n32 & ~n3313 ;
  assign n3315 = ~n32 & n3313 ;
  assign n3316 = n3314 | n3315 ;
  assign n3317 = n3174 | n3176 ;
  assign n3318 = ~n3177 & n3317 ;
  assign n3319 = n3086 | n3172 ;
  assign n3320 = n3169 | n3319 ;
  assign n3321 = ~n3173 & n3320 ;
  assign n3322 = n2527 & n2549 ;
  assign n3323 = n2531 & n3020 ;
  assign n3324 = n2518 & n2544 ;
  assign n3325 = n3323 | n3324 ;
  assign n3326 = n2522 & n2552 ;
  assign n3327 = n3325 | n3326 ;
  assign n3328 = n3322 | n3327 ;
  assign n3329 = n32 & ~n3328 ;
  assign n3330 = ~n32 & n3328 ;
  assign n3331 = n3329 | n3330 ;
  assign n3332 = n3321 | n3331 ;
  assign n3333 = n3166 | n3168 ;
  assign n3334 = ~n3169 & n3333 ;
  assign n3335 = n2522 & ~n2555 ;
  assign n3336 = n2527 & n2552 ;
  assign n3337 = n3335 | n3336 ;
  assign n3338 = n2531 & n2953 ;
  assign n3339 = n2518 & n2549 ;
  assign n3340 = n3338 | n3339 ;
  assign n3341 = n3337 | n3340 ;
  assign n3342 = n32 & ~n3341 ;
  assign n3343 = ~n32 & n3341 ;
  assign n3344 = n3342 | n3343 ;
  assign n3345 = n3334 & n3344 ;
  assign n3346 = n3320 & n3331 ;
  assign n3347 = ~n3173 & n3346 ;
  assign n3348 = n3345 | n3347 ;
  assign n3349 = n3162 | n3164 ;
  assign n3350 = ~n3165 & n3349 ;
  assign n3351 = n2522 & n2558 ;
  assign n3352 = n2527 & ~n2555 ;
  assign n3353 = n3351 | n3352 ;
  assign n3354 = n2531 & ~n2777 ;
  assign n3355 = n2518 & n2552 ;
  assign n3356 = n3354 | n3355 ;
  assign n3357 = n3353 | n3356 ;
  assign n3358 = n32 & ~n3357 ;
  assign n3359 = ~n32 & n3357 ;
  assign n3360 = n3358 | n3359 ;
  assign n3361 = n3350 & n3360 ;
  assign n3362 = n2527 & n2558 ;
  assign n3363 = n2531 & ~n2806 ;
  assign n3364 = n2518 & ~n2555 ;
  assign n3365 = n3363 | n3364 ;
  assign n3366 = n2522 & n2561 ;
  assign n3367 = n3365 | n3366 ;
  assign n3368 = n3362 | n3367 ;
  assign n3369 = n32 & ~n3368 ;
  assign n3370 = ~n32 & n3368 ;
  assign n3371 = n3369 | n3370 ;
  assign n3372 = ~n3139 & n3145 ;
  assign n3373 = n3155 | n3372 ;
  assign n3374 = ~n3157 & n3373 ;
  assign n3375 = n2518 & n2558 ;
  assign n3376 = n2522 & n2566 ;
  assign n3377 = n2527 & n2561 ;
  assign n3378 = n3376 | n3377 ;
  assign n3379 = n2531 & n2821 ;
  assign n3380 = n3378 | n3379 ;
  assign n3381 = n3375 | n3380 ;
  assign n3382 = n32 & ~n3381 ;
  assign n3383 = ~n32 & n3381 ;
  assign n3384 = n3382 | n3383 ;
  assign n3385 = n3374 | n3384 ;
  assign n3386 = n2518 & n2561 ;
  assign n3387 = n2522 & n2569 ;
  assign n3388 = n2527 & n2566 ;
  assign n3389 = n3387 | n3388 ;
  assign n3390 = n3386 | n3389 ;
  assign n3391 = n2531 & n2759 ;
  assign n3392 = n3390 | n3391 ;
  assign n3393 = n32 & ~n3392 ;
  assign n3394 = ~n32 & n3392 ;
  assign n3395 = n3393 | n3394 ;
  assign n3396 = n3140 | n3143 ;
  assign n3397 = ~n3144 & n3396 ;
  assign n3398 = n3395 & n3397 ;
  assign n3399 = ~n3118 & n3133 ;
  assign n3400 = n3141 | n3399 ;
  assign n3401 = ~n3143 & n3400 ;
  assign n3402 = n2518 & n2566 ;
  assign n3403 = n2531 & n2687 ;
  assign n3404 = n2522 & ~n2572 ;
  assign n3405 = n3403 | n3404 ;
  assign n3406 = n2527 & n2569 ;
  assign n3407 = n3405 | n3406 ;
  assign n3408 = n3402 | n3407 ;
  assign n3409 = n32 & ~n3408 ;
  assign n3410 = ~n32 & n3408 ;
  assign n3411 = n3409 | n3410 ;
  assign n3412 = n3401 | n3411 ;
  assign n3413 = n3395 | n3397 ;
  assign n3414 = n3412 & n3413 ;
  assign n3415 = n3401 & n3411 ;
  assign n3416 = n2518 & n2576 ;
  assign n3417 = ~n2656 & n2708 ;
  assign n3418 = n2531 & ~n3417 ;
  assign n3419 = n3416 | n3418 ;
  assign n3420 = pi0 | n2514 ;
  assign n3421 = n2578 & n3420 ;
  assign n3422 = n32 & ~n3421 ;
  assign n3423 = n2518 & ~n2572 ;
  assign n3424 = n2522 & n2578 ;
  assign n3425 = n2527 & n2576 ;
  assign n3426 = n3424 | n3425 ;
  assign n3427 = n3423 | n3426 ;
  assign n3428 = n3422 & ~n3427 ;
  assign n3429 = ~n3419 & n3428 ;
  assign n3430 = n3134 & n3429 ;
  assign n3431 = n3134 | n3429 ;
  assign n3432 = n2531 & ~n2730 ;
  assign n3433 = n2527 & ~n2572 ;
  assign n3434 = n2518 & n2569 ;
  assign n3435 = n2522 & n2576 ;
  assign n3436 = n3434 | n3435 ;
  assign n3437 = n3433 | n3436 ;
  assign n3438 = n3432 | n3437 ;
  assign n3439 = n32 & ~n3438 ;
  assign n3440 = ~n32 & n3438 ;
  assign n3441 = n3439 | n3440 ;
  assign n3442 = n3431 & n3441 ;
  assign n3443 = n3430 | n3442 ;
  assign n3444 = n3415 | n3443 ;
  assign n3445 = n3414 & n3444 ;
  assign n3446 = ~n3157 & n3384 ;
  assign n3447 = n3373 & n3446 ;
  assign n3448 = n3445 | n3447 ;
  assign n3449 = n3398 | n3448 ;
  assign n3450 = n3385 & n3449 ;
  assign n3451 = n3371 & n3450 ;
  assign n3452 = n3361 | n3451 ;
  assign n3453 = n3371 | n3450 ;
  assign n3454 = n3158 | n3160 ;
  assign n3455 = ~n3161 & n3454 ;
  assign n3456 = n3453 & n3455 ;
  assign n3457 = n3452 | n3456 ;
  assign n3458 = n3334 | n3344 ;
  assign n3459 = n3350 | n3360 ;
  assign n3460 = n3458 & n3459 ;
  assign n3461 = n3457 & n3460 ;
  assign n3462 = n3348 | n3461 ;
  assign n3463 = n3332 & n3462 ;
  assign n3464 = n3318 | n3463 ;
  assign n3465 = n3318 & n3463 ;
  assign n3466 = n2527 & n2544 ;
  assign n3467 = n2531 & ~n3008 ;
  assign n3468 = n3466 | n3467 ;
  assign n3469 = n2522 & n2549 ;
  assign n3470 = n2518 & ~n2541 ;
  assign n3471 = n3469 | n3470 ;
  assign n3472 = n3468 | n3471 ;
  assign n3473 = n32 & ~n3472 ;
  assign n3474 = ~n32 & n3472 ;
  assign n3475 = n3473 | n3474 ;
  assign n3476 = n3465 | n3475 ;
  assign n3477 = n3464 & n3476 ;
  assign n3478 = n2531 & ~n2991 ;
  assign n3479 = n2518 & n2538 ;
  assign n3480 = n2522 & n2544 ;
  assign n3481 = n2527 & ~n2541 ;
  assign n3482 = n3480 | n3481 ;
  assign n3483 = n3479 | n3482 ;
  assign n3484 = n3478 | n3483 ;
  assign n3485 = n32 & ~n3484 ;
  assign n3486 = ~n32 & n3484 ;
  assign n3487 = n3485 | n3486 ;
  assign n3488 = n3477 & n3487 ;
  assign n3489 = n3477 | n3487 ;
  assign n3490 = ~n3045 & n3047 ;
  assign n3491 = n3178 | n3490 ;
  assign n3492 = ~n3180 & n3491 ;
  assign n3493 = n3489 & n3492 ;
  assign n3494 = n3488 | n3493 ;
  assign n3495 = n3316 & n3494 ;
  assign n3496 = n3181 | n3184 ;
  assign n3497 = n3316 | n3494 ;
  assign n3498 = ~n3185 & n3497 ;
  assign n3499 = n3496 & n3498 ;
  assign n3500 = n3495 | n3499 ;
  assign n3501 = n3306 & n3500 ;
  assign n3502 = n3304 | n3501 ;
  assign n3503 = n3285 | n3287 ;
  assign n3504 = ~n3288 & n3503 ;
  assign n3505 = n3502 & n3504 ;
  assign n3506 = n3288 | n3505 ;
  assign n3507 = n3269 & n3506 ;
  assign n3508 = n3269 | n3506 ;
  assign n3509 = ~n3507 & n3508 ;
  assign n3510 = n320 | n342 ;
  assign n3511 = n200 | n2445 ;
  assign n3512 = n477 | n3511 ;
  assign n3513 = n177 | n191 ;
  assign n3514 = n247 | n3513 ;
  assign n3515 = n433 | n3514 ;
  assign n3516 = n271 | n3515 ;
  assign n3517 = n153 | n512 ;
  assign n3518 = n190 | n3517 ;
  assign n3519 = n3516 | n3518 ;
  assign n3520 = n274 | n3519 ;
  assign n3521 = n444 | n3520 ;
  assign n3522 = n3512 | n3521 ;
  assign n3523 = n140 | n248 ;
  assign n3524 = n124 | n3523 ;
  assign n3525 = n157 | n336 ;
  assign n3526 = n503 | n513 ;
  assign n3527 = n170 | n2086 ;
  assign n3528 = n179 | n281 ;
  assign n3529 = n142 | n186 ;
  assign n3530 = n194 | n3529 ;
  assign n3531 = n3528 | n3530 ;
  assign n3532 = n227 | n3531 ;
  assign n3533 = n204 | n3532 ;
  assign n3534 = n3527 | n3533 ;
  assign n3535 = n3526 | n3534 ;
  assign n3536 = n3525 | n3535 ;
  assign n3537 = n3524 | n3536 ;
  assign n3538 = n392 | n3537 ;
  assign n3539 = n284 | n304 ;
  assign n3540 = n167 | n3539 ;
  assign n3541 = n3538 | n3540 ;
  assign n3542 = n382 | n3541 ;
  assign n3543 = n106 | n3542 ;
  assign n3544 = n1980 | n3543 ;
  assign n3545 = n3522 | n3544 ;
  assign n3546 = n3510 | n3545 ;
  assign n3547 = n145 | n164 ;
  assign n3548 = n255 | n3547 ;
  assign n3549 = n3546 | n3548 ;
  assign n3550 = n269 | n3549 ;
  assign n3551 = n3509 & n3550 ;
  assign n3552 = n3509 | n3550 ;
  assign n3553 = ~n3551 & n3552 ;
  assign n3554 = n251 | n282 ;
  assign n3555 = n238 | n3554 ;
  assign n3556 = n158 | n615 ;
  assign n3557 = n239 | n263 ;
  assign n3558 = n337 | n392 ;
  assign n3559 = n296 | n1032 ;
  assign n3560 = n3558 | n3559 ;
  assign n3561 = n3557 | n3560 ;
  assign n3562 = n248 | n317 ;
  assign n3563 = n232 | n234 ;
  assign n3564 = n3562 | n3563 ;
  assign n3565 = n135 | n145 ;
  assign n3566 = n399 | n499 ;
  assign n3567 = n3565 | n3566 ;
  assign n3568 = n3564 | n3567 ;
  assign n3569 = n3561 | n3568 ;
  assign n3570 = n328 | n3569 ;
  assign n3571 = n3556 | n3570 ;
  assign n3572 = n179 | n321 ;
  assign n3573 = n3571 | n3572 ;
  assign n3574 = n148 | n170 ;
  assign n3575 = n109 | n3574 ;
  assign n3576 = n3573 | n3575 ;
  assign n3577 = n209 | n305 ;
  assign n3578 = n208 | n618 ;
  assign n3579 = n331 | n342 ;
  assign n3580 = n403 | n589 ;
  assign n3581 = n3579 | n3580 ;
  assign n3582 = n146 | n151 ;
  assign n3583 = n3581 | n3582 ;
  assign n3584 = n3578 | n3583 ;
  assign n3585 = n255 | n3584 ;
  assign n3586 = n293 | n3585 ;
  assign n3587 = n3577 | n3586 ;
  assign n3588 = n180 | n201 ;
  assign n3589 = n273 | n2111 ;
  assign n3590 = n3588 | n3589 ;
  assign n3591 = n205 | n314 ;
  assign n3592 = n1046 | n3591 ;
  assign n3593 = n275 | n3592 ;
  assign n3594 = n3590 | n3593 ;
  assign n3595 = n3587 | n3594 ;
  assign n3596 = n3576 | n3595 ;
  assign n3597 = n3555 | n3596 ;
  assign n3598 = n3502 | n3504 ;
  assign n3599 = ~n3505 & n3598 ;
  assign n3600 = n3597 & n3599 ;
  assign n3601 = n3306 | n3500 ;
  assign n3602 = ~n3501 & n3601 ;
  assign n3603 = n137 | n146 ;
  assign n3604 = n405 | n3603 ;
  assign n3605 = n140 | n195 ;
  assign n3606 = n176 | n2007 ;
  assign n3607 = n109 | n3606 ;
  assign n3608 = n626 | n3607 ;
  assign n3609 = n298 | n3608 ;
  assign n3610 = n2231 | n3609 ;
  assign n3611 = n243 | n343 ;
  assign n3612 = n252 | n3611 ;
  assign n3613 = n202 | n2160 ;
  assign n3614 = n163 | n3613 ;
  assign n3615 = n2127 | n3614 ;
  assign n3616 = n3612 | n3615 ;
  assign n3617 = n2249 | n2304 ;
  assign n3618 = n422 | n3617 ;
  assign n3619 = n3616 | n3618 ;
  assign n3620 = n3610 | n3619 ;
  assign n3621 = n3605 | n3620 ;
  assign n3622 = n3604 | n3621 ;
  assign n3623 = n157 | n3622 ;
  assign n3624 = n334 | n3623 ;
  assign n3625 = n3597 | n3599 ;
  assign n3626 = n3624 & n3625 ;
  assign n3627 = n3602 & n3626 ;
  assign n3628 = n3600 | n3627 ;
  assign n3629 = n3553 & n3628 ;
  assign n3630 = n3553 | n3628 ;
  assign n3631 = ~n3629 & n3630 ;
  assign n3632 = n3551 | n3629 ;
  assign n3633 = n3267 | n3507 ;
  assign n3634 = n200 | n234 ;
  assign n3635 = n192 | n484 ;
  assign n3636 = n3634 | n3635 ;
  assign n3637 = n164 | n205 ;
  assign n3638 = n230 | n3526 ;
  assign n3639 = n3637 | n3638 ;
  assign n3640 = n3636 | n3639 ;
  assign n3641 = n672 | n3640 ;
  assign n3642 = n268 | n460 ;
  assign n3643 = n186 | n3642 ;
  assign n3644 = n2003 | n3643 ;
  assign n3645 = n1067 | n3644 ;
  assign n3646 = n3641 | n3645 ;
  assign n3647 = n170 | n1319 ;
  assign n3648 = n1064 & ~n2112 ;
  assign n3649 = ~n157 & n3648 ;
  assign n3650 = ~n3647 & n3649 ;
  assign n3651 = ~n3646 & n3650 ;
  assign n3652 = ~n227 & n3651 ;
  assign n3653 = ~n447 & n3652 ;
  assign n3654 = n2510 & n3653 ;
  assign n3655 = n2510 | n3653 ;
  assign n3656 = ~n3654 & n3655 ;
  assign n3657 = n2518 & ~n3656 ;
  assign n3658 = n2522 & n2526 ;
  assign n3659 = n2511 & n2527 ;
  assign n3660 = n3658 | n3659 ;
  assign n3661 = n3657 | n3660 ;
  assign n3662 = ~n2511 & n3656 ;
  assign n3663 = n2511 & ~n3656 ;
  assign n3664 = n3662 | n3663 ;
  assign n3665 = n2533 | n2632 ;
  assign n3666 = n3664 | n3665 ;
  assign n3667 = n2533 | n2633 ;
  assign n3668 = n3664 | n3667 ;
  assign n3669 = ( n2628 & n3666 ) | ( n2628 & n3668 ) | ( n3666 & n3668 );
  assign n3670 = ~n3664 & n3669 ;
  assign n3671 = ( n2628 & n3665 ) | ( n2628 & n3667 ) | ( n3665 & n3667 );
  assign n3672 = ( n3669 & n3670 ) | ( n3669 & ~n3671 ) | ( n3670 & ~n3671 );
  assign n3673 = n2531 & ~n3672 ;
  assign n3674 = n3661 | n3673 ;
  assign n3675 = n32 & ~n3674 ;
  assign n3676 = ~n32 & n3674 ;
  assign n3677 = n3675 | n3676 ;
  assign n3678 = n3262 | n3264 ;
  assign n3679 = n3240 | n3243 ;
  assign n3680 = n224 & n2572 ;
  assign n3681 = n2561 & n2651 ;
  assign n3682 = n2569 & n2745 ;
  assign n3683 = n2566 & n2649 ;
  assign n3684 = n3682 | n3683 ;
  assign n3685 = n3681 | n3684 ;
  assign n3686 = n2657 & n2759 ;
  assign n3687 = n3685 | n3686 ;
  assign n3688 = n3680 & n3687 ;
  assign n3689 = n3680 | n3687 ;
  assign n3690 = ~n3688 & n3689 ;
  assign n3691 = n224 & ~n3207 ;
  assign n3692 = n2576 & n3691 ;
  assign n3693 = n3211 | n3692 ;
  assign n3694 = n3690 & n3693 ;
  assign n3695 = n3690 | n3693 ;
  assign n3696 = ~n3694 & n3695 ;
  assign n3697 = n2552 & n2680 ;
  assign n3698 = n2558 & n2676 ;
  assign n3699 = ~n2555 & n2678 ;
  assign n3700 = n3698 | n3699 ;
  assign n3701 = n3697 | n3700 ;
  assign n3702 = n2684 & ~n2777 ;
  assign n3703 = n3701 | n3702 ;
  assign n3704 = n375 | n3703 ;
  assign n3705 = n375 & n3703 ;
  assign n3706 = n3704 & ~n3705 ;
  assign n3707 = n3696 & n3706 ;
  assign n3708 = n3696 | n3706 ;
  assign n3709 = ~n3707 & n3708 ;
  assign n3710 = n3224 | n3227 ;
  assign n3711 = n3709 & n3710 ;
  assign n3712 = n3709 | n3710 ;
  assign n3713 = ~n3711 & n3712 ;
  assign n3714 = n2784 & ~n3008 ;
  assign n3715 = ~n2541 & n2786 ;
  assign n3716 = n2544 & n2791 ;
  assign n3717 = n2549 & n2794 ;
  assign n3718 = n3716 | n3717 ;
  assign n3719 = n3715 | n3718 ;
  assign n3720 = n3714 | n3719 ;
  assign n3721 = n906 & ~n3720 ;
  assign n3722 = ~n906 & n3720 ;
  assign n3723 = n3721 | n3722 ;
  assign n3724 = n3713 & n3723 ;
  assign n3725 = n3713 | n3723 ;
  assign n3726 = ~n3724 & n3725 ;
  assign n3727 = n3679 & n3726 ;
  assign n3728 = n3240 | n3726 ;
  assign n3729 = n3243 | n3728 ;
  assign n3730 = ~n3727 & n3729 ;
  assign n3731 = ~n2521 & n2976 ;
  assign n3732 = n2538 & n2982 ;
  assign n3733 = n2618 & n2984 ;
  assign n3734 = n3732 | n3733 ;
  assign n3735 = n3731 | n3734 ;
  assign n3736 = n2988 & ~n3296 ;
  assign n3737 = n3735 | n3736 ;
  assign n3738 = n1190 | n3737 ;
  assign n3739 = n1190 & n3737 ;
  assign n3740 = n3738 & ~n3739 ;
  assign n3741 = n3730 | n3740 ;
  assign n3742 = n3729 & n3740 ;
  assign n3743 = ~n3727 & n3742 ;
  assign n3744 = n3741 & ~n3743 ;
  assign n3745 = n3678 & n3744 ;
  assign n3746 = n3678 | n3744 ;
  assign n3747 = ~n3745 & n3746 ;
  assign n3748 = n3677 & n3747 ;
  assign n3749 = n3677 | n3747 ;
  assign n3750 = ~n3748 & n3749 ;
  assign n3751 = n3633 & n3750 ;
  assign n3752 = n3267 | n3750 ;
  assign n3753 = n3507 | n3752 ;
  assign n3754 = ~n3751 & n3753 ;
  assign n3755 = n618 | n1322 ;
  assign n3756 = n970 | n3526 ;
  assign n3757 = n3755 | n3756 ;
  assign n3758 = n2174 | n3757 ;
  assign n3759 = n3511 | n3758 ;
  assign n3760 = n418 | n3759 ;
  assign n3761 = n439 | n3760 ;
  assign n3762 = n135 | n654 ;
  assign n3763 = n312 | n3762 ;
  assign n3764 = n3761 | n3763 ;
  assign n3765 = n3754 | n3764 ;
  assign n3766 = n3753 & n3764 ;
  assign n3767 = ~n3751 & n3766 ;
  assign n3768 = n3765 & ~n3767 ;
  assign n3769 = n3632 & n3768 ;
  assign n3770 = n3632 | n3768 ;
  assign n3771 = ~n3769 & n3770 ;
  assign n3772 = n3631 & n3771 ;
  assign n3773 = n3631 | n3771 ;
  assign n3774 = ~n3772 & n3773 ;
  assign n3775 = pi22 & ~pi23 ;
  assign n3776 = ~pi22 & pi23 ;
  assign n3777 = n3775 | n3776 ;
  assign n3778 = n3774 & n3777 ;
  assign n3779 = n3767 | n3769 ;
  assign n3780 = n3748 | n3751 ;
  assign n3781 = n229 | n274 ;
  assign n3782 = n2035 | n2086 ;
  assign n3783 = n289 | n341 ;
  assign n3784 = n2304 | n3783 ;
  assign n3785 = n3782 | n3784 ;
  assign n3786 = n320 | n3785 ;
  assign n3787 = n3781 | n3786 ;
  assign n3788 = n504 | n804 ;
  assign n3789 = n628 | n3788 ;
  assign n3790 = n1339 & ~n3789 ;
  assign n3791 = ~n3787 & n3790 ;
  assign n3792 = n858 | n2303 ;
  assign n3793 = n3791 & ~n3792 ;
  assign n3794 = ~n317 & n3793 ;
  assign n3795 = n238 | n401 ;
  assign n3796 = n263 | n3795 ;
  assign n3797 = n3794 & ~n3796 ;
  assign n3798 = n3654 | n3797 ;
  assign n3799 = n3654 & n3797 ;
  assign n3800 = n3798 & ~n3799 ;
  assign n3801 = n3656 | n3800 ;
  assign n3802 = n3656 & n3800 ;
  assign n3803 = n3801 & ~n3802 ;
  assign n3804 = ~n3663 & n3664 ;
  assign n3805 = ( n2511 & n2533 ) | ( n2511 & ~n3656 ) | ( n2533 & ~n3656 );
  assign n3806 = ( n2633 & ~n3804 ) | ( n2633 & n3805 ) | ( ~n3804 & n3805 );
  assign n3807 = ( n2632 & ~n3804 ) | ( n2632 & n3805 ) | ( ~n3804 & n3805 );
  assign n3808 = ( n2628 & n3806 ) | ( n2628 & n3807 ) | ( n3806 & n3807 );
  assign n3809 = n3803 | n3808 ;
  assign n3810 = n3803 & n3808 ;
  assign n3811 = n3809 & ~n3810 ;
  assign n3812 = n2531 & n3811 ;
  assign n3813 = n2518 & ~n3800 ;
  assign n3814 = n2511 & n2522 ;
  assign n3815 = n2527 & ~n3656 ;
  assign n3816 = n3814 | n3815 ;
  assign n3817 = n3813 | n3816 ;
  assign n3818 = n3812 | n3817 ;
  assign n3819 = n32 & ~n3818 ;
  assign n3820 = ~n32 & n3818 ;
  assign n3821 = n3819 | n3820 ;
  assign n3822 = n3743 | n3745 ;
  assign n3823 = n3724 | n3727 ;
  assign n3824 = n3707 | n3711 ;
  assign n3825 = n224 & ~n2569 ;
  assign n3826 = n2558 & n2651 ;
  assign n3827 = n2566 & n2745 ;
  assign n3828 = n2561 & n2649 ;
  assign n3829 = n3827 | n3828 ;
  assign n3830 = n3826 | n3829 ;
  assign n3831 = n2657 & n2821 ;
  assign n3832 = n3830 | n3831 ;
  assign n3833 = n3825 & n3832 ;
  assign n3834 = n3825 | n3832 ;
  assign n3835 = ~n3833 & n3834 ;
  assign n3836 = n224 & ~n3687 ;
  assign n3837 = ~n2572 & n3836 ;
  assign n3838 = n3694 | n3837 ;
  assign n3839 = n3835 & n3838 ;
  assign n3840 = n3835 | n3838 ;
  assign n3841 = ~n3839 & n3840 ;
  assign n3842 = n2549 & n2680 ;
  assign n3843 = ~n2555 & n2676 ;
  assign n3844 = n2552 & n2678 ;
  assign n3845 = n3843 | n3844 ;
  assign n3846 = n3842 | n3845 ;
  assign n3847 = n2684 & n2953 ;
  assign n3848 = n3846 | n3847 ;
  assign n3849 = n375 | n3848 ;
  assign n3850 = n375 & n3848 ;
  assign n3851 = n3849 & ~n3850 ;
  assign n3852 = n3841 & n3851 ;
  assign n3853 = n3841 | n3851 ;
  assign n3854 = ~n3852 & n3853 ;
  assign n3855 = n3824 & n3854 ;
  assign n3856 = n3824 | n3854 ;
  assign n3857 = ~n3855 & n3856 ;
  assign n3858 = n2784 & ~n2991 ;
  assign n3859 = n2538 & n2786 ;
  assign n3860 = n2544 & n2794 ;
  assign n3861 = ~n2541 & n2791 ;
  assign n3862 = n3860 | n3861 ;
  assign n3863 = n3859 | n3862 ;
  assign n3864 = n3858 | n3863 ;
  assign n3865 = n906 & ~n3864 ;
  assign n3866 = ~n906 & n3864 ;
  assign n3867 = n3865 | n3866 ;
  assign n3868 = n3857 & n3867 ;
  assign n3869 = n3857 | n3867 ;
  assign n3870 = ~n3868 & n3869 ;
  assign n3871 = n3823 & n3870 ;
  assign n3872 = n3724 | n3870 ;
  assign n3873 = n3727 | n3872 ;
  assign n3874 = ~n3871 & n3873 ;
  assign n3875 = n2526 & n2976 ;
  assign n3876 = n2618 & n2982 ;
  assign n3877 = ~n2521 & n2984 ;
  assign n3878 = n3876 | n3877 ;
  assign n3879 = n3875 | n3878 ;
  assign n3880 = n2988 & ~n3280 ;
  assign n3881 = n3879 | n3880 ;
  assign n3882 = n1190 | n3881 ;
  assign n3883 = n1190 & n3881 ;
  assign n3884 = n3882 & ~n3883 ;
  assign n3885 = n3874 | n3884 ;
  assign n3886 = n3873 & n3884 ;
  assign n3887 = ~n3871 & n3886 ;
  assign n3888 = n3885 & ~n3887 ;
  assign n3889 = n3822 & n3888 ;
  assign n3890 = n3822 | n3888 ;
  assign n3891 = ~n3889 & n3890 ;
  assign n3892 = n3821 & n3891 ;
  assign n3893 = n3821 | n3891 ;
  assign n3894 = ~n3892 & n3893 ;
  assign n3895 = n3780 & n3894 ;
  assign n3896 = n3748 | n3894 ;
  assign n3897 = n3751 | n3896 ;
  assign n3898 = ~n3895 & n3897 ;
  assign n3899 = n2136 | n2194 ;
  assign n3900 = n434 | n3899 ;
  assign n3901 = n2035 | n3900 ;
  assign n3902 = n121 | n209 ;
  assign n3903 = n1320 | n3902 ;
  assign n3904 = n3901 | n3903 ;
  assign n3905 = n2432 | n3511 ;
  assign n3906 = n3538 | n3905 ;
  assign n3907 = n3904 | n3906 ;
  assign n3908 = n185 | n3907 ;
  assign n3909 = n176 | n3908 ;
  assign n3910 = n201 | n3909 ;
  assign n3911 = n234 | n320 ;
  assign n3912 = n247 | n3911 ;
  assign n3913 = n3910 | n3912 ;
  assign n3914 = n3898 | n3913 ;
  assign n3915 = n3897 & n3913 ;
  assign n3916 = ~n3895 & n3915 ;
  assign n3917 = n3914 & ~n3916 ;
  assign n3918 = n3779 & n3917 ;
  assign n3919 = n3779 | n3917 ;
  assign n3920 = ~n3918 & n3919 ;
  assign n3921 = n3772 & n3920 ;
  assign n3922 = n3772 | n3920 ;
  assign n3923 = ~n3921 & n3922 ;
  assign n3924 = n3778 & ~n3923 ;
  assign n3925 = ~n3778 & n3923 ;
  assign n3926 = n3924 | n3925 ;
  assign n3927 = n3774 | n3923 ;
  assign n3928 = n3777 & n3927 ;
  assign n3929 = n3916 | n3918 ;
  assign n3930 = n273 | n331 ;
  assign n3931 = n138 | n607 ;
  assign n3932 = n3616 | n3931 ;
  assign n3933 = n129 | n194 ;
  assign n3934 = n106 | n3933 ;
  assign n3935 = n285 | n447 ;
  assign n3936 = n1995 | n3935 ;
  assign n3937 = n3934 | n3936 ;
  assign n3938 = n424 | n3937 ;
  assign n3939 = n3932 | n3938 ;
  assign n3940 = n205 | n3939 ;
  assign n3941 = n291 | n3940 ;
  assign n3942 = n328 | n401 ;
  assign n3943 = n3941 | n3942 ;
  assign n3944 = n335 | n3943 ;
  assign n3945 = n3930 | n3944 ;
  assign n3946 = n3892 | n3895 ;
  assign n3947 = n2522 & ~n3656 ;
  assign n3948 = n2527 & ~n3800 ;
  assign n3949 = n3947 | n3948 ;
  assign n3950 = ( n3800 & n3801 ) | ( n3800 & ~n3810 ) | ( n3801 & ~n3810 );
  assign n3951 = n3800 & ~n3810 ;
  assign n3952 = n3950 & ~n3951 ;
  assign n3953 = n2531 & n3952 ;
  assign n3954 = n3949 | n3953 ;
  assign n3955 = n32 & ~n3954 ;
  assign n3956 = ~n32 & n3954 ;
  assign n3957 = n3955 | n3956 ;
  assign n3958 = n3887 | n3889 ;
  assign n3959 = n3868 | n3871 ;
  assign n3960 = n3852 | n3855 ;
  assign n3961 = n224 & ~n2566 ;
  assign n3962 = ~n2555 & n2651 ;
  assign n3963 = n2561 & n2745 ;
  assign n3964 = n2558 & n2649 ;
  assign n3965 = n3963 | n3964 ;
  assign n3966 = n3962 | n3965 ;
  assign n3967 = n2657 & ~n2806 ;
  assign n3968 = n3966 | n3967 ;
  assign n3969 = n3961 & n3968 ;
  assign n3970 = n3961 | n3968 ;
  assign n3971 = ~n3969 & n3970 ;
  assign n3972 = n224 & ~n3832 ;
  assign n3973 = n2569 & n3972 ;
  assign n3974 = n3839 | n3973 ;
  assign n3975 = n3971 & n3974 ;
  assign n3976 = n3971 | n3974 ;
  assign n3977 = ~n3975 & n3976 ;
  assign n3978 = n2544 & n2680 ;
  assign n3979 = n2552 & n2676 ;
  assign n3980 = n2549 & n2678 ;
  assign n3981 = n3979 | n3980 ;
  assign n3982 = n3978 | n3981 ;
  assign n3983 = n2684 & n3020 ;
  assign n3984 = n3982 | n3983 ;
  assign n3985 = n375 | n3984 ;
  assign n3986 = n375 & n3984 ;
  assign n3987 = n3985 & ~n3986 ;
  assign n3988 = n3977 & n3987 ;
  assign n3989 = n3977 | n3987 ;
  assign n3990 = ~n3988 & n3989 ;
  assign n3991 = n3960 & n3990 ;
  assign n3992 = n3960 | n3990 ;
  assign n3993 = ~n3991 & n3992 ;
  assign n3994 = n2618 & n2786 ;
  assign n3995 = ~n2541 & n2794 ;
  assign n3996 = n2538 & n2791 ;
  assign n3997 = n3995 | n3996 ;
  assign n3998 = n3994 | n3997 ;
  assign n3999 = n2784 & n3254 ;
  assign n4000 = n3998 | n3999 ;
  assign n4001 = n906 & ~n4000 ;
  assign n4002 = ~n906 & n4000 ;
  assign n4003 = n4001 | n4002 ;
  assign n4004 = n3993 & n4003 ;
  assign n4005 = n3993 | n4003 ;
  assign n4006 = ~n4004 & n4005 ;
  assign n4007 = n3959 & n4006 ;
  assign n4008 = n3868 | n4006 ;
  assign n4009 = n3871 | n4008 ;
  assign n4010 = ~n4007 & n4009 ;
  assign n4011 = n2511 & n2976 ;
  assign n4012 = ~n2521 & n2982 ;
  assign n4013 = n2526 & n2984 ;
  assign n4014 = n4012 | n4013 ;
  assign n4015 = n4011 | n4014 ;
  assign n4016 = n2635 & n2988 ;
  assign n4017 = n4015 | n4016 ;
  assign n4018 = n1190 | n4017 ;
  assign n4019 = n1190 & n4017 ;
  assign n4020 = n4018 & ~n4019 ;
  assign n4021 = n4010 | n4020 ;
  assign n4022 = n4009 & n4020 ;
  assign n4023 = ~n4007 & n4022 ;
  assign n4024 = n4021 & ~n4023 ;
  assign n4025 = n3958 & n4024 ;
  assign n4026 = n3958 | n4024 ;
  assign n4027 = ~n4025 & n4026 ;
  assign n4028 = n3957 & n4027 ;
  assign n4029 = n3957 | n4027 ;
  assign n4030 = ~n4028 & n4029 ;
  assign n4031 = n3946 & n4030 ;
  assign n4032 = n3946 | n4030 ;
  assign n4033 = ~n4031 & n4032 ;
  assign n4034 = n3945 | n4033 ;
  assign n4035 = n3945 & n4033 ;
  assign n4036 = n4034 & ~n4035 ;
  assign n4037 = n3929 & n4036 ;
  assign n4038 = n3929 | n4036 ;
  assign n4039 = ~n4037 & n4038 ;
  assign n4040 = n3921 & n4039 ;
  assign n4041 = n3921 | n4039 ;
  assign n4042 = ~n4040 & n4041 ;
  assign n4043 = n3928 & ~n4042 ;
  assign n4044 = ~n3928 & n4042 ;
  assign n4045 = n4043 | n4044 ;
  assign n4046 = n3927 | n4042 ;
  assign n4047 = n3777 & n4046 ;
  assign n4048 = n4035 | n4037 ;
  assign n4049 = n185 | n296 ;
  assign n4050 = n2194 | n3581 ;
  assign n4051 = n830 | n4050 ;
  assign n4052 = n661 | n1331 ;
  assign n4053 = n4051 | n4052 ;
  assign n4054 = n462 | n2056 ;
  assign n4055 = n202 | n4054 ;
  assign n4056 = n4053 | n4055 ;
  assign n4057 = n4049 | n4056 ;
  assign n4058 = n405 | n4057 ;
  assign n4059 = n269 | n4058 ;
  assign n4060 = n503 | n4059 ;
  assign n4061 = n622 | n4060 ;
  assign n4062 = n4028 | n4031 ;
  assign n4063 = n4023 | n4025 ;
  assign n4064 = n4004 | n4007 ;
  assign n4065 = n3988 | n3991 ;
  assign n4066 = n224 & ~n2561 ;
  assign n4067 = n2552 & n2651 ;
  assign n4068 = n2558 & n2745 ;
  assign n4069 = ~n2555 & n2649 ;
  assign n4070 = n4068 | n4069 ;
  assign n4071 = n4067 | n4070 ;
  assign n4072 = n2657 & ~n2777 ;
  assign n4073 = n4071 | n4072 ;
  assign n4074 = n4066 & n4073 ;
  assign n4075 = n4066 | n4073 ;
  assign n4076 = ~n4074 & n4075 ;
  assign n4077 = n224 & ~n3968 ;
  assign n4078 = n2566 & n4077 ;
  assign n4079 = n3975 | n4078 ;
  assign n4080 = n4076 & n4079 ;
  assign n4081 = n4076 | n4079 ;
  assign n4082 = ~n4080 & n4081 ;
  assign n4083 = ~n2541 & n2680 ;
  assign n4084 = n2549 & n2676 ;
  assign n4085 = n2544 & n2678 ;
  assign n4086 = n4084 | n4085 ;
  assign n4087 = n4083 | n4086 ;
  assign n4088 = n2684 & ~n3008 ;
  assign n4089 = n4087 | n4088 ;
  assign n4090 = n375 | n4089 ;
  assign n4091 = n375 & n4089 ;
  assign n4092 = n4090 & ~n4091 ;
  assign n4093 = n4082 & n4092 ;
  assign n4094 = n4082 | n4092 ;
  assign n4095 = ~n4093 & n4094 ;
  assign n4096 = n4065 & n4095 ;
  assign n4097 = n4065 | n4095 ;
  assign n4098 = ~n4096 & n4097 ;
  assign n4099 = ~n2521 & n2786 ;
  assign n4100 = n2538 & n2794 ;
  assign n4101 = n2618 & n2791 ;
  assign n4102 = n4100 | n4101 ;
  assign n4103 = n4099 | n4102 ;
  assign n4104 = n2784 & ~n3296 ;
  assign n4105 = n4103 | n4104 ;
  assign n4106 = n906 & ~n4105 ;
  assign n4107 = ~n906 & n4105 ;
  assign n4108 = n4106 | n4107 ;
  assign n4109 = n4098 & n4108 ;
  assign n4110 = n4098 | n4108 ;
  assign n4111 = ~n4109 & n4110 ;
  assign n4112 = n4064 & n4111 ;
  assign n4113 = n4004 | n4111 ;
  assign n4114 = n4007 | n4113 ;
  assign n4115 = ~n4112 & n4114 ;
  assign n4116 = n2988 & ~n3669 ;
  assign n4117 = n2988 & n3671 ;
  assign n4118 = ( ~n3670 & n4116 ) | ( ~n3670 & n4117 ) | ( n4116 & n4117 );
  assign n4119 = n2976 & ~n3656 ;
  assign n4120 = n2526 & n2982 ;
  assign n4121 = n2511 & n2984 ;
  assign n4122 = n4120 | n4121 ;
  assign n4123 = n4119 | n4122 ;
  assign n4124 = n1190 | n4123 ;
  assign n4125 = n4118 | n4124 ;
  assign n4126 = n1190 & n4123 ;
  assign n4127 = ( n1190 & n4118 ) | ( n1190 & n4126 ) | ( n4118 & n4126 );
  assign n4128 = n4125 & ~n4127 ;
  assign n4129 = n4115 | n4128 ;
  assign n4130 = n4114 & n4128 ;
  assign n4131 = ~n4112 & n4130 ;
  assign n4132 = n4129 & ~n4131 ;
  assign n4133 = n2522 & ~n3800 ;
  assign n4134 = n2531 & ~n3950 ;
  assign n4135 = n4133 | n4134 ;
  assign n4136 = n32 & ~n4135 ;
  assign n4137 = ~n32 & n4135 ;
  assign n4138 = n4136 | n4137 ;
  assign n4139 = n4132 | n4138 ;
  assign n4140 = ~n4131 & n4138 ;
  assign n4141 = n4129 & n4140 ;
  assign n4142 = n4139 & ~n4141 ;
  assign n4143 = n4063 | n4142 ;
  assign n4144 = n4063 & ~n4141 ;
  assign n4145 = n4139 & n4144 ;
  assign n4146 = n4143 & ~n4145 ;
  assign n4147 = n4062 & n4146 ;
  assign n4148 = n4062 | n4146 ;
  assign n4149 = ~n4147 & n4148 ;
  assign n4150 = n4061 | n4149 ;
  assign n4151 = n4061 & n4149 ;
  assign n4152 = n4150 & ~n4151 ;
  assign n4153 = n4048 & n4152 ;
  assign n4154 = n4048 | n4152 ;
  assign n4155 = ~n4153 & n4154 ;
  assign n4156 = n4040 & n4155 ;
  assign n4157 = n4040 | n4155 ;
  assign n4158 = ~n4156 & n4157 ;
  assign n4159 = n4047 & ~n4158 ;
  assign n4160 = ~n4047 & n4158 ;
  assign n4161 = n4159 | n4160 ;
  assign n4162 = n4151 | n4153 ;
  assign n4163 = n322 | n382 ;
  assign n4164 = n654 | n2111 ;
  assign n4165 = n2331 | n4164 ;
  assign n4166 = n4163 | n4165 ;
  assign n4167 = n146 | n2326 ;
  assign n4168 = n293 | n4167 ;
  assign n4169 = n209 | n2321 ;
  assign n4170 = n4168 | n4169 ;
  assign n4171 = n290 | n2334 ;
  assign n4172 = n447 | n4171 ;
  assign n4173 = n4170 | n4172 ;
  assign n4174 = n4166 | n4173 ;
  assign n4175 = n381 | n4174 ;
  assign n4176 = n892 | n1319 ;
  assign n4177 = n181 | n4176 ;
  assign n4178 = n649 | n4177 ;
  assign n4179 = n4175 | n4178 ;
  assign n4180 = n177 | n4179 ;
  assign n4181 = n483 | n4180 ;
  assign n4182 = n4145 | n4147 ;
  assign n4183 = n4131 | n4141 ;
  assign n4184 = n4093 | n4096 ;
  assign n4185 = n224 & ~n4073 ;
  assign n4186 = n2561 & n4185 ;
  assign n4187 = n4080 | n4186 ;
  assign n4188 = n2549 & n2651 ;
  assign n4189 = ~n2555 & n2745 ;
  assign n4190 = n2552 & n2649 ;
  assign n4191 = n4189 | n4190 ;
  assign n4192 = n4188 | n4191 ;
  assign n4193 = n2657 & n2953 ;
  assign n4194 = n4192 | n4193 ;
  assign n4195 = n224 & ~n4194 ;
  assign n4196 = n224 & ~n4195 ;
  assign n4197 = ( n4194 & n4195 ) | ( n4194 & ~n4196 ) | ( n4195 & ~n4196 );
  assign n4198 = n32 & n224 ;
  assign n4199 = n2558 & n4198 ;
  assign n4200 = n32 & ~n4199 ;
  assign n4201 = n2558 & ~n4199 ;
  assign n4202 = n224 & n4201 ;
  assign n4203 = n4200 | n4202 ;
  assign n4204 = n4197 & n4203 ;
  assign n4205 = n4197 & ~n4204 ;
  assign n4206 = n4203 & ~n4204 ;
  assign n4207 = n4205 | n4206 ;
  assign n4208 = n4187 & ~n4207 ;
  assign n4209 = ~n4187 & n4207 ;
  assign n4210 = n4208 | n4209 ;
  assign n4211 = n2538 & n2680 ;
  assign n4212 = n2544 & n2676 ;
  assign n4213 = ~n2541 & n2678 ;
  assign n4214 = n4212 | n4213 ;
  assign n4215 = n4211 | n4214 ;
  assign n4216 = n2684 & ~n2991 ;
  assign n4217 = n4215 | n4216 ;
  assign n4218 = n375 & n4217 ;
  assign n4219 = n375 | n4217 ;
  assign n4220 = ~n4218 & n4219 ;
  assign n4221 = n4210 & n4220 ;
  assign n4222 = n4210 | n4220 ;
  assign n4223 = ~n4221 & n4222 ;
  assign n4224 = n4184 & n4223 ;
  assign n4225 = n4184 | n4223 ;
  assign n4226 = ~n4224 & n4225 ;
  assign n4227 = n2526 & n2786 ;
  assign n4228 = n2618 & n2794 ;
  assign n4229 = ~n2521 & n2791 ;
  assign n4230 = n4228 | n4229 ;
  assign n4231 = n4227 | n4230 ;
  assign n4232 = n2784 & ~n3277 ;
  assign n4233 = ~n2526 & n2784 ;
  assign n4234 = ( n3279 & n4232 ) | ( n3279 & n4233 ) | ( n4232 & n4233 );
  assign n4235 = n4231 | n4234 ;
  assign n4236 = n906 & ~n4231 ;
  assign n4237 = ~n4234 & n4236 ;
  assign n4238 = n906 & ~n4236 ;
  assign n4239 = ( n906 & n4234 ) | ( n906 & n4238 ) | ( n4234 & n4238 );
  assign n4240 = ( n4235 & n4237 ) | ( n4235 & ~n4239 ) | ( n4237 & ~n4239 );
  assign n4241 = n4226 & n4240 ;
  assign n4242 = n4226 | n4240 ;
  assign n4243 = ~n4241 & n4242 ;
  assign n4244 = n4109 | n4112 ;
  assign n4245 = n4243 & n4244 ;
  assign n4246 = n4243 | n4244 ;
  assign n4247 = ~n4245 & n4246 ;
  assign n4248 = n2976 & ~n3800 ;
  assign n4249 = n2511 & n2982 ;
  assign n4250 = n2984 & ~n3656 ;
  assign n4251 = n4249 | n4250 ;
  assign n4252 = n4248 | n4251 ;
  assign n4253 = n2988 & n3811 ;
  assign n4254 = n4252 | n4253 ;
  assign n4255 = n1190 & n4254 ;
  assign n4256 = n1190 | n4254 ;
  assign n4257 = ~n4255 & n4256 ;
  assign n4258 = n4247 & n4257 ;
  assign n4259 = n4247 | n4257 ;
  assign n4260 = ~n4258 & n4259 ;
  assign n4261 = n4183 & n4260 ;
  assign n4262 = n4183 | n4260 ;
  assign n4263 = ~n4261 & n4262 ;
  assign n4264 = n4182 & n4263 ;
  assign n4265 = n4145 | n4263 ;
  assign n4266 = n4147 | n4265 ;
  assign n4267 = ~n4264 & n4266 ;
  assign n4268 = n4181 | n4267 ;
  assign n4269 = n4181 & n4267 ;
  assign n4270 = n4268 & ~n4269 ;
  assign n4271 = n4162 & n4270 ;
  assign n4272 = n4162 | n4270 ;
  assign n4273 = ~n4271 & n4272 ;
  assign n4274 = n4156 | n4273 ;
  assign n4275 = n4156 & n4273 ;
  assign n4276 = n4274 & ~n4275 ;
  assign n4277 = n4046 | n4158 ;
  assign n4278 = n3777 & n4277 ;
  assign n4279 = ~n4276 & n4278 ;
  assign n4280 = n4276 & ~n4278 ;
  assign n4281 = n4279 | n4280 ;
  assign n4282 = n4269 | n4271 ;
  assign n4283 = n158 | n181 ;
  assign n4284 = n251 | n2444 ;
  assign n4285 = n255 | n4284 ;
  assign n4286 = n153 | n608 ;
  assign n4287 = n206 | n4286 ;
  assign n4288 = n264 | n405 ;
  assign n4289 = n314 | n4288 ;
  assign n4290 = n2164 | n4289 ;
  assign n4291 = n3787 | n4290 ;
  assign n4292 = n4287 | n4291 ;
  assign n4293 = n3903 | n4292 ;
  assign n4294 = n4285 | n4293 ;
  assign n4295 = n128 | n4294 ;
  assign n4296 = n4283 | n4295 ;
  assign n4297 = n1981 | n4296 ;
  assign n4298 = n513 | n4297 ;
  assign n4299 = n4261 | n4264 ;
  assign n4300 = n4245 | n4258 ;
  assign n4301 = n4224 | n4241 ;
  assign n4302 = n4187 & n4207 ;
  assign n4303 = n4221 | n4302 ;
  assign n4304 = n4199 | n4204 ;
  assign n4305 = ~n2555 & n4198 ;
  assign n4306 = n32 & ~n4305 ;
  assign n4307 = n2555 | n4305 ;
  assign n4308 = n224 & ~n4307 ;
  assign n4309 = n4306 | n4308 ;
  assign n4310 = n4304 & n4309 ;
  assign n4311 = n4304 & ~n4310 ;
  assign n4312 = n4309 & ~n4310 ;
  assign n4313 = n4311 | n4312 ;
  assign n4314 = n2544 & n2651 ;
  assign n4315 = n2552 & n2745 ;
  assign n4316 = n2549 & n2649 ;
  assign n4317 = n4315 | n4316 ;
  assign n4318 = n4314 | n4317 ;
  assign n4319 = n2657 & n3020 ;
  assign n4320 = n4318 | n4319 ;
  assign n4321 = n224 | n4320 ;
  assign n4322 = n224 & n4320 ;
  assign n4323 = n4321 & ~n4322 ;
  assign n4324 = n4313 & n4323 ;
  assign n4325 = n4313 | n4323 ;
  assign n4326 = ~n4324 & n4325 ;
  assign n4327 = n2618 & n2680 ;
  assign n4328 = ~n2541 & n2676 ;
  assign n4329 = n2538 & n2678 ;
  assign n4330 = n4328 | n4329 ;
  assign n4331 = n4327 | n4330 ;
  assign n4332 = n2684 & n3254 ;
  assign n4333 = n4331 | n4332 ;
  assign n4334 = n375 & ~n4333 ;
  assign n4335 = ~n375 & n4333 ;
  assign n4336 = n4334 | n4335 ;
  assign n4337 = n4326 & n4336 ;
  assign n4338 = n4326 | n4336 ;
  assign n4339 = ~n4337 & n4338 ;
  assign n4340 = n4303 & n4339 ;
  assign n4341 = n4303 | n4339 ;
  assign n4342 = ~n4340 & n4341 ;
  assign n4343 = n2511 & n2786 ;
  assign n4344 = ~n2521 & n2794 ;
  assign n4345 = n2526 & n2791 ;
  assign n4346 = n4344 | n4345 ;
  assign n4347 = n4343 | n4346 ;
  assign n4348 = n2635 & n2784 ;
  assign n4349 = n4347 | n4348 ;
  assign n4350 = n906 & ~n4349 ;
  assign n4351 = n906 & ~n4350 ;
  assign n4352 = ( n4349 & n4350 ) | ( n4349 & ~n4351 ) | ( n4350 & ~n4351 );
  assign n4353 = n4342 & n4352 ;
  assign n4354 = n4342 | n4352 ;
  assign n4355 = ~n4353 & n4354 ;
  assign n4356 = n4301 & n4355 ;
  assign n4357 = n4301 | n4355 ;
  assign n4358 = ~n4356 & n4357 ;
  assign n4359 = n2982 & ~n3656 ;
  assign n4360 = n2984 & ~n3800 ;
  assign n4361 = n4359 | n4360 ;
  assign n4362 = n2988 & n3952 ;
  assign n4363 = n4361 | n4362 ;
  assign n4364 = n1190 & ~n4363 ;
  assign n4365 = ~n1190 & n4363 ;
  assign n4366 = n4364 | n4365 ;
  assign n4367 = n4358 & n4366 ;
  assign n4368 = n4358 | n4366 ;
  assign n4369 = ~n4367 & n4368 ;
  assign n4370 = n4300 & n4369 ;
  assign n4371 = n4300 | n4369 ;
  assign n4372 = ~n4370 & n4371 ;
  assign n4373 = n4299 & n4372 ;
  assign n4374 = n4299 | n4372 ;
  assign n4375 = ~n4373 & n4374 ;
  assign n4376 = n4298 | n4375 ;
  assign n4377 = n4298 & n4375 ;
  assign n4378 = n4376 & ~n4377 ;
  assign n4379 = n4282 & n4378 ;
  assign n4380 = n4269 | n4378 ;
  assign n4381 = n4271 | n4380 ;
  assign n4382 = ~n4379 & n4381 ;
  assign n4383 = n4275 | n4382 ;
  assign n4384 = n4275 & n4382 ;
  assign n4385 = n4383 & ~n4384 ;
  assign n4386 = n4276 | n4277 ;
  assign n4387 = n3777 & n4386 ;
  assign n4388 = ~n4385 & n4387 ;
  assign n4389 = n4385 & ~n4387 ;
  assign n4390 = n4388 | n4389 ;
  assign n4391 = n4377 | n4379 ;
  assign n4392 = n885 | n2327 ;
  assign n4393 = n3542 | n4392 ;
  assign n4394 = n2487 | n4393 ;
  assign n4395 = n146 | n4394 ;
  assign n4396 = n507 | n4395 ;
  assign n4397 = n858 | n1981 ;
  assign n4398 = n1991 | n2194 ;
  assign n4399 = n804 | n2291 ;
  assign n4400 = n1010 | n4399 ;
  assign n4401 = n481 | n4400 ;
  assign n4402 = n4398 | n4401 ;
  assign n4403 = n4397 | n4402 ;
  assign n4404 = n330 | n4403 ;
  assign n4405 = n196 | n4404 ;
  assign n4406 = n2102 | n4405 ;
  assign n4407 = n4396 | n4406 ;
  assign n4408 = n4370 | n4373 ;
  assign n4409 = n4356 | n4367 ;
  assign n4410 = n4340 | n4353 ;
  assign n4411 = n2982 & ~n3800 ;
  assign n4412 = n2988 & ~n3950 ;
  assign n4413 = n4411 | n4412 ;
  assign n4414 = ~n1190 & n4413 ;
  assign n4415 = n1190 & ~n4413 ;
  assign n4416 = n4414 | n4415 ;
  assign n4417 = n4410 & n4416 ;
  assign n4418 = n4410 | n4416 ;
  assign n4419 = ~n4417 & n4418 ;
  assign n4420 = n4324 | n4337 ;
  assign n4421 = n4305 | n4310 ;
  assign n4422 = n2552 & n4198 ;
  assign n4423 = n32 & ~n4422 ;
  assign n4424 = n2552 & ~n4422 ;
  assign n4425 = n224 & n4424 ;
  assign n4426 = n4423 | n4425 ;
  assign n4427 = n4421 & n4426 ;
  assign n4428 = n4421 & ~n4427 ;
  assign n4429 = n4426 & ~n4427 ;
  assign n4430 = n4428 | n4429 ;
  assign n4431 = ~n2541 & n2651 ;
  assign n4432 = n2549 & n2745 ;
  assign n4433 = n2544 & n2649 ;
  assign n4434 = n4432 | n4433 ;
  assign n4435 = n4431 | n4434 ;
  assign n4436 = n2657 & ~n3008 ;
  assign n4437 = n4435 | n4436 ;
  assign n4438 = n224 | n4437 ;
  assign n4439 = n224 & n4437 ;
  assign n4440 = n4438 & ~n4439 ;
  assign n4441 = n4430 & n4440 ;
  assign n4442 = n4430 | n4440 ;
  assign n4443 = ~n4441 & n4442 ;
  assign n4444 = ~n2521 & n2680 ;
  assign n4445 = n2538 & n2676 ;
  assign n4446 = n2618 & n2678 ;
  assign n4447 = n4445 | n4446 ;
  assign n4448 = n4444 | n4447 ;
  assign n4449 = n2684 & ~n3296 ;
  assign n4450 = n4448 | n4449 ;
  assign n4451 = n375 & ~n4450 ;
  assign n4452 = ~n375 & n4450 ;
  assign n4453 = n4451 | n4452 ;
  assign n4454 = n4443 & n4453 ;
  assign n4455 = n4443 | n4453 ;
  assign n4456 = ~n4454 & n4455 ;
  assign n4457 = n4420 & n4456 ;
  assign n4458 = n4420 | n4456 ;
  assign n4459 = ~n4457 & n4458 ;
  assign n4460 = n2786 & ~n3656 ;
  assign n4461 = n2526 & n2794 ;
  assign n4462 = n2511 & n2791 ;
  assign n4463 = n4461 | n4462 ;
  assign n4464 = n4460 | n4463 ;
  assign n4465 = ( n2784 & ~n3672 ) | ( n2784 & n4464 ) | ( ~n3672 & n4464 );
  assign n4466 = ( n906 & n4464 ) | ( n906 & ~n4465 ) | ( n4464 & ~n4465 );
  assign n4467 = n4465 | n4466 ;
  assign n4468 = ~n4464 & n4466 ;
  assign n4469 = ( ~n906 & n4467 ) | ( ~n906 & n4468 ) | ( n4467 & n4468 );
  assign n4470 = n4459 & n4469 ;
  assign n4471 = n4459 | n4469 ;
  assign n4472 = ~n4470 & n4471 ;
  assign n4473 = n4419 & n4472 ;
  assign n4474 = n4419 | n4472 ;
  assign n4475 = ~n4473 & n4474 ;
  assign n4476 = n4409 & n4475 ;
  assign n4477 = n4409 | n4475 ;
  assign n4478 = ~n4476 & n4477 ;
  assign n4479 = n4408 & n4478 ;
  assign n4480 = n4408 | n4478 ;
  assign n4481 = ~n4479 & n4480 ;
  assign n4482 = n4407 | n4481 ;
  assign n4483 = n4407 & n4481 ;
  assign n4484 = n4482 & ~n4483 ;
  assign n4485 = n4391 & n4484 ;
  assign n4486 = n4377 | n4484 ;
  assign n4487 = n4379 | n4486 ;
  assign n4488 = ~n4485 & n4487 ;
  assign n4489 = n4384 & n4488 ;
  assign n4490 = n4384 | n4488 ;
  assign n4491 = ~n4489 & n4490 ;
  assign n4492 = n4385 | n4386 ;
  assign n4493 = n3777 & n4492 ;
  assign n4494 = ~n4491 & n4493 ;
  assign n4495 = n4491 & ~n4493 ;
  assign n4496 = n4494 | n4495 ;
  assign n4497 = n157 | n229 ;
  assign n4498 = n623 | n4289 ;
  assign n4499 = n106 | n4498 ;
  assign n4500 = n208 | n2088 ;
  assign n4501 = n233 | n4500 ;
  assign n4502 = n240 | n285 ;
  assign n4503 = n2018 | n4502 ;
  assign n4504 = n115 | n290 ;
  assign n4505 = n2001 | n4504 ;
  assign n4506 = n4503 | n4505 ;
  assign n4507 = n4501 | n4506 ;
  assign n4508 = n2085 | n3588 ;
  assign n4509 = n329 | n462 ;
  assign n4510 = n148 | n434 ;
  assign n4511 = n4509 | n4510 ;
  assign n4512 = n4508 | n4511 ;
  assign n4513 = n4507 | n4512 ;
  assign n4514 = n671 | n4513 ;
  assign n4515 = n2260 | n4514 ;
  assign n4516 = n4499 | n4515 ;
  assign n4517 = n4497 | n4516 ;
  assign n4518 = n177 | n4404 ;
  assign n4519 = n109 | n971 ;
  assign n4520 = n4518 | n4519 ;
  assign n4521 = n4517 | n4520 ;
  assign n4522 = n234 | n4521 ;
  assign n4523 = n4476 | n4479 ;
  assign n4524 = n4417 | n4473 ;
  assign n4525 = n4457 | n4470 ;
  assign n4526 = n2786 & ~n3800 ;
  assign n4527 = n2511 & n2794 ;
  assign n4528 = n2791 & ~n3656 ;
  assign n4529 = n4527 | n4528 ;
  assign n4530 = n4526 | n4529 ;
  assign n4531 = n2784 & n3811 ;
  assign n4532 = n4530 | n4531 ;
  assign n4533 = n906 | n4532 ;
  assign n4534 = n906 & n4532 ;
  assign n4535 = n4533 & ~n4534 ;
  assign n4536 = n4525 & n4535 ;
  assign n4537 = n4525 | n4535 ;
  assign n4538 = ~n4536 & n4537 ;
  assign n4539 = n4441 | n4454 ;
  assign n4540 = n2526 & n2680 ;
  assign n4541 = n2618 & n2676 ;
  assign n4542 = ~n2521 & n2678 ;
  assign n4543 = n4541 | n4542 ;
  assign n4544 = n4540 | n4543 ;
  assign n4545 = n2684 & ~n3280 ;
  assign n4546 = n4544 | n4545 ;
  assign n4547 = n375 | n4546 ;
  assign n4548 = n375 & n4546 ;
  assign n4549 = n4547 & ~n4548 ;
  assign n4550 = n224 & n2549 ;
  assign n4551 = n32 | n1190 ;
  assign n4552 = n32 & n1190 ;
  assign n4553 = n4551 & ~n4552 ;
  assign n4554 = n4550 & n4553 ;
  assign n4555 = n4550 | n4553 ;
  assign n4556 = ~n4554 & n4555 ;
  assign n4557 = n2538 & n2651 ;
  assign n4558 = n2544 & n2745 ;
  assign n4559 = ~n2541 & n2649 ;
  assign n4560 = n4558 | n4559 ;
  assign n4561 = n4557 | n4560 ;
  assign n4562 = n2657 & ~n2991 ;
  assign n4563 = n4561 | n4562 ;
  assign n4564 = n224 & ~n4563 ;
  assign n4565 = ~n224 & n4563 ;
  assign n4566 = n4564 | n4565 ;
  assign n4567 = n4556 & n4566 ;
  assign n4568 = n4556 | n4566 ;
  assign n4569 = ~n4567 & n4568 ;
  assign n4570 = n4422 | n4427 ;
  assign n4571 = n4569 & n4570 ;
  assign n4572 = n4569 | n4570 ;
  assign n4573 = ~n4571 & n4572 ;
  assign n4574 = n4549 & n4573 ;
  assign n4575 = n4549 | n4573 ;
  assign n4576 = ~n4574 & n4575 ;
  assign n4577 = n4539 & n4576 ;
  assign n4578 = n4539 | n4576 ;
  assign n4579 = ~n4577 & n4578 ;
  assign n4580 = n4538 & n4579 ;
  assign n4581 = n4538 | n4579 ;
  assign n4582 = ~n4580 & n4581 ;
  assign n4583 = n4524 & n4582 ;
  assign n4584 = n4524 | n4582 ;
  assign n4585 = ~n4583 & n4584 ;
  assign n4586 = n4523 & n4585 ;
  assign n4587 = n4523 | n4585 ;
  assign n4588 = ~n4586 & n4587 ;
  assign n4589 = n4522 & n4588 ;
  assign n4590 = n4522 | n4588 ;
  assign n4591 = ~n4589 & n4590 ;
  assign n4592 = n4483 | n4485 ;
  assign n4593 = n4591 & n4592 ;
  assign n4594 = n4591 | n4592 ;
  assign n4595 = ~n4593 & n4594 ;
  assign n4596 = n4489 & n4595 ;
  assign n4597 = n4489 | n4595 ;
  assign n4598 = ~n4596 & n4597 ;
  assign n4599 = n4491 | n4492 ;
  assign n4600 = n3777 & n4599 ;
  assign n4601 = ~n4598 & n4600 ;
  assign n4602 = n4598 & ~n4600 ;
  assign n4603 = n4601 | n4602 ;
  assign n4604 = n4589 | n4593 ;
  assign n4605 = n190 | n305 ;
  assign n4606 = n142 | n4605 ;
  assign n4607 = n477 | n2039 ;
  assign n4608 = n406 | n4607 ;
  assign n4609 = n204 | n4608 ;
  assign n4610 = n140 | n4609 ;
  assign n4611 = n4606 | n4610 ;
  assign n4612 = n269 | n4611 ;
  assign n4613 = n382 | n4612 ;
  assign n4614 = n3571 | n4613 ;
  assign n4615 = n861 | n2196 ;
  assign n4616 = n850 | n4615 ;
  assign n4617 = n4614 | n4616 ;
  assign n4618 = n200 | n401 ;
  assign n4619 = n129 | n4618 ;
  assign n4620 = n281 | n4619 ;
  assign n4621 = n2041 | n4620 ;
  assign n4622 = n4617 | n4621 ;
  assign n4623 = n230 | n4622 ;
  assign n4624 = n4536 | n4580 ;
  assign n4625 = n4574 | n4577 ;
  assign n4626 = n4567 | n4571 ;
  assign n4627 = n2618 & n2651 ;
  assign n4628 = ~n2541 & n2745 ;
  assign n4629 = n2538 & n2649 ;
  assign n4630 = n4628 | n4629 ;
  assign n4631 = n4627 | n4630 ;
  assign n4632 = n2657 & n3254 ;
  assign n4633 = n4631 | n4632 ;
  assign n4634 = n224 | n4633 ;
  assign n4635 = n224 & n4633 ;
  assign n4636 = n4634 & ~n4635 ;
  assign n4637 = n224 & n2544 ;
  assign n4638 = n4551 & ~n4554 ;
  assign n4639 = n4637 | n4638 ;
  assign n4640 = n4637 & n4638 ;
  assign n4641 = n4639 & ~n4640 ;
  assign n4642 = n4636 & n4641 ;
  assign n4643 = n4636 | n4641 ;
  assign n4644 = ~n4642 & n4643 ;
  assign n4645 = n4626 & n4644 ;
  assign n4646 = n4626 | n4644 ;
  assign n4647 = ~n4645 & n4646 ;
  assign n4648 = n2511 & n2680 ;
  assign n4649 = ~n2521 & n2676 ;
  assign n4650 = n2526 & n2678 ;
  assign n4651 = n4649 | n4650 ;
  assign n4652 = n4648 | n4651 ;
  assign n4653 = n2635 & n2684 ;
  assign n4654 = n4652 | n4653 ;
  assign n4655 = n375 & n4654 ;
  assign n4656 = n375 | n4654 ;
  assign n4657 = ~n4655 & n4656 ;
  assign n4658 = n4647 & n4657 ;
  assign n4659 = n4647 | n4657 ;
  assign n4660 = ~n4658 & n4659 ;
  assign n4661 = n4625 & n4660 ;
  assign n4662 = n4625 | n4660 ;
  assign n4663 = ~n4661 & n4662 ;
  assign n4664 = n2794 & ~n3656 ;
  assign n4665 = n2791 & ~n3800 ;
  assign n4666 = n4664 | n4665 ;
  assign n4667 = ( n2784 & n3952 ) | ( n2784 & n4666 ) | ( n3952 & n4666 );
  assign n4668 = ( n906 & n4666 ) | ( n906 & ~n4667 ) | ( n4666 & ~n4667 );
  assign n4669 = n4667 | n4668 ;
  assign n4670 = ~n4666 & n4668 ;
  assign n4671 = ( ~n906 & n4669 ) | ( ~n906 & n4670 ) | ( n4669 & n4670 );
  assign n4672 = n4663 & n4671 ;
  assign n4673 = n4663 | n4671 ;
  assign n4674 = ~n4672 & n4673 ;
  assign n4675 = n4624 & n4674 ;
  assign n4676 = n4624 | n4674 ;
  assign n4677 = ~n4675 & n4676 ;
  assign n4678 = n4583 | n4586 ;
  assign n4679 = n4677 & n4678 ;
  assign n4680 = n4677 | n4678 ;
  assign n4681 = ~n4679 & n4680 ;
  assign n4682 = n4623 | n4681 ;
  assign n4683 = n4623 & n4681 ;
  assign n4684 = n4682 & ~n4683 ;
  assign n4685 = n4604 & n4684 ;
  assign n4686 = n4604 | n4684 ;
  assign n4687 = ~n4685 & n4686 ;
  assign n4688 = n4596 | n4687 ;
  assign n4689 = n4596 & n4687 ;
  assign n4690 = n4688 & ~n4689 ;
  assign n4691 = n4598 | n4599 ;
  assign n4692 = n3777 & n4691 ;
  assign n4693 = ~n4690 & n4692 ;
  assign n4694 = n4690 & ~n4692 ;
  assign n4695 = n4693 | n4694 ;
  assign n4696 = n4683 | n4685 ;
  assign n4697 = n196 | n2303 ;
  assign n4698 = n312 | n623 ;
  assign n4699 = n192 | n4698 ;
  assign n4700 = n675 | n4699 ;
  assign n4701 = n3520 | n4700 ;
  assign n4702 = n2487 | n4701 ;
  assign n4703 = n2432 | n4702 ;
  assign n4704 = n4697 | n4703 ;
  assign n4705 = n313 | n4704 ;
  assign n4706 = n142 | n4705 ;
  assign n4707 = n3588 | n4706 ;
  assign n4708 = n243 | n4707 ;
  assign n4709 = n336 | n4708 ;
  assign n4710 = n4675 | n4679 ;
  assign n4711 = n4661 | n4672 ;
  assign n4712 = n4645 | n4658 ;
  assign n4713 = n2794 & ~n3800 ;
  assign n4714 = n2784 & ~n3950 ;
  assign n4715 = n4713 | n4714 ;
  assign n4716 = n906 & ~n4715 ;
  assign n4717 = ~n906 & n4715 ;
  assign n4718 = n4716 | n4717 ;
  assign n4719 = n4712 & n4718 ;
  assign n4720 = n4712 | n4718 ;
  assign n4721 = ~n4719 & n4720 ;
  assign n4722 = n4639 & ~n4642 ;
  assign n4723 = n224 & ~n2547 ;
  assign n4724 = ~n2521 & n2651 ;
  assign n4725 = n2538 & n2745 ;
  assign n4726 = n2618 & n2649 ;
  assign n4727 = n4725 | n4726 ;
  assign n4728 = n4724 | n4727 ;
  assign n4729 = n2657 & ~n3296 ;
  assign n4730 = n4728 | n4729 ;
  assign n4731 = n224 & ~n4730 ;
  assign n4732 = ~n224 & n4730 ;
  assign n4733 = n4731 | n4732 ;
  assign n4734 = ~n4723 & n4733 ;
  assign n4735 = n4723 & ~n4733 ;
  assign n4736 = n4734 | n4735 ;
  assign n4737 = n4722 | n4736 ;
  assign n4738 = n4722 & n4736 ;
  assign n4739 = n4737 & ~n4738 ;
  assign n4740 = n2680 & ~n3656 ;
  assign n4741 = n2526 & n2676 ;
  assign n4742 = n2511 & n2678 ;
  assign n4743 = n4741 | n4742 ;
  assign n4744 = n4740 | n4743 ;
  assign n4745 = n2684 & ~n3672 ;
  assign n4746 = n4744 | n4745 ;
  assign n4747 = n375 & ~n4746 ;
  assign n4748 = ~n375 & n4746 ;
  assign n4749 = n4747 | n4748 ;
  assign n4750 = n4739 & n4749 ;
  assign n4751 = n4739 | n4749 ;
  assign n4752 = ~n4750 & n4751 ;
  assign n4753 = n4721 & n4752 ;
  assign n4754 = n4721 | n4752 ;
  assign n4755 = ~n4753 & n4754 ;
  assign n4756 = n4711 & n4755 ;
  assign n4757 = n4711 | n4755 ;
  assign n4758 = ~n4756 & n4757 ;
  assign n4759 = n4710 & n4758 ;
  assign n4760 = n4710 | n4758 ;
  assign n4761 = ~n4759 & n4760 ;
  assign n4762 = n4709 & n4761 ;
  assign n4763 = n4708 | n4761 ;
  assign n4764 = n336 | n4763 ;
  assign n4765 = ~n4762 & n4764 ;
  assign n4766 = n4696 | n4765 ;
  assign n4767 = n4696 & n4764 ;
  assign n4768 = ~n4762 & n4767 ;
  assign n4769 = n4766 & ~n4768 ;
  assign n4770 = n4689 | n4769 ;
  assign n4771 = n4689 & n4769 ;
  assign n4772 = n4770 & ~n4771 ;
  assign n4773 = n4690 | n4691 ;
  assign n4774 = n3777 & n4773 ;
  assign n4775 = ~n4772 & n4774 ;
  assign n4776 = n4772 & ~n4774 ;
  assign n4777 = n4775 | n4776 ;
  assign n4778 = n4762 | n4768 ;
  assign n4779 = n184 | n191 ;
  assign n4780 = n440 | n1980 ;
  assign n4781 = n859 | n2487 ;
  assign n4782 = n4780 | n4781 ;
  assign n4783 = n250 | n453 ;
  assign n4784 = n3585 | n3591 ;
  assign n4785 = n473 | n4784 ;
  assign n4786 = n3511 | n4785 ;
  assign n4787 = n4783 | n4786 ;
  assign n4788 = n337 | n4787 ;
  assign n4789 = n4782 | n4788 ;
  assign n4790 = n983 | n4789 ;
  assign n4791 = n4779 | n4790 ;
  assign n4792 = n319 | n4791 ;
  assign n4793 = n4719 | n4753 ;
  assign n4794 = n4737 & ~n4750 ;
  assign n4795 = n2680 & ~n3800 ;
  assign n4796 = n2511 & n2676 ;
  assign n4797 = n2678 & ~n3656 ;
  assign n4798 = n4796 | n4797 ;
  assign n4799 = n4795 | n4798 ;
  assign n4800 = n2684 & n3811 ;
  assign n4801 = n4799 | n4800 ;
  assign n4802 = n375 | n4801 ;
  assign n4803 = n375 & n4801 ;
  assign n4804 = n4802 & ~n4803 ;
  assign n4805 = ~n4794 & n4804 ;
  assign n4806 = n4794 & ~n4804 ;
  assign n4807 = n4805 | n4806 ;
  assign n4808 = n224 & n2538 ;
  assign n4809 = ~n906 & n4808 ;
  assign n4810 = n906 & ~n4808 ;
  assign n4811 = n4637 & ~n4810 ;
  assign n4812 = ~n4809 & n4811 ;
  assign n4813 = n4637 & ~n4812 ;
  assign n4814 = n4809 | n4812 ;
  assign n4815 = n4810 | n4814 ;
  assign n4816 = ~n4813 & n4815 ;
  assign n4817 = n224 & ~n2541 ;
  assign n4818 = ~n2544 & n4817 ;
  assign n4819 = n4734 | n4818 ;
  assign n4820 = ~n4816 & n4819 ;
  assign n4821 = n4816 & ~n4819 ;
  assign n4822 = n4820 | n4821 ;
  assign n4823 = n2526 & n2651 ;
  assign n4824 = n2618 & n2745 ;
  assign n4825 = ~n2521 & n2649 ;
  assign n4826 = n4824 | n4825 ;
  assign n4827 = n4823 | n4826 ;
  assign n4828 = n2657 & ~n3280 ;
  assign n4829 = n4827 | n4828 ;
  assign n4830 = n224 & ~n4829 ;
  assign n4831 = ~n224 & n4829 ;
  assign n4832 = n4830 | n4831 ;
  assign n4833 = ~n4822 & n4832 ;
  assign n4834 = n4822 & ~n4832 ;
  assign n4835 = n4833 | n4834 ;
  assign n4836 = n4807 | n4835 ;
  assign n4837 = n4807 & n4835 ;
  assign n4838 = n4836 & ~n4837 ;
  assign n4839 = n4793 & n4838 ;
  assign n4840 = n4793 | n4838 ;
  assign n4841 = ~n4839 & n4840 ;
  assign n4842 = n4756 | n4759 ;
  assign n4843 = n4841 & n4842 ;
  assign n4844 = n4841 | n4842 ;
  assign n4845 = ~n4843 & n4844 ;
  assign n4846 = n4792 | n4845 ;
  assign n4847 = n4792 & n4845 ;
  assign n4848 = n4846 & ~n4847 ;
  assign n4849 = n4778 & n4848 ;
  assign n4850 = n4778 | n4848 ;
  assign n4851 = ~n4849 & n4850 ;
  assign n4852 = n4771 | n4851 ;
  assign n4853 = n4771 & n4851 ;
  assign n4854 = n4852 & ~n4853 ;
  assign n4855 = n4772 | n4773 ;
  assign n4856 = n3777 & n4855 ;
  assign n4857 = ~n4854 & n4856 ;
  assign n4858 = n4854 & ~n4856 ;
  assign n4859 = n4857 | n4858 ;
  assign n4860 = n4847 | n4849 ;
  assign n4861 = n200 | n417 ;
  assign n4862 = n2189 | n4861 ;
  assign n4863 = n109 | n2188 ;
  assign n4864 = n196 | n286 ;
  assign n4865 = n124 | n238 ;
  assign n4866 = n4864 | n4865 ;
  assign n4867 = n164 | n513 ;
  assign n4868 = n382 | n393 ;
  assign n4869 = n4867 | n4868 ;
  assign n4870 = n4866 | n4869 ;
  assign n4871 = n234 | n503 ;
  assign n4872 = n247 | n251 ;
  assign n4873 = n4871 | n4872 ;
  assign n4874 = n167 | n383 ;
  assign n4875 = n205 | n305 ;
  assign n4876 = n4874 | n4875 ;
  assign n4877 = n4873 | n4876 ;
  assign n4878 = n4870 | n4877 ;
  assign n4879 = n210 | n400 ;
  assign n4880 = n389 | n4879 ;
  assign n4881 = n165 | n170 ;
  assign n4882 = n207 | n328 ;
  assign n4883 = n4881 | n4882 ;
  assign n4884 = n4880 | n4883 ;
  assign n4885 = n484 | n887 ;
  assign n4886 = n391 | n4885 ;
  assign n4887 = n325 | n399 ;
  assign n4888 = n192 | n195 ;
  assign n4889 = n4887 | n4888 ;
  assign n4890 = n4886 | n4889 ;
  assign n4891 = n4884 | n4890 ;
  assign n4892 = n4878 | n4891 ;
  assign n4893 = n4863 | n4892 ;
  assign n4894 = n4862 | n4893 ;
  assign n4895 = n117 | n280 ;
  assign n4896 = n4894 | n4895 ;
  assign n4897 = n4839 | n4843 ;
  assign n4898 = ~n4805 & n4836 ;
  assign n4899 = n4820 | n4833 ;
  assign n4900 = n224 & n2618 ;
  assign n4901 = n4814 & n4900 ;
  assign n4902 = n4814 | n4900 ;
  assign n4903 = ~n4901 & n4902 ;
  assign n4904 = n2511 & n2651 ;
  assign n4905 = ~n2521 & n2745 ;
  assign n4906 = n2526 & n2649 ;
  assign n4907 = n4905 | n4906 ;
  assign n4908 = n4904 | n4907 ;
  assign n4909 = n2635 & n2657 ;
  assign n4910 = n4908 | n4909 ;
  assign n4911 = n224 | n4910 ;
  assign n4912 = n224 & n4910 ;
  assign n4913 = n4911 & ~n4912 ;
  assign n4914 = ~n4903 & n4913 ;
  assign n4915 = n4903 & ~n4913 ;
  assign n4916 = n4914 | n4915 ;
  assign n4917 = n4899 & ~n4916 ;
  assign n4918 = ~n4899 & n4916 ;
  assign n4919 = n4917 | n4918 ;
  assign n4920 = n2684 & n3952 ;
  assign n4921 = n2676 & ~n3656 ;
  assign n4922 = n2678 & ~n3800 ;
  assign n4923 = n4921 | n4922 ;
  assign n4924 = n4920 | n4923 ;
  assign n4925 = n375 & n4924 ;
  assign n4926 = n375 | n4924 ;
  assign n4927 = ~n4925 & n4926 ;
  assign n4928 = ~n4919 & n4927 ;
  assign n4929 = n4919 & ~n4927 ;
  assign n4930 = n4928 | n4929 ;
  assign n4931 = n4898 | n4930 ;
  assign n4932 = n4898 & n4930 ;
  assign n4933 = n4931 & ~n4932 ;
  assign n4934 = n4897 & n4933 ;
  assign n4935 = n4897 | n4933 ;
  assign n4936 = ~n4934 & n4935 ;
  assign n4937 = n4896 | n4936 ;
  assign n4938 = n4896 & n4936 ;
  assign n4939 = n4937 & ~n4938 ;
  assign n4940 = n4860 & n4939 ;
  assign n4941 = n4860 | n4939 ;
  assign n4942 = ~n4940 & n4941 ;
  assign n4943 = n4853 | n4942 ;
  assign n4944 = n4853 & n4942 ;
  assign n4945 = n4943 & ~n4944 ;
  assign n4946 = n4854 | n4855 ;
  assign n4947 = n3777 & n4946 ;
  assign n4948 = ~n4945 & n4947 ;
  assign n4949 = n4945 & ~n4947 ;
  assign n4950 = n4948 | n4949 ;
  assign n4951 = n4938 | n4940 ;
  assign n4952 = n73 & n127 ;
  assign n4953 = n256 | n321 ;
  assign n4954 = n151 | n4953 ;
  assign n4955 = n200 | n4954 ;
  assign n4956 = n313 | n4955 ;
  assign n4957 = n2228 | n4956 ;
  assign n4958 = n830 | n4957 ;
  assign n4959 = n2110 | n3937 ;
  assign n4960 = n4958 | n4959 ;
  assign n4961 = n4952 | n4960 ;
  assign n4962 = n180 | n392 ;
  assign n4963 = n382 | n4962 ;
  assign n4964 = n297 | n4963 ;
  assign n4965 = n4961 | n4964 ;
  assign n4966 = n263 | n318 ;
  assign n4967 = n255 | n1985 ;
  assign n4968 = n314 | n4967 ;
  assign n4969 = n4966 | n4968 ;
  assign n4970 = n243 | n329 ;
  assign n4971 = n227 | n232 ;
  assign n4972 = n4970 | n4971 ;
  assign n4973 = n4969 | n4972 ;
  assign n4974 = n330 | n449 ;
  assign n4975 = n195 | n4974 ;
  assign n4976 = n4973 | n4975 ;
  assign n4977 = n4965 | n4976 ;
  assign n4978 = n4931 & ~n4934 ;
  assign n4979 = n4917 | n4928 ;
  assign n4980 = n4814 & ~n4900 ;
  assign n4981 = n4914 | n4980 ;
  assign n4982 = n224 & ~n2521 ;
  assign n4983 = n4900 & ~n4982 ;
  assign n4984 = ~n4900 & n4982 ;
  assign n4985 = n4981 & ~n4984 ;
  assign n4986 = ~n4983 & n4985 ;
  assign n4987 = n4981 & ~n4986 ;
  assign n4988 = n4983 | n4986 ;
  assign n4989 = n4984 | n4988 ;
  assign n4990 = ~n4987 & n4989 ;
  assign n4991 = n2651 & ~n3656 ;
  assign n4992 = n2526 & n2745 ;
  assign n4993 = n2511 & n2649 ;
  assign n4994 = n4992 | n4993 ;
  assign n4995 = n4991 | n4994 ;
  assign n4996 = n2657 & ~n3672 ;
  assign n4997 = n4995 | n4996 ;
  assign n4998 = n224 & ~n4997 ;
  assign n4999 = ~n224 & n4997 ;
  assign n5000 = n4998 | n4999 ;
  assign n5001 = n2676 & ~n3800 ;
  assign n5002 = n2684 & ~n3950 ;
  assign n5003 = n5001 | n5002 ;
  assign n5004 = n375 & ~n5003 ;
  assign n5005 = ~n375 & n5003 ;
  assign n5006 = n5004 | n5005 ;
  assign n5007 = n5000 & n5006 ;
  assign n5008 = n5000 | n5006 ;
  assign n5009 = ~n5007 & n5008 ;
  assign n5010 = ~n4990 & n5009 ;
  assign n5011 = n4990 & ~n5009 ;
  assign n5012 = n5010 | n5011 ;
  assign n5013 = n4979 & ~n5012 ;
  assign n5014 = ~n4979 & n5012 ;
  assign n5015 = n5013 | n5014 ;
  assign n5016 = n4978 | n5015 ;
  assign n5017 = n4978 & n5015 ;
  assign n5018 = n5016 & ~n5017 ;
  assign n5019 = n4977 | n5018 ;
  assign n5020 = n4977 & n5018 ;
  assign n5021 = n5019 & ~n5020 ;
  assign n5022 = n4951 & n5021 ;
  assign n5023 = n4951 | n5021 ;
  assign n5024 = ~n5022 & n5023 ;
  assign n5025 = n4944 | n5024 ;
  assign n5026 = n4944 & n5024 ;
  assign n5027 = n5025 & ~n5026 ;
  assign n5028 = n4945 | n4946 ;
  assign n5029 = n3777 & n5028 ;
  assign n5030 = ~n5027 & n5029 ;
  assign n5031 = n5027 & ~n5029 ;
  assign n5032 = n5030 | n5031 ;
  assign n5033 = n5020 | n5022 ;
  assign n5034 = n115 | n433 ;
  assign n5035 = n1332 | n2034 ;
  assign n5036 = n202 | n5035 ;
  assign n5037 = n252 | n270 ;
  assign n5038 = n990 | n2158 ;
  assign n5039 = n163 | n5038 ;
  assign n5040 = n5037 | n5039 ;
  assign n5041 = n5036 | n5040 ;
  assign n5042 = n229 | n1991 ;
  assign n5043 = n3903 | n5042 ;
  assign n5044 = n399 | n513 ;
  assign n5045 = n377 | n5044 ;
  assign n5046 = n5043 | n5045 ;
  assign n5047 = n135 | n320 ;
  assign n5048 = n177 | n5047 ;
  assign n5049 = n243 | n862 ;
  assign n5050 = n233 | n336 ;
  assign n5051 = n5049 | n5050 ;
  assign n5052 = n5048 | n5051 ;
  assign n5053 = n5046 | n5052 ;
  assign n5054 = n5041 | n5053 ;
  assign n5055 = n5034 | n5054 ;
  assign n5056 = n238 | n341 ;
  assign n5057 = n287 | n5056 ;
  assign n5058 = n5055 | n5057 ;
  assign n5059 = n400 | n5058 ;
  assign n5060 = ~n5013 & n5016 ;
  assign n5061 = n5007 | n5010 ;
  assign n5062 = n2651 & ~n3800 ;
  assign n5063 = n2511 & n2745 ;
  assign n5064 = n2649 & ~n3656 ;
  assign n5065 = n5063 | n5064 ;
  assign n5066 = n5062 | n5065 ;
  assign n5067 = n2657 & n3811 ;
  assign n5068 = n5066 | n5067 ;
  assign n5069 = n224 & ~n5068 ;
  assign n5070 = ~n224 & n5068 ;
  assign n5071 = n5069 | n5070 ;
  assign n5072 = n224 & n2526 ;
  assign n5073 = ~n375 & n4982 ;
  assign n5074 = n375 & ~n4982 ;
  assign n5075 = n5073 | n5074 ;
  assign n5076 = n5072 & ~n5075 ;
  assign n5077 = ~n5072 & n5075 ;
  assign n5078 = n5076 | n5077 ;
  assign n5079 = n5071 & ~n5078 ;
  assign n5080 = ~n5071 & n5078 ;
  assign n5081 = n5079 | n5080 ;
  assign n5082 = n4988 & ~n5081 ;
  assign n5083 = ~n4988 & n5081 ;
  assign n5084 = n5082 | n5083 ;
  assign n5085 = n5061 & ~n5084 ;
  assign n5086 = ~n5061 & n5084 ;
  assign n5087 = n5085 | n5086 ;
  assign n5088 = n5060 | n5087 ;
  assign n5089 = ~n5013 & n5087 ;
  assign n5090 = n5016 & n5089 ;
  assign n5091 = n5088 & ~n5090 ;
  assign n5092 = n5059 & n5091 ;
  assign n5093 = n5059 | n5091 ;
  assign n5094 = ~n5092 & n5093 ;
  assign n5095 = n5033 & n5094 ;
  assign n5096 = n5033 | n5094 ;
  assign n5097 = ~n5095 & n5096 ;
  assign n5098 = n5026 | n5097 ;
  assign n5099 = n5026 & n5097 ;
  assign n5100 = n5098 & ~n5099 ;
  assign n5101 = n5027 | n5028 ;
  assign n5102 = n3777 & n5101 ;
  assign n5103 = ~n5100 & n5102 ;
  assign n5104 = n5100 & ~n5102 ;
  assign n5105 = n5103 | n5104 ;
  assign n5106 = n5092 | n5095 ;
  assign n5107 = n286 | n296 ;
  assign n5108 = n117 | n5107 ;
  assign n5109 = n258 | n2041 ;
  assign n5110 = n243 | n2040 ;
  assign n5111 = n856 | n5110 ;
  assign n5112 = n5109 | n5111 ;
  assign n5113 = n158 | n1347 ;
  assign n5114 = n399 | n5113 ;
  assign n5115 = n2037 | n5114 ;
  assign n5116 = n2228 | n2304 ;
  assign n5117 = n328 | n499 ;
  assign n5118 = n170 | n5117 ;
  assign n5119 = n5116 | n5118 ;
  assign n5120 = n5115 | n5119 ;
  assign n5121 = n2321 | n3933 ;
  assign n5122 = n275 | n447 ;
  assign n5123 = n473 | n5122 ;
  assign n5124 = n5121 | n5123 ;
  assign n5125 = n5120 | n5124 ;
  assign n5126 = n2043 | n5125 ;
  assign n5127 = n122 | n2487 ;
  assign n5128 = n5126 | n5127 ;
  assign n5129 = n5112 | n5128 ;
  assign n5130 = n145 | n168 ;
  assign n5131 = n5129 | n5130 ;
  assign n5132 = n5108 | n5131 ;
  assign n5133 = n331 | n5132 ;
  assign n5134 = ~n5085 & n5088 ;
  assign n5135 = n224 & n2511 ;
  assign n5136 = n5072 | n5073 ;
  assign n5137 = ( n5073 & ~n5075 ) | ( n5073 & n5136 ) | ( ~n5075 & n5136 );
  assign n5138 = n2649 & ~n3800 ;
  assign n5139 = n2648 | n3656 ;
  assign n5140 = n2744 & ~n5139 ;
  assign n5141 = n5138 | n5140 ;
  assign n5142 = n2657 & n3952 ;
  assign n5143 = n224 & ~n5142 ;
  assign n5144 = ~n5141 & n5143 ;
  assign n5145 = n224 & ~n5144 ;
  assign n5146 = ( n5135 & n5137 ) | ( n5135 & n5144 ) | ( n5137 & n5144 );
  assign n5147 = n5141 | n5142 ;
  assign n5148 = ( n5135 & n5137 ) | ( n5135 & n5147 ) | ( n5137 & n5147 );
  assign n5149 = ( ~n5145 & n5146 ) | ( ~n5145 & n5148 ) | ( n5146 & n5148 );
  assign n5150 = ( n5135 & n5137 ) | ( n5135 & ~n5149 ) | ( n5137 & ~n5149 );
  assign n5151 = n5079 | n5082 ;
  assign n5152 = n5149 & n5151 ;
  assign n5153 = ( n5144 & ~n5145 ) | ( n5144 & n5147 ) | ( ~n5145 & n5147 );
  assign n5154 = n5151 & ~n5153 ;
  assign n5155 = ( ~n5150 & n5152 ) | ( ~n5150 & n5154 ) | ( n5152 & n5154 );
  assign n5156 = n5149 | n5151 ;
  assign n5157 = ~n5151 & n5153 ;
  assign n5158 = ( n5150 & ~n5156 ) | ( n5150 & n5157 ) | ( ~n5156 & n5157 );
  assign n5159 = n5155 | n5158 ;
  assign n5160 = n5134 | n5159 ;
  assign n5161 = n5134 & n5159 ;
  assign n5162 = n5160 & ~n5161 ;
  assign n5163 = n5133 | n5162 ;
  assign n5164 = n5133 & n5162 ;
  assign n5165 = n5163 & ~n5164 ;
  assign n5166 = n5106 & n5165 ;
  assign n5167 = n5106 | n5165 ;
  assign n5168 = ~n5166 & n5167 ;
  assign n5169 = n5099 | n5168 ;
  assign n5170 = n5099 & n5168 ;
  assign n5171 = n5169 & ~n5170 ;
  assign n5172 = n5100 | n5101 ;
  assign n5173 = n3777 & n5172 ;
  assign n5174 = ~n5171 & n5173 ;
  assign n5175 = n5171 & ~n5173 ;
  assign n5176 = n5174 | n5175 ;
  assign n5177 = n5164 | n5166 ;
  assign n5178 = n286 | n335 ;
  assign n5179 = n1014 | n5178 ;
  assign n5180 = n233 | n343 ;
  assign n5181 = n152 | n239 ;
  assign n5182 = n5180 | n5181 ;
  assign n5183 = n5179 | n5182 ;
  assign n5184 = n230 | n318 ;
  assign n5185 = n788 | n5184 ;
  assign n5186 = n168 | n251 ;
  assign n5187 = n464 | n5186 ;
  assign n5188 = n5185 | n5187 ;
  assign n5189 = n5183 | n5188 ;
  assign n5190 = n377 | n3526 ;
  assign n5191 = n2237 | n5190 ;
  assign n5192 = n389 | n814 ;
  assign n5193 = n282 | n448 ;
  assign n5194 = n1045 | n5193 ;
  assign n5195 = n196 | n5194 ;
  assign n5196 = n1043 | n5195 ;
  assign n5197 = n201 | n5196 ;
  assign n5198 = n5192 | n5197 ;
  assign n5199 = n177 | n654 ;
  assign n5200 = n135 | n4956 ;
  assign n5201 = n5199 | n5200 ;
  assign n5202 = n5198 | n5201 ;
  assign n5203 = n5191 | n5202 ;
  assign n5204 = n5189 | n5203 ;
  assign n5205 = n145 | n243 ;
  assign n5206 = n331 | n5205 ;
  assign n5207 = n5204 | n5206 ;
  assign n5208 = n459 | n5207 ;
  assign n5209 = n588 | n5208 ;
  assign n5210 = n224 & ~n3664 ;
  assign n5211 = n2657 & ~n3950 ;
  assign n5212 = n2648 | n3800 ;
  assign n5213 = n2744 & ~n5212 ;
  assign n5214 = n5211 | n5213 ;
  assign n5215 = n224 & ~n5214 ;
  assign n5216 = ~n224 & n5214 ;
  assign n5217 = n5215 | n5216 ;
  assign n5218 = ~n5210 & n5217 ;
  assign n5219 = n5210 & ~n5217 ;
  assign n5220 = n5218 | n5219 ;
  assign n5221 = ( ~n5135 & n5137 ) | ( ~n5135 & n5144 ) | ( n5137 & n5144 );
  assign n5222 = ( ~n5135 & n5137 ) | ( ~n5135 & n5147 ) | ( n5137 & n5147 );
  assign n5223 = ( ~n5145 & n5221 ) | ( ~n5145 & n5222 ) | ( n5221 & n5222 );
  assign n5224 = n5220 & ~n5223 ;
  assign n5225 = ~n5220 & n5223 ;
  assign n5226 = n5224 | n5225 ;
  assign n5227 = n5134 & ~n5155 ;
  assign n5228 = ( ~n5155 & n5159 ) | ( ~n5155 & n5227 ) | ( n5159 & n5227 );
  assign n5229 = n5226 & n5228 ;
  assign n5230 = n5226 | n5228 ;
  assign n5231 = ~n5229 & n5230 ;
  assign n5232 = n5209 & n5231 ;
  assign n5233 = n5209 | n5231 ;
  assign n5234 = ~n5232 & n5233 ;
  assign n5235 = n5177 & n5234 ;
  assign n5236 = n5177 | n5234 ;
  assign n5237 = ~n5235 & n5236 ;
  assign n5238 = n5170 | n5237 ;
  assign n5239 = n5170 & n5237 ;
  assign n5240 = n5238 & ~n5239 ;
  assign n5241 = n5171 | n5172 ;
  assign n5242 = n3777 & n5241 ;
  assign n5243 = ~n5240 & n5242 ;
  assign n5244 = n5240 & ~n5242 ;
  assign n5245 = n5243 | n5244 ;
  assign n5246 = n5240 | n5241 ;
  assign n5247 = n3777 & n5246 ;
  assign n5248 = n5232 | n5235 ;
  assign n5249 = n297 | n399 ;
  assign n5250 = n435 | n2097 ;
  assign n5251 = n207 | n249 ;
  assign n5252 = n5250 | n5251 ;
  assign n5253 = n5249 | n5252 ;
  assign n5254 = n2166 | n3532 ;
  assign n5255 = n3608 | n5048 ;
  assign n5256 = n5254 | n5255 ;
  assign n5257 = n5253 | n5256 ;
  assign n5258 = n5037 | n5257 ;
  assign n5259 = ~n2511 & n3800 ;
  assign n5260 = ( n224 & n2511 ) | ( n224 & n5259 ) | ( n2511 & n5259 );
  assign n5261 = ( ~n3800 & n5259 ) | ( ~n3800 & n5260 ) | ( n5259 & n5260 );
  assign n5262 = n224 & ~n3656 ;
  assign n5263 = ~n5135 & n5262 ;
  assign n5264 = n5210 & ~n5263 ;
  assign n5265 = ( n5217 & n5263 ) | ( n5217 & ~n5264 ) | ( n5263 & ~n5264 );
  assign n5266 = ( n5223 & ~n5261 ) | ( n5223 & n5265 ) | ( ~n5261 & n5265 );
  assign n5267 = ~n5261 & n5265 ;
  assign n5268 = ( ~n5220 & n5266 ) | ( ~n5220 & n5267 ) | ( n5266 & n5267 );
  assign n5269 = n5261 & ~n5265 ;
  assign n5270 = ( n5226 & ~n5268 ) | ( n5226 & n5269 ) | ( ~n5268 & n5269 );
  assign n5271 = ( n5228 & ~n5268 ) | ( n5228 & n5270 ) | ( ~n5268 & n5270 );
  assign n5272 = ~n5225 & n5226 ;
  assign n5273 = ( ~n5225 & n5228 ) | ( ~n5225 & n5272 ) | ( n5228 & n5272 );
  assign n5274 = ( n5265 & n5271 ) | ( n5265 & ~n5273 ) | ( n5271 & ~n5273 );
  assign n5275 = ( ~n5261 & n5271 ) | ( ~n5261 & n5274 ) | ( n5271 & n5274 );
  assign n5276 = n5258 | n5275 ;
  assign n5277 = n5258 & n5275 ;
  assign n5278 = n5276 & ~n5277 ;
  assign n5279 = n5248 & n5278 ;
  assign n5280 = n5248 | n5278 ;
  assign n5281 = ~n5279 & n5280 ;
  assign n5282 = n5239 & n5281 ;
  assign n5283 = n5239 | n5281 ;
  assign n5284 = ~n5282 & n5283 ;
  assign n5285 = n5247 & ~n5284 ;
  assign n5286 = ~n5247 & n5284 ;
  assign n5287 = n5285 | n5286 ;
  assign n5288 = n5277 | n5279 ;
  assign n5289 = n149 | n1991 ;
  assign n5290 = n812 | n5289 ;
  assign n5291 = n232 | n2444 ;
  assign n5292 = n167 | n334 ;
  assign n5293 = n5291 | n5292 ;
  assign n5294 = n255 | n275 ;
  assign n5295 = n121 | n251 ;
  assign n5296 = n5294 | n5295 ;
  assign n5297 = n5293 | n5296 ;
  assign n5298 = n5290 | n5297 ;
  assign n5299 = n524 | n1980 ;
  assign n5300 = n208 | n862 ;
  assign n5301 = n200 | n5300 ;
  assign n5302 = n5299 | n5301 ;
  assign n5303 = n5298 | n5302 ;
  assign n5304 = n466 | n5303 ;
  assign n5305 = n392 | n5304 ;
  assign n5306 = n5288 & n5305 ;
  assign n5307 = n5277 | n5305 ;
  assign n5308 = n5279 | n5307 ;
  assign n5309 = ~n5306 & n5308 ;
  assign n5310 = ~n5282 & n5309 ;
  assign n5311 = n5282 & ~n5309 ;
  assign n5312 = n5310 | n5311 ;
  assign n5313 = n5246 | n5284 ;
  assign n5314 = n3777 & n5313 ;
  assign n5315 = ~n5312 & n5314 ;
  assign n5316 = n5312 & ~n5314 ;
  assign n5317 = n5315 | n5316 ;
  assign n5318 = n5312 | n5313 ;
  assign n5319 = n3777 & n5318 ;
  assign n5320 = n5282 & n5309 ;
  assign n5321 = n200 | n330 ;
  assign n5322 = n503 | n5321 ;
  assign n5323 = n1059 | n2027 ;
  assign n5324 = n424 | n479 ;
  assign n5325 = n1037 | n5324 ;
  assign n5326 = n5323 | n5325 ;
  assign n5327 = n179 | n5326 ;
  assign n5328 = n168 | n3569 ;
  assign n5329 = n5327 | n5328 ;
  assign n5330 = n870 | n5329 ;
  assign n5331 = n5322 | n5330 ;
  assign n5332 = n5306 | n5331 ;
  assign n5333 = n5320 & n5332 ;
  assign n5334 = n5320 | n5332 ;
  assign n5335 = n5305 & n5331 ;
  assign n5336 = n5288 & n5335 ;
  assign n5337 = n5334 & ~n5336 ;
  assign n5338 = ~n5333 & n5337 ;
  assign n5339 = n5319 & ~n5338 ;
  assign n5340 = ~n5319 & n5338 ;
  assign n5341 = n5339 | n5340 ;
  assign n5342 = n316 | n328 ;
  assign n5343 = n393 | n4289 ;
  assign n5344 = n5196 | n5343 ;
  assign n5345 = n5342 | n5344 ;
  assign n5346 = n798 | n2410 ;
  assign n5347 = n148 | n3577 ;
  assign n5348 = n207 | n5347 ;
  assign n5349 = n5346 | n5348 ;
  assign n5350 = n5345 | n5349 ;
  assign n5351 = n163 | n5350 ;
  assign n5352 = n5336 | n5351 ;
  assign n5353 = n5336 & n5351 ;
  assign n5354 = n5352 & ~n5353 ;
  assign n5355 = n5333 | n5354 ;
  assign n5356 = n5333 & n5354 ;
  assign n5357 = n5355 & ~n5356 ;
  assign n5358 = n5318 | n5338 ;
  assign n5359 = n3777 & n5358 ;
  assign n5360 = ~n5357 & n5359 ;
  assign n5361 = n5357 & ~n5359 ;
  assign n5362 = n5360 | n5361 ;
  assign n5363 = n5357 | n5358 ;
  assign n5364 = n3777 & n5363 ;
  assign n5365 = n124 | n4613 ;
  assign n5366 = n157 | n3539 ;
  assign n5367 = n179 | n5366 ;
  assign n5368 = n5365 | n5367 ;
  assign n5369 = n153 | n184 ;
  assign n5370 = n177 | n291 ;
  assign n5371 = n377 | n5370 ;
  assign n5372 = n227 | n246 ;
  assign n5373 = n168 | n274 ;
  assign n5374 = n5372 | n5373 ;
  assign n5375 = n5371 | n5374 ;
  assign n5376 = n186 | n1981 ;
  assign n5377 = n877 | n5376 ;
  assign n5378 = n5375 | n5377 ;
  assign n5379 = n871 | n875 ;
  assign n5380 = n327 | n790 ;
  assign n5381 = n290 | n5380 ;
  assign n5382 = n865 | n5381 ;
  assign n5383 = n5379 | n5382 ;
  assign n5384 = n5378 | n5383 ;
  assign n5385 = n5369 | n5384 ;
  assign n5386 = n5368 | n5385 ;
  assign n5387 = n389 | n5386 ;
  assign n5388 = n5353 & n5387 ;
  assign n5389 = n5353 | n5387 ;
  assign n5390 = ~n5388 & n5389 ;
  assign n5391 = n5356 | n5390 ;
  assign n5392 = n5331 & n5389 ;
  assign n5393 = n5354 & n5392 ;
  assign n5394 = n5320 & n5393 ;
  assign n5395 = n5391 & ~n5394 ;
  assign n5396 = n5364 & ~n5395 ;
  assign n5397 = ~n5364 & n5395 ;
  assign n5398 = n5396 | n5397 ;
  assign n5399 = n5363 | n5395 ;
  assign n5400 = n3777 & n5399 ;
  assign n5401 = n171 | n448 ;
  assign n5402 = n229 | n5401 ;
  assign n5403 = n167 | n1029 ;
  assign n5404 = n318 | n5403 ;
  assign n5405 = n316 | n5404 ;
  assign n5406 = n5402 | n5405 ;
  assign n5407 = n323 | n655 ;
  assign n5408 = n294 | n852 ;
  assign n5409 = n163 | n5408 ;
  assign n5410 = n262 | n5409 ;
  assign n5411 = n5407 | n5410 ;
  assign n5412 = n135 | n230 ;
  assign n5413 = n134 | n153 ;
  assign n5414 = n238 | n313 ;
  assign n5415 = n166 | n5414 ;
  assign n5416 = n216 | n5415 ;
  assign n5417 = n5413 | n5416 ;
  assign n5418 = n148 | n233 ;
  assign n5419 = n145 | n433 ;
  assign n5420 = n137 | n264 ;
  assign n5421 = n5419 | n5420 ;
  assign n5422 = n5418 | n5421 ;
  assign n5423 = n5417 | n5422 ;
  assign n5424 = n5412 | n5423 ;
  assign n5425 = n5411 | n5424 ;
  assign n5426 = n263 | n317 ;
  assign n5427 = n142 | n158 ;
  assign n5428 = n177 | n5427 ;
  assign n5429 = n5426 | n5428 ;
  assign n5430 = n312 | n5429 ;
  assign n5431 = n5425 | n5430 ;
  assign n5432 = n5406 | n5431 ;
  assign n5433 = n405 | n5432 ;
  assign n5434 = n2123 | n5433 ;
  assign n5435 = n5388 | n5434 ;
  assign n5436 = n5388 & n5434 ;
  assign n5437 = n5435 & ~n5436 ;
  assign n5438 = n5394 & n5437 ;
  assign n5439 = n5394 | n5437 ;
  assign n5440 = ~n5438 & n5439 ;
  assign n5441 = n5400 & n5440 ;
  assign n5442 = n5400 | n5440 ;
  assign n5443 = ~n5441 & n5442 ;
  assign n5444 = n5399 | n5440 ;
  assign n5445 = n3777 & n5444 ;
  assign n5446 = n5394 | n5436 ;
  assign n5447 = n5435 & n5446 ;
  assign n5448 = n148 | n345 ;
  assign n5449 = n138 | n306 ;
  assign n5450 = n5401 | n5449 ;
  assign n5451 = n5448 | n5450 ;
  assign n5452 = n157 | n189 ;
  assign n5453 = n176 | n215 ;
  assign n5454 = n140 | n249 ;
  assign n5455 = n5453 | n5454 ;
  assign n5456 = n153 | n5455 ;
  assign n5457 = n340 | n5419 ;
  assign n5458 = n5403 | n5457 ;
  assign n5459 = n5456 | n5458 ;
  assign n5460 = n134 | n303 ;
  assign n5461 = n163 | n405 ;
  assign n5462 = n258 | n5461 ;
  assign n5463 = n166 | n5462 ;
  assign n5464 = n5460 | n5463 ;
  assign n5465 = n5459 | n5464 ;
  assign n5466 = n5452 | n5465 ;
  assign n5467 = n5451 | n5466 ;
  assign n5468 = n5428 | n5467 ;
  assign n5469 = n5447 & n5468 ;
  assign n5470 = n5447 | n5468 ;
  assign n5471 = ~n5469 & n5470 ;
  assign n5472 = n5445 & n5471 ;
  assign n5473 = n5445 | n5471 ;
  assign n5474 = ~n5472 & n5473 ;
  assign n5475 = ~n5445 & n5469 ;
  assign n5476 = pi21 | n65 ;
  assign n5477 = pi22 | n5476 ;
  assign n5478 = ~n5475 & n5477 ;
  assign n5479 = n4599 | n5468 ;
  assign n5480 = n4598 | n5479 ;
  assign n5481 = n4690 | n5480 ;
  assign n5482 = n4772 | n5481 ;
  assign n5483 = n4854 | n5482 ;
  assign n5484 = n4945 | n5483 ;
  assign n5485 = n5027 | n5484 ;
  assign n5486 = n5100 | n5485 ;
  assign n5487 = n5171 | n5486 ;
  assign n5488 = n5240 | n5487 ;
  assign n5489 = n5284 | n5488 ;
  assign n5490 = n5312 | n5489 ;
  assign n5491 = n5357 | n5490 ;
  assign n5492 = n5440 | n5491 ;
  assign n5493 = n5338 | n5395 ;
  assign n5494 = n5447 | n5493 ;
  assign n5495 = n5492 | n5494 ;
  assign n5496 = n3777 & n5495 ;
  assign n5497 = ~n5469 & n5496 ;
  assign n5498 = n5478 & ~n5497 ;
  assign n5499 = n5477 & ~n5495 ;
  assign n5500 = n3777 & ~n5499 ;
  assign po0 = n3774 ;
  assign po1 = n3926 ;
  assign po2 = n4045 ;
  assign po3 = n4161 ;
  assign po4 = n4281 ;
  assign po5 = n4390 ;
  assign po6 = n4496 ;
  assign po7 = n4603 ;
  assign po8 = n4695 ;
  assign po9 = n4777 ;
  assign po10 = n4859 ;
  assign po11 = n4950 ;
  assign po12 = n5032 ;
  assign po13 = n5105 ;
  assign po14 = n5176 ;
  assign po15 = n5245 ;
  assign po16 = n5287 ;
  assign po17 = n5317 ;
  assign po18 = n5341 ;
  assign po19 = n5362 ;
  assign po20 = n5398 ;
  assign po21 = n5443 ;
  assign po22 = n5474 ;
  assign po23 = ~n5498 ;
  assign po24 = n5500 ;
endmodule
