module top(G7 , G121 , G119 , G147 , G53 , G86 , G43 , G96 , G32 , G76 , G64 , G106 , G146 , G145 , G89 , G99 , G79 , G109 , G115 , G124 , G137 , G139 , G140 , G141 , G142 , G11 , G2 , G74 , G88 , G98 , G78 , G108 , G90 , G100 , G80 , G110 , G120 , G117 , G57 , G46 , G36 , G68 , G58 , G47 , G37 , G69 , G59 , G48 , G38 , G70 , G122 , G52 , G42 , G31 , G63 , G28 , G116 , G1 , G3 , G60 , G49 , G39 , G71 , G56 , G35 , G67 , G55 , G45 , G34 , G66 , G54 , G44 , G33 , G65 , G61 , G50 , G40 , G72 , G123 , G118 , G144 , G143 , G87 , G97 , G77 , G107 , G155 , G154 , G125 , G126 , G153 , G152 , G151 , G150 , G149 , G148 , G10 , G157 , G138 , G133 , G134 , G135 , G136 , G131 , G132 , G129 , G130 , G156 , G128 , G9 , G22 , G23 , G27 , G24 , G93 , G103 , G83 , G113 , G20 , G92 , G102 , G82 , G112 , G25 , G91 , G101 , G81 , G111 , G21 , G26 , G16 , G12 , G17 , G6 , G18 , G19 , G85 , G95 , G75 , G105 , G13 , G4 , G14 , G5 , G15 , G62 , G51 , G41 , G73 , G94 , G104 , G84 , G114 , G29 , G30 , G127 , G8 , G2551 , G2552 , G2553 , G2554 , G2555 , G2556 , G2557 , G2531 , G2532 , G2533 , G2534 , G2535 , G2536 , G2537 , G2538 , G2539 , G2540 , G2541 , G2542 , G2543 , G2544 , G2545 , G2546 , G2547 , G2548 , G2549 , G2550 , G2558 , G2559 , G2560 , G2561 , G2562 , G2563 , G2564 , G2565 , G2566 , G2567 , G2568 , G2569 , G2570 , G2571 , G2572 , G2573 , G2574 , G2575 , G2576 , G2577 , G2578 , G2579 , G2580 , G2581 , G2582 , G2583 , G2584 , G2585 , G2586 , G2587 , G2588 , G2589 , G2590 , G2591 , G2592 , G2593 , G2594 );
  input G7 , G121 , G119 , G147 , G53 , G86 , G43 , G96 , G32 , G76 , G64 , G106 , G146 , G145 , G89 , G99 , G79 , G109 , G115 , G124 , G137 , G139 , G140 , G141 , G142 , G11 , G2 , G74 , G88 , G98 , G78 , G108 , G90 , G100 , G80 , G110 , G120 , G117 , G57 , G46 , G36 , G68 , G58 , G47 , G37 , G69 , G59 , G48 , G38 , G70 , G122 , G52 , G42 , G31 , G63 , G28 , G116 , G1 , G3 , G60 , G49 , G39 , G71 , G56 , G35 , G67 , G55 , G45 , G34 , G66 , G54 , G44 , G33 , G65 , G61 , G50 , G40 , G72 , G123 , G118 , G144 , G143 , G87 , G97 , G77 , G107 , G155 , G154 , G125 , G126 , G153 , G152 , G151 , G150 , G149 , G148 , G10 , G157 , G138 , G133 , G134 , G135 , G136 , G131 , G132 , G129 , G130 , G156 , G128 , G9 , G22 , G23 , G27 , G24 , G93 , G103 , G83 , G113 , G20 , G92 , G102 , G82 , G112 , G25 , G91 , G101 , G81 , G111 , G21 , G26 , G16 , G12 , G17 , G6 , G18 , G19 , G85 , G95 , G75 , G105 , G13 , G4 , G14 , G5 , G15 , G62 , G51 , G41 , G73 , G94 , G104 , G84 , G114 , G29 , G30 , G127 , G8 ;
  output G2551 , G2552 , G2553 , G2554 , G2555 , G2556 , G2557 , G2531 , G2532 , G2533 , G2534 , G2535 , G2536 , G2537 , G2538 , G2539 , G2540 , G2541 , G2542 , G2543 , G2544 , G2545 , G2546 , G2547 , G2548 , G2549 , G2550 , G2558 , G2559 , G2560 , G2561 , G2562 , G2563 , G2564 , G2565 , G2566 , G2567 , G2568 , G2569 , G2570 , G2571 , G2572 , G2573 , G2574 , G2575 , G2576 , G2577 , G2578 , G2579 , G2580 , G2581 , G2582 , G2583 , G2584 , G2585 , G2586 , G2587 , G2588 , G2589 , G2590 , G2591 , G2592 , G2593 , G2594 ;
  wire n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650;
  assign n158 = G7 & G121 ;
  assign n159 = G119 & n158 ;
  assign n160 = G147 & n158 ;
  assign n161 = G53 & G86 ;
  assign n162 = G43 & G96 ;
  assign n163 = n161 & n162 ;
  assign n164 = G32 & G76 ;
  assign n165 = G64 & G106 ;
  assign n166 = n164 & n165 ;
  assign n167 = n163 & n166 ;
  assign n168 = G147 & ~n166 ;
  assign n169 = G119 & ~n163 ;
  assign n170 = n168 | n169 ;
  assign n171 = ( G146 & G145 ) | ( G146 & ~G99 ) | ( G145 & ~G99 );
  assign n172 = ( ~G146 & G145 ) | ( ~G146 & G89 ) | ( G145 & G89 );
  assign n173 = ~n171 & n172 ;
  assign n174 = ( G146 & ~G145 ) | ( G146 & G109 ) | ( ~G145 & G109 );
  assign n175 = ( G146 & G145 ) | ( G146 & G79 ) | ( G145 & G79 );
  assign n176 = n174 & n175 ;
  assign n177 = n173 | n176 ;
  assign n178 = G139 & G140 ;
  assign n179 = G141 & G142 ;
  assign n180 = n178 & n179 ;
  assign n181 = G11 & G2 ;
  assign n182 = G121 & n181 ;
  assign n183 = ~G115 & G74 ;
  assign n184 = ( G146 & G145 ) | ( G146 & ~G98 ) | ( G145 & ~G98 );
  assign n185 = ( ~G146 & G145 ) | ( ~G146 & G88 ) | ( G145 & G88 );
  assign n186 = ~n184 & n185 ;
  assign n187 = ( G146 & ~G145 ) | ( G146 & G108 ) | ( ~G145 & G108 );
  assign n188 = ( G146 & G145 ) | ( G146 & G78 ) | ( G145 & G78 );
  assign n189 = n187 & n188 ;
  assign n190 = n186 | n189 ;
  assign n191 = ( G146 & G145 ) | ( G146 & ~G100 ) | ( G145 & ~G100 );
  assign n192 = ( ~G146 & G145 ) | ( ~G146 & G90 ) | ( G145 & G90 );
  assign n193 = ~n191 & n192 ;
  assign n194 = ( G146 & ~G145 ) | ( G146 & G110 ) | ( ~G145 & G110 );
  assign n195 = ( G146 & G145 ) | ( G146 & G80 ) | ( G145 & G80 );
  assign n196 = n194 & n195 ;
  assign n197 = n193 | n196 ;
  assign n198 = ( G120 & G117 ) | ( G120 & ~G46 ) | ( G117 & ~G46 );
  assign n199 = ( ~G120 & G117 ) | ( ~G120 & G57 ) | ( G117 & G57 );
  assign n200 = ~n198 & n199 ;
  assign n201 = ( G120 & ~G117 ) | ( G120 & G68 ) | ( ~G117 & G68 );
  assign n202 = ( G120 & G117 ) | ( G120 & G36 ) | ( G117 & G36 );
  assign n203 = n201 & n202 ;
  assign n204 = n200 | n203 ;
  assign n205 = ( G120 & G117 ) | ( G120 & ~G47 ) | ( G117 & ~G47 );
  assign n206 = ( ~G120 & G117 ) | ( ~G120 & G58 ) | ( G117 & G58 );
  assign n207 = ~n205 & n206 ;
  assign n208 = ( G120 & ~G117 ) | ( G120 & G69 ) | ( ~G117 & G69 );
  assign n209 = ( G120 & G117 ) | ( G120 & G37 ) | ( G117 & G37 );
  assign n210 = n208 & n209 ;
  assign n211 = n207 | n210 ;
  assign n212 = ( G120 & G117 ) | ( G120 & ~G48 ) | ( G117 & ~G48 );
  assign n213 = ( ~G120 & G117 ) | ( ~G120 & G59 ) | ( G117 & G59 );
  assign n214 = ~n212 & n213 ;
  assign n215 = ( G120 & ~G117 ) | ( G120 & G70 ) | ( ~G117 & G70 );
  assign n216 = ( G120 & G117 ) | ( G120 & G38 ) | ( G117 & G38 );
  assign n217 = n215 & n216 ;
  assign n218 = n214 | n217 ;
  assign n219 = ( G120 & G117 ) | ( G120 & ~G42 ) | ( G117 & ~G42 );
  assign n220 = ( ~G120 & G117 ) | ( ~G120 & G52 ) | ( G117 & G52 );
  assign n221 = ~n219 & n220 ;
  assign n222 = ( G120 & ~G117 ) | ( G120 & G63 ) | ( ~G117 & G63 );
  assign n223 = ( G120 & G117 ) | ( G120 & G31 ) | ( G117 & G31 );
  assign n224 = n222 & n223 ;
  assign n225 = n221 | n224 ;
  assign n226 = G122 & n225 ;
  assign n227 = G122 & ~n226 ;
  assign n228 = ~G121 & G116 ;
  assign n229 = G28 & ~n170 ;
  assign n230 = n228 & n229 ;
  assign n231 = G1 & G3 ;
  assign n232 = n170 | n231 ;
  assign n233 = n228 & ~n232 ;
  assign n234 = ( G120 & G117 ) | ( G120 & ~G49 ) | ( G117 & ~G49 );
  assign n235 = ( ~G120 & G117 ) | ( ~G120 & G60 ) | ( G117 & G60 );
  assign n236 = ~n234 & n235 ;
  assign n237 = ( G120 & ~G117 ) | ( G120 & G71 ) | ( ~G117 & G71 );
  assign n238 = ( G120 & G117 ) | ( G120 & G39 ) | ( G117 & G39 );
  assign n239 = n237 & n238 ;
  assign n240 = n236 | n239 ;
  assign n241 = G117 | G56 ;
  assign n242 = ~G120 & n241 ;
  assign n243 = ( G120 & ~G117 ) | ( G120 & G67 ) | ( ~G117 & G67 );
  assign n244 = ( G120 & G117 ) | ( G120 & G35 ) | ( G117 & G35 );
  assign n245 = n243 & n244 ;
  assign n246 = n242 | n245 ;
  assign n247 = ( G120 & G117 ) | ( G120 & ~G45 ) | ( G117 & ~G45 );
  assign n248 = ( ~G120 & G117 ) | ( ~G120 & G55 ) | ( G117 & G55 );
  assign n249 = ~n247 & n248 ;
  assign n250 = ( G120 & ~G117 ) | ( G120 & G66 ) | ( ~G117 & G66 );
  assign n251 = ( G120 & G117 ) | ( G120 & G34 ) | ( G117 & G34 );
  assign n252 = n250 & n251 ;
  assign n253 = n249 | n252 ;
  assign n254 = ( G120 & G117 ) | ( G120 & ~G44 ) | ( G117 & ~G44 );
  assign n255 = ( ~G120 & G117 ) | ( ~G120 & G54 ) | ( G117 & G54 );
  assign n256 = ~n254 & n255 ;
  assign n257 = ( G120 & ~G117 ) | ( G120 & G65 ) | ( ~G117 & G65 );
  assign n258 = ( G120 & G117 ) | ( G120 & G33 ) | ( G117 & G33 );
  assign n259 = n257 & n258 ;
  assign n260 = n256 | n259 ;
  assign n261 = G123 & ~n218 ;
  assign n262 = ( G120 & G117 ) | ( G120 & ~G50 ) | ( G117 & ~G50 );
  assign n263 = ( ~G120 & G117 ) | ( ~G120 & G61 ) | ( G117 & G61 );
  assign n264 = ~n262 & n263 ;
  assign n265 = ( G120 & ~G117 ) | ( G120 & G72 ) | ( ~G117 & G72 );
  assign n266 = ( G120 & G117 ) | ( G120 & G40 ) | ( G117 & G40 );
  assign n267 = n265 & n266 ;
  assign n268 = n264 | n267 ;
  assign n269 = ~G123 & n268 ;
  assign n270 = n261 | n269 ;
  assign n271 = G123 | n240 ;
  assign n272 = G123 & n211 ;
  assign n273 = n271 & ~n272 ;
  assign n274 = ~G122 & G118 ;
  assign n275 = n268 | n274 ;
  assign n276 = G118 | n268 ;
  assign n277 = G123 & n276 ;
  assign n278 = ~G123 & n225 ;
  assign n279 = n277 | n278 ;
  assign n280 = ( G146 & G145 ) | ( G146 & ~G97 ) | ( G145 & ~G97 );
  assign n281 = ( ~G146 & G145 ) | ( ~G146 & G87 ) | ( G145 & G87 );
  assign n282 = ~n280 & n281 ;
  assign n283 = ( G146 & ~G145 ) | ( G146 & G107 ) | ( ~G145 & G107 );
  assign n284 = ( G146 & G145 ) | ( G146 & G77 ) | ( G145 & G77 );
  assign n285 = n283 & n284 ;
  assign n286 = n282 | n285 ;
  assign n287 = G143 & ~n286 ;
  assign n288 = ( G144 & G143 ) | ( G144 & ~n287 ) | ( G143 & ~n287 );
  assign n289 = ( n286 & n287 ) | ( n286 & ~n288 ) | ( n287 & ~n288 );
  assign n290 = G149 & ~G148 ;
  assign n291 = ~G149 & G148 ;
  assign n292 = n290 | n291 ;
  assign n293 = G153 & ~G152 ;
  assign n294 = ~G153 & G152 ;
  assign n295 = n293 | n294 ;
  assign n296 = G151 & ~G150 ;
  assign n297 = ~G151 & G150 ;
  assign n298 = n296 | n297 ;
  assign n299 = ( n292 & n295 ) | ( n292 & ~n298 ) | ( n295 & ~n298 );
  assign n300 = ( ~n295 & n298 ) | ( ~n295 & n299 ) | ( n298 & n299 );
  assign n301 = ( ~n292 & n299 ) | ( ~n292 & n300 ) | ( n299 & n300 );
  assign n302 = ~G125 & G126 ;
  assign n303 = G125 & ~G126 ;
  assign n304 = n302 | n303 ;
  assign n305 = ( ~G155 & G154 ) | ( ~G155 & n304 ) | ( G154 & n304 );
  assign n306 = ( G155 & ~G154 ) | ( G155 & n305 ) | ( ~G154 & n305 );
  assign n307 = ( ~n304 & n305 ) | ( ~n304 & n306 ) | ( n305 & n306 );
  assign n308 = ~n299 & n307 ;
  assign n309 = n292 & n307 ;
  assign n310 = ( ~n300 & n308 ) | ( ~n300 & n309 ) | ( n308 & n309 );
  assign n311 = ( G10 & ~n307 ) | ( G10 & n310 ) | ( ~n307 & n310 );
  assign n312 = ( n301 & n310 ) | ( n301 & n311 ) | ( n310 & n311 );
  assign n313 = G157 & G138 ;
  assign n314 = G157 | G138 ;
  assign n315 = ~n313 & n314 ;
  assign n316 = ~G141 & G142 ;
  assign n317 = G141 & ~G142 ;
  assign n318 = n316 | n317 ;
  assign n319 = ~G139 & G140 ;
  assign n320 = G139 & ~G140 ;
  assign n321 = n319 | n320 ;
  assign n322 = ( n315 & n318 ) | ( n315 & ~n321 ) | ( n318 & ~n321 );
  assign n323 = ( ~n318 & n321 ) | ( ~n318 & n322 ) | ( n321 & n322 );
  assign n324 = ( ~n315 & n322 ) | ( ~n315 & n323 ) | ( n322 & n323 );
  assign n325 = ( ~G144 & G143 ) | ( ~G144 & n324 ) | ( G143 & n324 );
  assign n326 = ( G144 & ~G143 ) | ( G144 & n325 ) | ( ~G143 & n325 );
  assign n327 = ( ~n324 & n325 ) | ( ~n324 & n326 ) | ( n325 & n326 );
  assign n328 = ~G135 & G136 ;
  assign n329 = G135 & ~G136 ;
  assign n330 = n328 | n329 ;
  assign n331 = ( G133 & ~G134 ) | ( G133 & n330 ) | ( ~G134 & n330 );
  assign n332 = ( ~G133 & G134 ) | ( ~G133 & n331 ) | ( G134 & n331 );
  assign n333 = ( ~n330 & n331 ) | ( ~n330 & n332 ) | ( n331 & n332 );
  assign n334 = G156 & G128 ;
  assign n335 = G156 | G128 ;
  assign n336 = ~n334 & n335 ;
  assign n337 = ~G131 & G132 ;
  assign n338 = G131 & ~G132 ;
  assign n339 = n337 | n338 ;
  assign n340 = ~G129 & G130 ;
  assign n341 = G129 & ~G130 ;
  assign n342 = n340 | n341 ;
  assign n343 = ( n336 & n339 ) | ( n336 & ~n342 ) | ( n339 & ~n342 );
  assign n344 = ( ~n339 & n342 ) | ( ~n339 & n343 ) | ( n342 & n343 );
  assign n345 = ( ~n336 & n343 ) | ( ~n336 & n344 ) | ( n343 & n344 );
  assign n346 = n333 & ~n345 ;
  assign n347 = ~n333 & n345 ;
  assign n348 = n346 | n347 ;
  assign n349 = G12 & G6 ;
  assign n350 = ~G12 & n253 ;
  assign n351 = n349 | n350 ;
  assign n352 = G12 & G18 ;
  assign n353 = ~G12 & n260 ;
  assign n354 = n352 | n353 ;
  assign n355 = G23 & G19 ;
  assign n356 = ( G146 & G145 ) | ( G146 & ~G95 ) | ( G145 & ~G95 );
  assign n357 = ( ~G146 & G145 ) | ( ~G146 & G85 ) | ( G145 & G85 );
  assign n358 = ~n356 & n357 ;
  assign n359 = ( G146 & ~G145 ) | ( G146 & G105 ) | ( ~G145 & G105 );
  assign n360 = ( G146 & G145 ) | ( G146 & G75 ) | ( G145 & G75 );
  assign n361 = n359 & n360 ;
  assign n362 = n358 | n361 ;
  assign n363 = ~G23 & n362 ;
  assign n364 = n355 | n363 ;
  assign n365 = G135 & ~n364 ;
  assign n366 = ( G134 & ~n354 ) | ( G134 & n365 ) | ( ~n354 & n365 );
  assign n367 = ~G135 & n364 ;
  assign n368 = ( ~G134 & n354 ) | ( ~G134 & n367 ) | ( n354 & n367 );
  assign n369 = n366 | n368 ;
  assign n370 = ( ~G133 & n351 ) | ( ~G133 & n369 ) | ( n351 & n369 );
  assign n371 = G16 & G12 ;
  assign n372 = ~G12 & n204 ;
  assign n373 = n371 | n372 ;
  assign n374 = G12 & G17 ;
  assign n375 = ~G12 & n246 ;
  assign n376 = n374 | n375 ;
  assign n377 = G132 & ~n376 ;
  assign n378 = ( G131 & ~n373 ) | ( G131 & n377 ) | ( ~n373 & n377 );
  assign n379 = ~G132 & n376 ;
  assign n380 = ( ~G131 & n373 ) | ( ~G131 & n379 ) | ( n373 & n379 );
  assign n381 = n378 | n380 ;
  assign n382 = ( G133 & ~n351 ) | ( G133 & n381 ) | ( ~n351 & n381 );
  assign n383 = n370 | n382 ;
  assign n384 = G12 & G14 ;
  assign n385 = ~G12 & n240 ;
  assign n386 = n384 | n385 ;
  assign n387 = G12 & G5 ;
  assign n388 = ~G12 & n218 ;
  assign n389 = n387 | n388 ;
  assign n390 = G12 & G15 ;
  assign n391 = ~G12 & n211 ;
  assign n392 = n390 | n391 ;
  assign n393 = G130 & ~n392 ;
  assign n394 = ( G129 & ~n389 ) | ( G129 & n393 ) | ( ~n389 & n393 );
  assign n395 = ~G130 & n392 ;
  assign n396 = ( ~G129 & n389 ) | ( ~G129 & n395 ) | ( n389 & n395 );
  assign n397 = n394 | n396 ;
  assign n398 = ( ~G128 & n386 ) | ( ~G128 & n397 ) | ( n386 & n397 );
  assign n399 = G12 & G13 ;
  assign n400 = ~G12 & n225 ;
  assign n401 = n399 | n400 ;
  assign n402 = G12 & G4 ;
  assign n403 = ~G12 & n268 ;
  assign n404 = n402 | n403 ;
  assign n405 = G126 & ~n404 ;
  assign n406 = ( G125 & ~n401 ) | ( G125 & n405 ) | ( ~n401 & n405 );
  assign n407 = ~G126 & n404 ;
  assign n408 = ( ~G125 & n401 ) | ( ~G125 & n407 ) | ( n401 & n407 );
  assign n409 = n406 | n408 ;
  assign n410 = ( G128 & ~n386 ) | ( G128 & n409 ) | ( ~n386 & n409 );
  assign n411 = n398 | n410 ;
  assign n412 = n383 | n411 ;
  assign n413 = G23 & G27 ;
  assign n414 = ~G23 & n190 ;
  assign n415 = n413 | n414 ;
  assign n416 = G22 & G23 ;
  assign n417 = ~G23 & n286 ;
  assign n418 = n416 | n417 ;
  assign n419 = ( ~G142 & n415 ) | ( ~G142 & n418 ) | ( n415 & n418 );
  assign n420 = G23 & G24 ;
  assign n421 = ( G146 & G145 ) | ( G146 & ~G103 ) | ( G145 & ~G103 );
  assign n422 = ( ~G146 & G145 ) | ( ~G146 & G93 ) | ( G145 & G93 );
  assign n423 = ~n421 & n422 ;
  assign n424 = ( G146 & ~G145 ) | ( G146 & G113 ) | ( ~G145 & G113 );
  assign n425 = ( G146 & G145 ) | ( G146 & G83 ) | ( G145 & G83 );
  assign n426 = n424 & n425 ;
  assign n427 = n423 | n426 ;
  assign n428 = ~G23 & n427 ;
  assign n429 = n420 | n428 ;
  assign n430 = G136 & ~n429 ;
  assign n431 = G23 & G20 ;
  assign n432 = ( G146 & G145 ) | ( G146 & ~G102 ) | ( G145 & ~G102 );
  assign n433 = ( ~G146 & G145 ) | ( ~G146 & G92 ) | ( G145 & G92 );
  assign n434 = ~n432 & n433 ;
  assign n435 = ( G146 & ~G145 ) | ( G146 & G112 ) | ( ~G145 & G112 );
  assign n436 = ( G146 & G145 ) | ( G146 & G82 ) | ( G145 & G82 );
  assign n437 = n435 & n436 ;
  assign n438 = n434 | n437 ;
  assign n439 = ~G23 & n438 ;
  assign n440 = n431 | n439 ;
  assign n441 = ( G138 & n430 ) | ( G138 & ~n440 ) | ( n430 & ~n440 );
  assign n442 = ~G136 & n429 ;
  assign n443 = ( ~G138 & n440 ) | ( ~G138 & n442 ) | ( n440 & n442 );
  assign n444 = n441 | n443 ;
  assign n445 = G23 & G25 ;
  assign n446 = ( G146 & G145 ) | ( G146 & ~G101 ) | ( G145 & ~G101 );
  assign n447 = ( ~G146 & G145 ) | ( ~G146 & G91 ) | ( G145 & G91 );
  assign n448 = ~n446 & n447 ;
  assign n449 = ( G146 & ~G145 ) | ( G146 & G111 ) | ( ~G145 & G111 );
  assign n450 = ( G146 & G145 ) | ( G146 & G81 ) | ( G145 & G81 );
  assign n451 = n449 & n450 ;
  assign n452 = n448 | n451 ;
  assign n453 = ~G23 & n452 ;
  assign n454 = n445 | n453 ;
  assign n455 = ( G139 & n444 ) | ( G139 & ~n454 ) | ( n444 & ~n454 );
  assign n456 = G23 & G21 ;
  assign n457 = ~G23 & n197 ;
  assign n458 = n456 | n457 ;
  assign n459 = G23 & G26 ;
  assign n460 = ~G23 & n177 ;
  assign n461 = n459 | n460 ;
  assign n462 = G141 & ~n461 ;
  assign n463 = ( G140 & ~n458 ) | ( G140 & n462 ) | ( ~n458 & n462 );
  assign n464 = ~G141 & n461 ;
  assign n465 = ( ~G140 & n458 ) | ( ~G140 & n464 ) | ( n458 & n464 );
  assign n466 = n463 | n465 ;
  assign n467 = ( ~G139 & n454 ) | ( ~G139 & n466 ) | ( n454 & n466 );
  assign n468 = n455 | n467 ;
  assign n469 = ( ~G142 & n415 ) | ( ~G142 & n468 ) | ( n415 & n468 );
  assign n470 = n419 & ~n469 ;
  assign n471 = ~n412 & n470 ;
  assign n472 = G9 & n471 ;
  assign n473 = ( G120 & G117 ) | ( G120 & ~G51 ) | ( G117 & ~G51 );
  assign n474 = ( ~G120 & G117 ) | ( ~G120 & G62 ) | ( G117 & G62 );
  assign n475 = ~n473 & n474 ;
  assign n476 = ( G120 & ~G117 ) | ( G120 & G73 ) | ( ~G117 & G73 );
  assign n477 = ( G120 & G117 ) | ( G120 & G41 ) | ( G117 & G41 );
  assign n478 = n476 & n477 ;
  assign n479 = n475 | n478 ;
  assign n480 = G118 & ~n268 ;
  assign n481 = ( n225 & ~n479 ) | ( n225 & n480 ) | ( ~n479 & n480 );
  assign n482 = G122 | n481 ;
  assign n483 = ( n225 & n480 ) | ( n225 & ~n481 ) | ( n480 & ~n481 );
  assign n484 = G122 | n483 ;
  assign n485 = ( n479 & n482 ) | ( n479 & ~n484 ) | ( n482 & ~n484 );
  assign n486 = ( G146 & G145 ) | ( G146 & ~G104 ) | ( G145 & ~G104 );
  assign n487 = ( ~G146 & G145 ) | ( ~G146 & G94 ) | ( G145 & G94 );
  assign n488 = ~n486 & n487 ;
  assign n489 = ( G146 & ~G145 ) | ( G146 & G114 ) | ( ~G145 & G114 );
  assign n490 = ( G146 & G145 ) | ( G146 & G84 ) | ( G145 & G84 );
  assign n491 = n489 & n490 ;
  assign n492 = n488 | n491 ;
  assign n493 = n362 & n492 ;
  assign n494 = n362 | n492 ;
  assign n495 = ~n493 & n494 ;
  assign n496 = ( n197 & ~n452 ) | ( n197 & n495 ) | ( ~n452 & n495 );
  assign n497 = ( ~n197 & n452 ) | ( ~n197 & n495 ) | ( n452 & n495 );
  assign n498 = ( ~n495 & n496 ) | ( ~n495 & n497 ) | ( n496 & n497 );
  assign n499 = ~n427 & n438 ;
  assign n500 = n427 & ~n438 ;
  assign n501 = n499 | n500 ;
  assign n502 = ( n177 & ~n190 ) | ( n177 & n286 ) | ( ~n190 & n286 );
  assign n503 = ( ~n177 & n190 ) | ( ~n177 & n502 ) | ( n190 & n502 );
  assign n504 = ( ~n286 & n502 ) | ( ~n286 & n503 ) | ( n502 & n503 );
  assign n505 = ( n498 & n501 ) | ( n498 & ~n504 ) | ( n501 & ~n504 );
  assign n506 = ( n498 & ~n501 ) | ( n498 & n504 ) | ( ~n501 & n504 );
  assign n507 = ( ~n498 & n505 ) | ( ~n498 & n506 ) | ( n505 & n506 );
  assign n508 = ~G29 & n507 ;
  assign n509 = G123 | n479 ;
  assign n510 = ~n253 & n260 ;
  assign n511 = n253 & ~n260 ;
  assign n512 = n510 | n511 ;
  assign n513 = ( ~n204 & n246 ) | ( ~n204 & n512 ) | ( n246 & n512 );
  assign n514 = ( n204 & ~n246 ) | ( n204 & n513 ) | ( ~n246 & n513 );
  assign n515 = ( ~n512 & n513 ) | ( ~n512 & n514 ) | ( n513 & n514 );
  assign n516 = ~n225 & n479 ;
  assign n517 = n225 & ~n479 ;
  assign n518 = n516 | n517 ;
  assign n519 = n240 | n268 ;
  assign n520 = n240 & n268 ;
  assign n521 = n519 & ~n520 ;
  assign n522 = ( n276 & ~n518 ) | ( n276 & n521 ) | ( ~n518 & n521 );
  assign n523 = ( n276 & n521 ) | ( n276 & ~n522 ) | ( n521 & ~n522 );
  assign n524 = ( n518 & n522 ) | ( n518 & ~n523 ) | ( n522 & ~n523 );
  assign n525 = n515 & ~n524 ;
  assign n526 = ( G123 & n515 ) | ( G123 & ~n524 ) | ( n515 & ~n524 );
  assign n527 = ( n509 & n525 ) | ( n509 & ~n526 ) | ( n525 & ~n526 );
  assign n528 = n211 | n218 ;
  assign n529 = n211 & n218 ;
  assign n530 = n528 & ~n529 ;
  assign n531 = ( ~n518 & n521 ) | ( ~n518 & n530 ) | ( n521 & n530 );
  assign n532 = ( n518 & ~n521 ) | ( n518 & n531 ) | ( ~n521 & n531 );
  assign n533 = ( ~n530 & n531 ) | ( ~n530 & n532 ) | ( n531 & n532 );
  assign n534 = n515 & ~n533 ;
  assign n535 = ( G29 & n515 ) | ( G29 & ~n534 ) | ( n515 & ~n534 );
  assign n536 = ( n533 & n534 ) | ( n533 & ~n535 ) | ( n534 & ~n535 );
  assign n537 = G30 & ~n177 ;
  assign n538 = ~G127 & n197 ;
  assign n539 = n537 & ~n538 ;
  assign n540 = n537 & n538 ;
  assign n541 = G138 | n540 ;
  assign n542 = n539 & ~n541 ;
  assign n543 = ~n438 & n539 ;
  assign n544 = n542 & n543 ;
  assign n545 = n542 | n543 ;
  assign n546 = ~n544 & n545 ;
  assign n547 = G135 | n540 ;
  assign n548 = n539 & ~n547 ;
  assign n549 = n362 & n539 ;
  assign n550 = n548 & ~n549 ;
  assign n551 = n548 & ~n550 ;
  assign n552 = n549 | n550 ;
  assign n553 = ( n546 & ~n551 ) | ( n546 & n552 ) | ( ~n551 & n552 );
  assign n554 = ~G136 & n539 ;
  assign n555 = n427 & n539 ;
  assign n556 = n554 & ~n555 ;
  assign n557 = ( n549 & ~n554 ) | ( n549 & n555 ) | ( ~n554 & n555 );
  assign n558 = ( n548 & n556 ) | ( n548 & ~n557 ) | ( n556 & ~n557 );
  assign n559 = ( n542 & ~n543 ) | ( n542 & n558 ) | ( ~n543 & n558 );
  assign n560 = ~n260 & n539 ;
  assign n561 = ~G134 & n539 ;
  assign n562 = ~n560 & n561 ;
  assign n563 = n554 | n555 ;
  assign n564 = ( ~n554 & n556 ) | ( ~n554 & n563 ) | ( n556 & n563 );
  assign n565 = n562 & ~n564 ;
  assign n566 = n559 | n565 ;
  assign n567 = ( ~n553 & n559 ) | ( ~n553 & n566 ) | ( n559 & n566 );
  assign n568 = n561 & ~n562 ;
  assign n569 = n560 | n562 ;
  assign n570 = ( n564 & ~n568 ) | ( n564 & n569 ) | ( ~n568 & n569 );
  assign n571 = ( n553 & ~n567 ) | ( n553 & n570 ) | ( ~n567 & n570 );
  assign n572 = ~G140 & n540 ;
  assign n573 = G129 | n540 ;
  assign n574 = ~n572 & n573 ;
  assign n575 = n218 & ~n574 ;
  assign n576 = ( ~G8 & n246 ) | ( ~G8 & n540 ) | ( n246 & n540 );
  assign n577 = ( ~G132 & G8 ) | ( ~G132 & n540 ) | ( G8 & n540 );
  assign n578 = ~n576 & n577 ;
  assign n579 = ( ~G8 & n253 ) | ( ~G8 & n540 ) | ( n253 & n540 );
  assign n580 = ( ~G133 & G8 ) | ( ~G133 & n540 ) | ( G8 & n540 );
  assign n581 = ~n579 & n580 ;
  assign n582 = n578 | n581 ;
  assign n583 = n575 & ~n582 ;
  assign n584 = ( G141 & ~G8 ) | ( G141 & n540 ) | ( ~G8 & n540 );
  assign n585 = ( ~G130 & G8 ) | ( ~G130 & n540 ) | ( G8 & n540 );
  assign n586 = ~n584 & n585 ;
  assign n587 = ~n211 & n540 ;
  assign n588 = n211 | n540 ;
  assign n589 = ~n587 & n588 ;
  assign n590 = G8 & ~n589 ;
  assign n591 = n586 | n590 ;
  assign n592 = ~n204 & n540 ;
  assign n593 = n204 | n540 ;
  assign n594 = ~n592 & n593 ;
  assign n595 = G8 & ~n594 ;
  assign n596 = ( G142 & ~G8 ) | ( G142 & n540 ) | ( ~G8 & n540 );
  assign n597 = ( ~G131 & G8 ) | ( ~G131 & n540 ) | ( G8 & n540 );
  assign n598 = ~n596 & n597 ;
  assign n599 = n595 & n598 ;
  assign n600 = n595 | n598 ;
  assign n601 = ~n599 & n600 ;
  assign n602 = ( n586 & n590 ) | ( n586 & ~n591 ) | ( n590 & ~n591 );
  assign n603 = ( n591 & n601 ) | ( n591 & ~n602 ) | ( n601 & ~n602 );
  assign n604 = n583 & ~n603 ;
  assign n605 = ( n582 & n586 ) | ( n582 & ~n590 ) | ( n586 & ~n590 );
  assign n606 = ~n582 & n605 ;
  assign n607 = ~n601 & n606 ;
  assign n608 = ~n595 & n598 ;
  assign n609 = G133 & G132 ;
  assign n610 = G8 & ~n609 ;
  assign n611 = ~n540 & n610 ;
  assign n612 = n582 & ~n611 ;
  assign n613 = ( n608 & n611 ) | ( n608 & ~n612 ) | ( n611 & ~n612 );
  assign n614 = n607 | n613 ;
  assign n615 = n604 | n614 ;
  assign n616 = n571 | n615 ;
  assign n617 = ( ~n218 & n574 ) | ( ~n218 & n578 ) | ( n574 & n578 );
  assign n618 = n575 | n617 ;
  assign n619 = ( n581 & ~n603 ) | ( n581 & n618 ) | ( ~n603 & n618 );
  assign n620 = ~G138 & n540 ;
  assign n621 = G126 | n540 ;
  assign n622 = ~n620 & n621 ;
  assign n623 = n268 | n622 ;
  assign n624 = ~G139 & n540 ;
  assign n625 = G128 | n540 ;
  assign n626 = ~n624 & n625 ;
  assign n627 = ( ~n240 & n623 ) | ( ~n240 & n626 ) | ( n623 & n626 );
  assign n628 = n268 & n622 ;
  assign n629 = ( G136 & n225 ) | ( G136 & n540 ) | ( n225 & n540 );
  assign n630 = ( G125 & n225 ) | ( G125 & ~n540 ) | ( n225 & ~n540 );
  assign n631 = n629 | n630 ;
  assign n632 = n626 | n631 ;
  assign n633 = n240 & ~n631 ;
  assign n634 = ( n628 & n632 ) | ( n628 & ~n633 ) | ( n632 & ~n633 );
  assign n635 = n627 & n634 ;
  assign n636 = n603 | n635 ;
  assign n637 = n619 | n636 ;
  assign n638 = ( ~n567 & n571 ) | ( ~n567 & n637 ) | ( n571 & n637 );
  assign n639 = ~n567 & n571 ;
  assign n640 = ( ~n616 & n638 ) | ( ~n616 & n639 ) | ( n638 & n639 );
  assign n641 = ~n312 & n348 ;
  assign n642 = n327 & ~n536 ;
  assign n643 = n641 & n642 ;
  assign n644 = ~n170 & n643 ;
  assign n645 = G29 & n325 ;
  assign n646 = G29 & ~n324 ;
  assign n647 = ( n326 & n645 ) | ( n326 & n646 ) | ( n645 & n646 );
  assign n648 = n641 & n647 ;
  assign n649 = ~n170 & n648 ;
  assign n650 = ( ~n507 & n644 ) | ( ~n507 & n649 ) | ( n644 & n649 );
  assign G2551 = ~n158 ;
  assign G2552 = ~n159 ;
  assign G2553 = ~n160 ;
  assign G2554 = ~n167 ;
  assign G2555 = ~n167 ;
  assign G2556 = n170 ;
  assign G2557 = ~n177 ;
  assign G2531 = ~G115 ;
  assign G2532 = ~G115 ;
  assign G2533 = ~G115 ;
  assign G2534 = ~G124 ;
  assign G2535 = ~G124 ;
  assign G2536 = ~G137 ;
  assign G2537 = ~G137 ;
  assign G2538 = ~G137 ;
  assign G2539 = ~G32 ;
  assign G2540 = ~G106 ;
  assign G2541 = ~G64 ;
  assign G2542 = ~G76 ;
  assign G2543 = ~G53 ;
  assign G2544 = ~G96 ;
  assign G2545 = ~G43 ;
  assign G2546 = ~G86 ;
  assign G2547 = ~n180 ;
  assign G2548 = ~n182 ;
  assign G2549 = G115 ;
  assign G2550 = n183 ;
  assign G2558 = ~n190 ;
  assign G2559 = ~n197 ;
  assign G2560 = ~n204 ;
  assign G2561 = ~n211 ;
  assign G2562 = ~n218 ;
  assign G2563 = ~n227 ;
  assign G2564 = ~n230 ;
  assign G2565 = ~n233 ;
  assign G2566 = n240 ;
  assign G2567 = n218 ;
  assign G2568 = n211 ;
  assign G2569 = n204 ;
  assign G2570 = n246 ;
  assign G2571 = n253 ;
  assign G2572 = n260 ;
  assign G2573 = ~n270 ;
  assign G2574 = ~n270 ;
  assign G2575 = n273 ;
  assign G2576 = n273 ;
  assign G2577 = n275 ;
  assign G2578 = ~n279 ;
  assign G2579 = ~n279 ;
  assign G2580 = ~n289 ;
  assign G2581 = ~n312 ;
  assign G2582 = ~n327 ;
  assign G2583 = ~n348 ;
  assign G2584 = ~n472 ;
  assign G2585 = ~n472 ;
  assign G2586 = n485 ;
  assign G2587 = ~n508 ;
  assign G2588 = n527 ;
  assign G2589 = n527 ;
  assign G2590 = ~n536 ;
  assign G2591 = n640 ;
  assign G2592 = 1'b0 ;
  assign G2593 = ~n650 ;
  assign G2594 = ~n650 ;
endmodule
