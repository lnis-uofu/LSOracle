module top(G7 , G121 , G119 , G147 , G53 , G86 , G43 , G96 , G32 , G76 , G64 , G106 , G146 , G145 , G89 , G99 , G79 , G109 , G115 , G124 , G137 , G139 , G140 , G141 , G142 , G11 , G2 , G74 , G88 , G98 , G78 , G108 , G90 , G100 , G80 , G110 , G120 , G117 , G57 , G46 , G36 , G68 , G58 , G47 , G37 , G69 , G59 , G48 , G38 , G70 , G122 , G52 , G42 , G31 , G63 , G28 , G116 , G1 , G3 , G60 , G49 , G39 , G71 , G56 , G35 , G67 , G55 , G45 , G34 , G66 , G54 , G44 , G33 , G65 , G61 , G50 , G40 , G72 , G123 , G118 , G144 , G143 , G87 , G97 , G77 , G107 , G155 , G154 , G125 , G126 , G153 , G152 , G151 , G150 , G149 , G148 , G10 , G157 , G138 , G133 , G134 , G135 , G136 , G131 , G132 , G129 , G130 , G156 , G128 , G9 , G22 , G23 , G27 , G24 , G93 , G103 , G83 , G113 , G20 , G92 , G102 , G82 , G112 , G25 , G91 , G101 , G81 , G111 , G21 , G26 , G16 , G12 , G17 , G6 , G18 , G19 , G85 , G95 , G75 , G105 , G13 , G4 , G14 , G5 , G15 , G62 , G51 , G41 , G73 , G94 , G104 , G84 , G114 , G29 , G30 , G127 , G8 , G2551 , G2552 , G2553 , G2554 , G2555 , G2556 , G2557 , G2531 , G2532 , G2533 , G2534 , G2535 , G2536 , G2537 , G2538 , G2539 , G2540 , G2541 , G2542 , G2543 , G2544 , G2545 , G2546 , G2547 , G2548 , G2549 , G2550 , G2558 , G2559 , G2560 , G2561 , G2562 , G2563 , G2564 , G2565 , G2566 , G2567 , G2568 , G2569 , G2570 , G2571 , G2572 , G2573 , G2574 , G2575 , G2576 , G2577 , G2578 , G2579 , G2580 , G2581 , G2582 , G2583 , G2584 , G2585 , G2586 , G2587 , G2588 , G2589 , G2590 , G2591 , G2592 , G2593 , G2594 );
  input G7 , G121 , G119 , G147 , G53 , G86 , G43 , G96 , G32 , G76 , G64 , G106 , G146 , G145 , G89 , G99 , G79 , G109 , G115 , G124 , G137 , G139 , G140 , G141 , G142 , G11 , G2 , G74 , G88 , G98 , G78 , G108 , G90 , G100 , G80 , G110 , G120 , G117 , G57 , G46 , G36 , G68 , G58 , G47 , G37 , G69 , G59 , G48 , G38 , G70 , G122 , G52 , G42 , G31 , G63 , G28 , G116 , G1 , G3 , G60 , G49 , G39 , G71 , G56 , G35 , G67 , G55 , G45 , G34 , G66 , G54 , G44 , G33 , G65 , G61 , G50 , G40 , G72 , G123 , G118 , G144 , G143 , G87 , G97 , G77 , G107 , G155 , G154 , G125 , G126 , G153 , G152 , G151 , G150 , G149 , G148 , G10 , G157 , G138 , G133 , G134 , G135 , G136 , G131 , G132 , G129 , G130 , G156 , G128 , G9 , G22 , G23 , G27 , G24 , G93 , G103 , G83 , G113 , G20 , G92 , G102 , G82 , G112 , G25 , G91 , G101 , G81 , G111 , G21 , G26 , G16 , G12 , G17 , G6 , G18 , G19 , G85 , G95 , G75 , G105 , G13 , G4 , G14 , G5 , G15 , G62 , G51 , G41 , G73 , G94 , G104 , G84 , G114 , G29 , G30 , G127 , G8 ;
  output G2551 , G2552 , G2553 , G2554 , G2555 , G2556 , G2557 , G2531 , G2532 , G2533 , G2534 , G2535 , G2536 , G2537 , G2538 , G2539 , G2540 , G2541 , G2542 , G2543 , G2544 , G2545 , G2546 , G2547 , G2548 , G2549 , G2550 , G2558 , G2559 , G2560 , G2561 , G2562 , G2563 , G2564 , G2565 , G2566 , G2567 , G2568 , G2569 , G2570 , G2571 , G2572 , G2573 , G2574 , G2575 , G2576 , G2577 , G2578 , G2579 , G2580 , G2581 , G2582 , G2583 , G2584 , G2585 , G2586 , G2587 , G2588 , G2589 , G2590 , G2591 , G2592 , G2593 , G2594 ;
  wire n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873;
  assign n158 = G7 & G121 ;
  assign n159 = G119 & n158 ;
  assign n160 = G147 & n158 ;
  assign n161 = G53 & G86 ;
  assign n162 = G43 & G96 ;
  assign n163 = n161 & n162 ;
  assign n164 = G32 & G76 ;
  assign n165 = G64 & G106 ;
  assign n166 = n164 & n165 ;
  assign n167 = n163 & n166 ;
  assign n168 = G147 & ~n166 ;
  assign n169 = G119 & ~n163 ;
  assign n170 = ~n168 & ~n169 ;
  assign n171 = ~G145 & G89 ;
  assign n172 = ~G146 & n171 ;
  assign n173 = G145 & G99 ;
  assign n174 = ~G146 & n173 ;
  assign n175 = ~n172 & ~n174 ;
  assign n176 = ~G145 & G79 ;
  assign n177 = G146 & n176 ;
  assign n178 = G145 & G109 ;
  assign n179 = G146 & n178 ;
  assign n180 = ~n177 & ~n179 ;
  assign n181 = n175 & n180 ;
  assign n182 = G139 & G140 ;
  assign n183 = G141 & G142 ;
  assign n184 = n182 & n183 ;
  assign n185 = G11 & G2 ;
  assign n186 = G121 & n185 ;
  assign n187 = ~G115 & G74 ;
  assign n188 = ~G145 & G88 ;
  assign n189 = ~G146 & n188 ;
  assign n190 = G145 & G98 ;
  assign n191 = ~G146 & n190 ;
  assign n192 = ~n189 & ~n191 ;
  assign n193 = ~G145 & G78 ;
  assign n194 = G146 & n193 ;
  assign n195 = G145 & G108 ;
  assign n196 = G146 & n195 ;
  assign n197 = ~n194 & ~n196 ;
  assign n198 = n192 & n197 ;
  assign n199 = ~G145 & G90 ;
  assign n200 = ~G146 & n199 ;
  assign n201 = G145 & G100 ;
  assign n202 = ~G146 & n201 ;
  assign n203 = ~n200 & ~n202 ;
  assign n204 = ~G145 & G80 ;
  assign n205 = G146 & n204 ;
  assign n206 = G145 & G110 ;
  assign n207 = G146 & n206 ;
  assign n208 = ~n205 & ~n207 ;
  assign n209 = n203 & n208 ;
  assign n210 = ~G117 & G57 ;
  assign n211 = ~G120 & n210 ;
  assign n212 = G117 & G46 ;
  assign n213 = ~G120 & n212 ;
  assign n214 = ~n211 & ~n213 ;
  assign n215 = ~G117 & G36 ;
  assign n216 = G120 & n215 ;
  assign n217 = G117 & G68 ;
  assign n218 = G120 & n217 ;
  assign n219 = ~n216 & ~n218 ;
  assign n220 = n214 & n219 ;
  assign n221 = ~G117 & G58 ;
  assign n222 = ~G120 & n221 ;
  assign n223 = G117 & G47 ;
  assign n224 = ~G120 & n223 ;
  assign n225 = ~n222 & ~n224 ;
  assign n226 = ~G117 & G37 ;
  assign n227 = G120 & n226 ;
  assign n228 = G117 & G69 ;
  assign n229 = G120 & n228 ;
  assign n230 = ~n227 & ~n229 ;
  assign n231 = n225 & n230 ;
  assign n232 = ~G117 & G59 ;
  assign n233 = ~G120 & n232 ;
  assign n234 = G117 & G48 ;
  assign n235 = ~G120 & n234 ;
  assign n236 = ~n233 & ~n235 ;
  assign n237 = ~G117 & G38 ;
  assign n238 = G120 & n237 ;
  assign n239 = G117 & G70 ;
  assign n240 = G120 & n239 ;
  assign n241 = ~n238 & ~n240 ;
  assign n242 = n236 & n241 ;
  assign n243 = ~G117 & G52 ;
  assign n244 = ~G120 & n243 ;
  assign n245 = G117 & G42 ;
  assign n246 = ~G120 & n245 ;
  assign n247 = ~n244 & ~n246 ;
  assign n248 = ~G117 & G31 ;
  assign n249 = G120 & n248 ;
  assign n250 = G117 & G63 ;
  assign n251 = G120 & n250 ;
  assign n252 = ~n249 & ~n251 ;
  assign n253 = n247 & n252 ;
  assign n254 = G122 & ~n253 ;
  assign n255 = G122 & ~n254 ;
  assign n256 = G28 & n170 ;
  assign n257 = ~G121 & G116 ;
  assign n258 = n256 & n257 ;
  assign n259 = G1 & G3 ;
  assign n260 = n170 & ~n259 ;
  assign n261 = n257 & n260 ;
  assign n262 = ~G117 & G60 ;
  assign n263 = ~G120 & n262 ;
  assign n264 = G117 & G49 ;
  assign n265 = ~G120 & n264 ;
  assign n266 = ~n263 & ~n265 ;
  assign n267 = ~G117 & G39 ;
  assign n268 = G120 & n267 ;
  assign n269 = G117 & G71 ;
  assign n270 = G120 & n269 ;
  assign n271 = ~n268 & ~n270 ;
  assign n272 = n266 & n271 ;
  assign n273 = ~G117 & G56 ;
  assign n274 = ~G120 & n273 ;
  assign n275 = ~G120 & G117 ;
  assign n276 = ~n274 & ~n275 ;
  assign n277 = ~G117 & G35 ;
  assign n278 = G120 & n277 ;
  assign n279 = G117 & G67 ;
  assign n280 = G120 & n279 ;
  assign n281 = ~n278 & ~n280 ;
  assign n282 = n276 & n281 ;
  assign n283 = ~G117 & G55 ;
  assign n284 = ~G120 & n283 ;
  assign n285 = G117 & G45 ;
  assign n286 = ~G120 & n285 ;
  assign n287 = ~n284 & ~n286 ;
  assign n288 = ~G117 & G34 ;
  assign n289 = G120 & n288 ;
  assign n290 = G117 & G66 ;
  assign n291 = G120 & n290 ;
  assign n292 = ~n289 & ~n291 ;
  assign n293 = n287 & n292 ;
  assign n294 = ~G117 & G54 ;
  assign n295 = ~G120 & n294 ;
  assign n296 = G117 & G44 ;
  assign n297 = ~G120 & n296 ;
  assign n298 = ~n295 & ~n297 ;
  assign n299 = ~G117 & G33 ;
  assign n300 = G120 & n299 ;
  assign n301 = G117 & G65 ;
  assign n302 = G120 & n301 ;
  assign n303 = ~n300 & ~n302 ;
  assign n304 = n298 & n303 ;
  assign n305 = ~G117 & G61 ;
  assign n306 = ~G120 & n305 ;
  assign n307 = G117 & G50 ;
  assign n308 = ~G120 & n307 ;
  assign n309 = ~n306 & ~n308 ;
  assign n310 = ~G117 & G40 ;
  assign n311 = G120 & n310 ;
  assign n312 = G117 & G72 ;
  assign n313 = G120 & n312 ;
  assign n314 = ~n311 & ~n313 ;
  assign n315 = n309 & n314 ;
  assign n316 = ~G123 & ~n315 ;
  assign n317 = G123 & n242 ;
  assign n318 = ~n316 & ~n317 ;
  assign n319 = ~G123 & n272 ;
  assign n320 = G123 & ~n231 ;
  assign n321 = ~n319 & ~n320 ;
  assign n322 = ~G118 & n315 ;
  assign n323 = ~G122 & ~n322 ;
  assign n324 = G122 & ~n315 ;
  assign n325 = ~n323 & ~n324 ;
  assign n326 = ~G123 & ~n253 ;
  assign n327 = G123 & ~n322 ;
  assign n328 = ~n326 & ~n327 ;
  assign n329 = ~G146 & ~G145 ;
  assign n330 = ~G146 & G145 ;
  assign n331 = ~n329 & ~n330 ;
  assign n332 = G146 & ~G145 ;
  assign n333 = G146 & G145 ;
  assign n334 = ~n332 & ~n333 ;
  assign n335 = n331 & n334 ;
  assign n336 = ~G144 & ~n335 ;
  assign n337 = ~G144 & ~n336 ;
  assign n338 = ~n335 & ~n336 ;
  assign n339 = ~n337 & ~n338 ;
  assign n340 = ~G145 & G87 ;
  assign n341 = ~G146 & n340 ;
  assign n342 = G145 & G97 ;
  assign n343 = ~G146 & n342 ;
  assign n344 = ~n341 & ~n343 ;
  assign n345 = ~G145 & G77 ;
  assign n346 = G146 & n345 ;
  assign n347 = G145 & G107 ;
  assign n348 = G146 & n347 ;
  assign n349 = ~n346 & ~n348 ;
  assign n350 = n344 & n349 ;
  assign n351 = ~G143 & ~n350 ;
  assign n352 = ~G143 & ~n351 ;
  assign n353 = ~n350 & ~n351 ;
  assign n354 = ~n352 & ~n353 ;
  assign n355 = n339 & n354 ;
  assign n356 = G155 & ~G154 ;
  assign n357 = ~G155 & G154 ;
  assign n358 = ~n356 & ~n357 ;
  assign n359 = ~G125 & G126 ;
  assign n360 = G125 & ~G126 ;
  assign n361 = ~n359 & ~n360 ;
  assign n362 = ~n358 & n361 ;
  assign n363 = n358 & ~n361 ;
  assign n364 = ~n362 & ~n363 ;
  assign n365 = G153 & ~G152 ;
  assign n366 = ~G153 & G152 ;
  assign n367 = ~n365 & ~n366 ;
  assign n368 = G151 & ~G150 ;
  assign n369 = ~G151 & G150 ;
  assign n370 = ~n368 & ~n369 ;
  assign n371 = G149 & ~G148 ;
  assign n372 = ~G149 & G148 ;
  assign n373 = ~n371 & ~n372 ;
  assign n374 = n370 & ~n373 ;
  assign n375 = ~n367 & n374 ;
  assign n376 = n370 & n373 ;
  assign n377 = n367 & n376 ;
  assign n378 = ~n375 & ~n377 ;
  assign n379 = ~n370 & n373 ;
  assign n380 = ~n367 & n379 ;
  assign n381 = ~n370 & ~n373 ;
  assign n382 = n367 & n381 ;
  assign n383 = ~n380 & ~n382 ;
  assign n384 = n378 & n383 ;
  assign n385 = ~n364 & n384 ;
  assign n386 = n364 & ~n384 ;
  assign n387 = ~n385 & ~n386 ;
  assign n388 = G10 & n387 ;
  assign n389 = G144 & ~G143 ;
  assign n390 = ~G144 & G143 ;
  assign n391 = ~n389 & ~n390 ;
  assign n392 = ~G141 & G142 ;
  assign n393 = G141 & ~G142 ;
  assign n394 = ~n392 & ~n393 ;
  assign n395 = ~G139 & G140 ;
  assign n396 = G139 & ~G140 ;
  assign n397 = ~n395 & ~n396 ;
  assign n398 = G157 & G138 ;
  assign n399 = ~G157 & ~G138 ;
  assign n400 = ~n398 & ~n399 ;
  assign n401 = n397 & ~n400 ;
  assign n402 = ~n394 & n401 ;
  assign n403 = n397 & n400 ;
  assign n404 = n394 & n403 ;
  assign n405 = ~n402 & ~n404 ;
  assign n406 = ~n397 & n400 ;
  assign n407 = ~n394 & n406 ;
  assign n408 = ~n397 & ~n400 ;
  assign n409 = n394 & n408 ;
  assign n410 = ~n407 & ~n409 ;
  assign n411 = n405 & n410 ;
  assign n412 = ~n391 & n411 ;
  assign n413 = n391 & ~n411 ;
  assign n414 = ~n412 & ~n413 ;
  assign n415 = ~G133 & G134 ;
  assign n416 = G133 & ~G134 ;
  assign n417 = ~n415 & ~n416 ;
  assign n418 = ~G135 & G136 ;
  assign n419 = G135 & ~G136 ;
  assign n420 = ~n418 & ~n419 ;
  assign n421 = ~n417 & n420 ;
  assign n422 = n417 & ~n420 ;
  assign n423 = ~n421 & ~n422 ;
  assign n424 = ~G131 & G132 ;
  assign n425 = G131 & ~G132 ;
  assign n426 = ~n424 & ~n425 ;
  assign n427 = ~G129 & G130 ;
  assign n428 = G129 & ~G130 ;
  assign n429 = ~n427 & ~n428 ;
  assign n430 = G156 & G128 ;
  assign n431 = ~G156 & ~G128 ;
  assign n432 = ~n430 & ~n431 ;
  assign n433 = n429 & ~n432 ;
  assign n434 = ~n426 & n433 ;
  assign n435 = n429 & n432 ;
  assign n436 = n426 & n435 ;
  assign n437 = ~n434 & ~n436 ;
  assign n438 = ~n429 & n432 ;
  assign n439 = ~n426 & n438 ;
  assign n440 = ~n429 & ~n432 ;
  assign n441 = n426 & n440 ;
  assign n442 = ~n439 & ~n441 ;
  assign n443 = n437 & n442 ;
  assign n444 = ~n423 & n443 ;
  assign n445 = n423 & ~n443 ;
  assign n446 = ~n444 & ~n445 ;
  assign n447 = ~G123 & G9 ;
  assign n448 = G123 & G9 ;
  assign n449 = ~n447 & ~n448 ;
  assign n450 = G22 & G23 ;
  assign n451 = ~G23 & ~n350 ;
  assign n452 = ~n450 & ~n451 ;
  assign n453 = G23 & G27 ;
  assign n454 = ~G23 & ~n198 ;
  assign n455 = ~n453 & ~n454 ;
  assign n456 = ~G142 & ~n455 ;
  assign n457 = G142 & n455 ;
  assign n458 = ~n456 & ~n457 ;
  assign n459 = ~n452 & n458 ;
  assign n460 = G23 & G24 ;
  assign n461 = ~G145 & G93 ;
  assign n462 = ~G146 & n461 ;
  assign n463 = G145 & G103 ;
  assign n464 = ~G146 & n463 ;
  assign n465 = ~n462 & ~n464 ;
  assign n466 = ~G145 & G83 ;
  assign n467 = G146 & n466 ;
  assign n468 = G145 & G113 ;
  assign n469 = G146 & n468 ;
  assign n470 = ~n467 & ~n469 ;
  assign n471 = n465 & n470 ;
  assign n472 = ~G23 & ~n471 ;
  assign n473 = ~n460 & ~n472 ;
  assign n474 = ~G136 & ~n473 ;
  assign n475 = G136 & n473 ;
  assign n476 = ~n474 & ~n475 ;
  assign n477 = G23 & G20 ;
  assign n478 = ~G145 & G92 ;
  assign n479 = ~G146 & n478 ;
  assign n480 = G145 & G102 ;
  assign n481 = ~G146 & n480 ;
  assign n482 = ~n479 & ~n481 ;
  assign n483 = ~G145 & G82 ;
  assign n484 = G146 & n483 ;
  assign n485 = G145 & G112 ;
  assign n486 = G146 & n485 ;
  assign n487 = ~n484 & ~n486 ;
  assign n488 = n482 & n487 ;
  assign n489 = ~G23 & ~n488 ;
  assign n490 = ~n477 & ~n489 ;
  assign n491 = ~G138 & ~n490 ;
  assign n492 = G138 & n490 ;
  assign n493 = ~n491 & ~n492 ;
  assign n494 = n476 & n493 ;
  assign n495 = G23 & G25 ;
  assign n496 = ~G145 & G91 ;
  assign n497 = ~G146 & n496 ;
  assign n498 = G145 & G101 ;
  assign n499 = ~G146 & n498 ;
  assign n500 = ~n497 & ~n499 ;
  assign n501 = ~G145 & G81 ;
  assign n502 = G146 & n501 ;
  assign n503 = G145 & G111 ;
  assign n504 = G146 & n503 ;
  assign n505 = ~n502 & ~n504 ;
  assign n506 = n500 & n505 ;
  assign n507 = ~G23 & ~n506 ;
  assign n508 = ~n495 & ~n507 ;
  assign n509 = ~G139 & ~n508 ;
  assign n510 = G139 & n508 ;
  assign n511 = ~n509 & ~n510 ;
  assign n512 = G23 & G21 ;
  assign n513 = ~G23 & ~n209 ;
  assign n514 = ~n512 & ~n513 ;
  assign n515 = ~G140 & ~n514 ;
  assign n516 = G140 & n514 ;
  assign n517 = ~n515 & ~n516 ;
  assign n518 = G23 & G26 ;
  assign n519 = ~G23 & ~n181 ;
  assign n520 = ~n518 & ~n519 ;
  assign n521 = ~G141 & ~n520 ;
  assign n522 = G141 & n520 ;
  assign n523 = ~n521 & ~n522 ;
  assign n524 = n517 & n523 ;
  assign n525 = n511 & n524 ;
  assign n526 = n494 & n525 ;
  assign n527 = n459 & n526 ;
  assign n528 = G16 & G12 ;
  assign n529 = ~G12 & ~n220 ;
  assign n530 = ~n528 & ~n529 ;
  assign n531 = ~G131 & ~n530 ;
  assign n532 = G131 & n530 ;
  assign n533 = ~n531 & ~n532 ;
  assign n534 = G12 & G17 ;
  assign n535 = ~G12 & ~n282 ;
  assign n536 = ~n534 & ~n535 ;
  assign n537 = ~G132 & ~n536 ;
  assign n538 = G132 & n536 ;
  assign n539 = ~n537 & ~n538 ;
  assign n540 = n533 & n539 ;
  assign n541 = G12 & G6 ;
  assign n542 = ~G12 & ~n293 ;
  assign n543 = ~n541 & ~n542 ;
  assign n544 = ~G133 & ~n543 ;
  assign n545 = G133 & n543 ;
  assign n546 = ~n544 & ~n545 ;
  assign n547 = G12 & G18 ;
  assign n548 = ~G12 & ~n304 ;
  assign n549 = ~n547 & ~n548 ;
  assign n550 = ~G134 & ~n549 ;
  assign n551 = G134 & n549 ;
  assign n552 = ~n550 & ~n551 ;
  assign n553 = G23 & G19 ;
  assign n554 = ~G145 & G85 ;
  assign n555 = ~G146 & n554 ;
  assign n556 = G145 & G95 ;
  assign n557 = ~G146 & n556 ;
  assign n558 = ~n555 & ~n557 ;
  assign n559 = ~G145 & G75 ;
  assign n560 = G146 & n559 ;
  assign n561 = G145 & G105 ;
  assign n562 = G146 & n561 ;
  assign n563 = ~n560 & ~n562 ;
  assign n564 = n558 & n563 ;
  assign n565 = ~G23 & ~n564 ;
  assign n566 = ~n553 & ~n565 ;
  assign n567 = ~G135 & ~n566 ;
  assign n568 = G135 & n566 ;
  assign n569 = ~n567 & ~n568 ;
  assign n570 = n552 & n569 ;
  assign n571 = n546 & n570 ;
  assign n572 = n540 & n571 ;
  assign n573 = G12 & G13 ;
  assign n574 = ~G12 & ~n253 ;
  assign n575 = ~n573 & ~n574 ;
  assign n576 = ~G125 & ~n575 ;
  assign n577 = G125 & n575 ;
  assign n578 = ~n576 & ~n577 ;
  assign n579 = G12 & G4 ;
  assign n580 = ~G12 & ~n315 ;
  assign n581 = ~n579 & ~n580 ;
  assign n582 = ~G126 & ~n581 ;
  assign n583 = G126 & n581 ;
  assign n584 = ~n582 & ~n583 ;
  assign n585 = n578 & n584 ;
  assign n586 = G12 & G14 ;
  assign n587 = ~G12 & ~n272 ;
  assign n588 = ~n586 & ~n587 ;
  assign n589 = ~G128 & ~n588 ;
  assign n590 = G128 & n588 ;
  assign n591 = ~n589 & ~n590 ;
  assign n592 = G12 & G5 ;
  assign n593 = ~G12 & ~n242 ;
  assign n594 = ~n592 & ~n593 ;
  assign n595 = ~G129 & ~n594 ;
  assign n596 = G129 & n594 ;
  assign n597 = ~n595 & ~n596 ;
  assign n598 = G12 & G15 ;
  assign n599 = ~G12 & ~n231 ;
  assign n600 = ~n598 & ~n599 ;
  assign n601 = ~G130 & ~n600 ;
  assign n602 = G130 & n600 ;
  assign n603 = ~n601 & ~n602 ;
  assign n604 = n597 & n603 ;
  assign n605 = n591 & n604 ;
  assign n606 = n585 & n605 ;
  assign n607 = n572 & n606 ;
  assign n608 = n527 & n607 ;
  assign n609 = ~n449 & n608 ;
  assign n610 = n253 & n315 ;
  assign n611 = ~n253 & ~n315 ;
  assign n612 = ~n610 & ~n611 ;
  assign n613 = ~n322 & ~n612 ;
  assign n614 = n322 & n612 ;
  assign n615 = ~n613 & ~n614 ;
  assign n616 = ~G117 & G62 ;
  assign n617 = ~G120 & n616 ;
  assign n618 = G117 & G51 ;
  assign n619 = ~G120 & n618 ;
  assign n620 = ~n617 & ~n619 ;
  assign n621 = ~G117 & G41 ;
  assign n622 = G120 & n621 ;
  assign n623 = G117 & G73 ;
  assign n624 = G120 & n623 ;
  assign n625 = ~n622 & ~n624 ;
  assign n626 = n620 & n625 ;
  assign n627 = ~n615 & n626 ;
  assign n628 = n615 & ~n626 ;
  assign n629 = ~n627 & ~n628 ;
  assign n630 = ~G122 & ~n629 ;
  assign n631 = G122 & ~n626 ;
  assign n632 = ~n630 & ~n631 ;
  assign n633 = n181 & ~n198 ;
  assign n634 = ~n181 & n198 ;
  assign n635 = ~n633 & ~n634 ;
  assign n636 = ~n335 & n350 ;
  assign n637 = n335 & ~n350 ;
  assign n638 = ~n636 & ~n637 ;
  assign n639 = ~n635 & n638 ;
  assign n640 = n635 & ~n638 ;
  assign n641 = ~n639 & ~n640 ;
  assign n642 = ~n209 & n506 ;
  assign n643 = n209 & ~n506 ;
  assign n644 = ~n642 & ~n643 ;
  assign n645 = n471 & ~n488 ;
  assign n646 = ~n471 & n488 ;
  assign n647 = ~n645 & ~n646 ;
  assign n648 = ~G145 & G94 ;
  assign n649 = ~G146 & n648 ;
  assign n650 = G145 & G104 ;
  assign n651 = ~G146 & n650 ;
  assign n652 = ~n649 & ~n651 ;
  assign n653 = ~G145 & G84 ;
  assign n654 = G146 & n653 ;
  assign n655 = G145 & G114 ;
  assign n656 = G146 & n655 ;
  assign n657 = ~n654 & ~n656 ;
  assign n658 = n652 & n657 ;
  assign n659 = ~n564 & ~n658 ;
  assign n660 = n564 & n658 ;
  assign n661 = ~n659 & ~n660 ;
  assign n662 = n647 & ~n661 ;
  assign n663 = ~n644 & n662 ;
  assign n664 = n647 & n661 ;
  assign n665 = n644 & n664 ;
  assign n666 = ~n663 & ~n665 ;
  assign n667 = ~n647 & n661 ;
  assign n668 = ~n644 & n667 ;
  assign n669 = ~n647 & ~n661 ;
  assign n670 = n644 & n669 ;
  assign n671 = ~n668 & ~n670 ;
  assign n672 = n666 & n671 ;
  assign n673 = ~n641 & n672 ;
  assign n674 = n641 & ~n672 ;
  assign n675 = ~n673 & ~n674 ;
  assign n676 = ~G29 & n675 ;
  assign n677 = ~G123 & n626 ;
  assign n678 = n220 & ~n282 ;
  assign n679 = ~n220 & n282 ;
  assign n680 = ~n678 & ~n679 ;
  assign n681 = n293 & ~n304 ;
  assign n682 = ~n293 & n304 ;
  assign n683 = ~n681 & ~n682 ;
  assign n684 = ~n680 & n683 ;
  assign n685 = n680 & ~n683 ;
  assign n686 = ~n684 & ~n685 ;
  assign n687 = ~n272 & ~n315 ;
  assign n688 = n272 & n315 ;
  assign n689 = ~n687 & ~n688 ;
  assign n690 = n253 & ~n626 ;
  assign n691 = ~n253 & n626 ;
  assign n692 = ~n690 & ~n691 ;
  assign n693 = n322 & n692 ;
  assign n694 = ~n689 & n693 ;
  assign n695 = ~n322 & n692 ;
  assign n696 = n689 & n695 ;
  assign n697 = ~n694 & ~n696 ;
  assign n698 = ~n322 & ~n692 ;
  assign n699 = ~n689 & n698 ;
  assign n700 = n322 & ~n692 ;
  assign n701 = n689 & n700 ;
  assign n702 = ~n699 & ~n701 ;
  assign n703 = n697 & n702 ;
  assign n704 = ~n686 & n703 ;
  assign n705 = n686 & ~n703 ;
  assign n706 = ~n704 & ~n705 ;
  assign n707 = G123 & ~n706 ;
  assign n708 = ~n677 & ~n707 ;
  assign n709 = n231 & n242 ;
  assign n710 = ~n231 & ~n242 ;
  assign n711 = ~n709 & ~n710 ;
  assign n712 = n689 & ~n692 ;
  assign n713 = ~n711 & n712 ;
  assign n714 = n689 & n692 ;
  assign n715 = n711 & n714 ;
  assign n716 = ~n713 & ~n715 ;
  assign n717 = ~n689 & n692 ;
  assign n718 = ~n711 & n717 ;
  assign n719 = ~n689 & ~n692 ;
  assign n720 = n711 & n719 ;
  assign n721 = ~n718 & ~n720 ;
  assign n722 = n716 & n721 ;
  assign n723 = ~n686 & n722 ;
  assign n724 = n686 & ~n722 ;
  assign n725 = ~n723 & ~n724 ;
  assign n726 = ~G29 & n725 ;
  assign n727 = ~G127 & ~n209 ;
  assign n728 = n181 & n727 ;
  assign n729 = G30 & n728 ;
  assign n730 = ~n471 & ~n729 ;
  assign n731 = G30 & n181 ;
  assign n732 = ~n727 & n731 ;
  assign n733 = n730 & n732 ;
  assign n734 = ~G136 & ~n729 ;
  assign n735 = n732 & n734 ;
  assign n736 = n733 & n735 ;
  assign n737 = ~n733 & ~n735 ;
  assign n738 = ~n736 & ~n737 ;
  assign n739 = n304 & ~n729 ;
  assign n740 = n732 & n739 ;
  assign n741 = ~G134 & ~n729 ;
  assign n742 = n732 & n741 ;
  assign n743 = ~n740 & n742 ;
  assign n744 = ~n738 & n743 ;
  assign n745 = n488 & ~n729 ;
  assign n746 = n732 & n745 ;
  assign n747 = ~G138 & ~n729 ;
  assign n748 = n732 & n747 ;
  assign n749 = n746 & n748 ;
  assign n750 = ~n746 & ~n748 ;
  assign n751 = ~n749 & ~n750 ;
  assign n752 = ~n564 & ~n729 ;
  assign n753 = n732 & n752 ;
  assign n754 = ~G135 & ~n729 ;
  assign n755 = n732 & n754 ;
  assign n756 = n753 & n755 ;
  assign n757 = ~n753 & ~n755 ;
  assign n758 = ~n756 & ~n757 ;
  assign n759 = ~n751 & ~n758 ;
  assign n760 = n744 & n759 ;
  assign n761 = ~n753 & n755 ;
  assign n762 = ~n738 & ~n751 ;
  assign n763 = n761 & n762 ;
  assign n764 = ~n760 & ~n763 ;
  assign n765 = ~n733 & n735 ;
  assign n766 = ~n751 & n765 ;
  assign n767 = ~n746 & n748 ;
  assign n768 = ~n766 & ~n767 ;
  assign n769 = n764 & n768 ;
  assign n770 = n282 & n729 ;
  assign n771 = G8 & n770 ;
  assign n772 = ~G132 & ~n729 ;
  assign n773 = G8 & n772 ;
  assign n774 = n771 & n773 ;
  assign n775 = ~n771 & ~n773 ;
  assign n776 = ~n774 & ~n775 ;
  assign n777 = ~G140 & n729 ;
  assign n778 = ~G129 & ~n729 ;
  assign n779 = ~n777 & ~n778 ;
  assign n780 = ~n242 & ~n779 ;
  assign n781 = ~n776 & n780 ;
  assign n782 = n293 & n729 ;
  assign n783 = G8 & n782 ;
  assign n784 = ~G133 & ~n729 ;
  assign n785 = G8 & n784 ;
  assign n786 = n783 & n785 ;
  assign n787 = ~n783 & ~n785 ;
  assign n788 = ~n786 & ~n787 ;
  assign n789 = n220 & n729 ;
  assign n790 = n220 & ~n729 ;
  assign n791 = ~n789 & ~n790 ;
  assign n792 = G8 & ~n791 ;
  assign n793 = ~G142 & n729 ;
  assign n794 = ~G131 & ~n729 ;
  assign n795 = ~n793 & ~n794 ;
  assign n796 = G8 & ~n795 ;
  assign n797 = n792 & n796 ;
  assign n798 = ~n792 & ~n796 ;
  assign n799 = ~n797 & ~n798 ;
  assign n800 = n231 & n729 ;
  assign n801 = n231 & ~n729 ;
  assign n802 = ~n800 & ~n801 ;
  assign n803 = G8 & ~n802 ;
  assign n804 = ~G141 & n729 ;
  assign n805 = ~G130 & ~n729 ;
  assign n806 = ~n804 & ~n805 ;
  assign n807 = G8 & ~n806 ;
  assign n808 = n803 & n807 ;
  assign n809 = ~n803 & ~n807 ;
  assign n810 = ~n808 & ~n809 ;
  assign n811 = ~n799 & ~n810 ;
  assign n812 = ~n788 & n811 ;
  assign n813 = n781 & n812 ;
  assign n814 = ~n803 & n807 ;
  assign n815 = ~n776 & n814 ;
  assign n816 = ~n788 & ~n799 ;
  assign n817 = n815 & n816 ;
  assign n818 = ~n813 & ~n817 ;
  assign n819 = ~n792 & n796 ;
  assign n820 = ~n776 & ~n788 ;
  assign n821 = n819 & n820 ;
  assign n822 = ~n771 & n773 ;
  assign n823 = ~n788 & n822 ;
  assign n824 = ~n783 & n785 ;
  assign n825 = ~n823 & ~n824 ;
  assign n826 = ~n821 & n825 ;
  assign n827 = n818 & n826 ;
  assign n828 = ~n788 & ~n810 ;
  assign n829 = n242 & ~n779 ;
  assign n830 = ~n242 & n779 ;
  assign n831 = ~n829 & ~n830 ;
  assign n832 = ~n776 & ~n831 ;
  assign n833 = ~n799 & n832 ;
  assign n834 = n828 & n833 ;
  assign n835 = ~G136 & n729 ;
  assign n836 = ~G125 & ~n729 ;
  assign n837 = ~n835 & ~n836 ;
  assign n838 = n253 & ~n837 ;
  assign n839 = ~G139 & n729 ;
  assign n840 = ~G128 & ~n729 ;
  assign n841 = ~n839 & ~n840 ;
  assign n842 = n272 & ~n841 ;
  assign n843 = ~n272 & n841 ;
  assign n844 = ~n842 & ~n843 ;
  assign n845 = ~G138 & n729 ;
  assign n846 = ~G126 & ~n729 ;
  assign n847 = ~n845 & ~n846 ;
  assign n848 = ~n315 & ~n847 ;
  assign n849 = n315 & n847 ;
  assign n850 = ~n848 & ~n849 ;
  assign n851 = ~n844 & ~n850 ;
  assign n852 = n838 & n851 ;
  assign n853 = n315 & ~n847 ;
  assign n854 = ~n844 & n853 ;
  assign n855 = ~n272 & ~n841 ;
  assign n856 = ~n854 & ~n855 ;
  assign n857 = ~n852 & n856 ;
  assign n858 = n834 & ~n857 ;
  assign n859 = n827 & ~n858 ;
  assign n860 = ~n769 & n859 ;
  assign n861 = n740 & n742 ;
  assign n862 = ~n740 & ~n742 ;
  assign n863 = ~n861 & ~n862 ;
  assign n864 = ~n738 & ~n863 ;
  assign n865 = n759 & n864 ;
  assign n866 = n769 & ~n865 ;
  assign n867 = ~n859 & ~n866 ;
  assign n868 = ~n860 & ~n867 ;
  assign n869 = ~n388 & ~n446 ;
  assign n870 = ~n676 & ~n726 ;
  assign n871 = ~n414 & n870 ;
  assign n872 = n869 & n871 ;
  assign n873 = n170 & n872 ;
  assign G2551 = ~n158 ;
  assign G2552 = ~n159 ;
  assign G2553 = ~n160 ;
  assign G2554 = ~n167 ;
  assign G2555 = ~n167 ;
  assign G2556 = ~n170 ;
  assign G2557 = n181 ;
  assign G2531 = ~G115 ;
  assign G2532 = ~G115 ;
  assign G2533 = ~G115 ;
  assign G2534 = ~G124 ;
  assign G2535 = ~G124 ;
  assign G2536 = ~G137 ;
  assign G2537 = ~G137 ;
  assign G2538 = ~G137 ;
  assign G2539 = ~G32 ;
  assign G2540 = ~G106 ;
  assign G2541 = ~G64 ;
  assign G2542 = ~G76 ;
  assign G2543 = ~G53 ;
  assign G2544 = ~G96 ;
  assign G2545 = ~G43 ;
  assign G2546 = ~G86 ;
  assign G2547 = ~n184 ;
  assign G2548 = ~n186 ;
  assign G2549 = G115 ;
  assign G2550 = n187 ;
  assign G2558 = n198 ;
  assign G2559 = n209 ;
  assign G2560 = n220 ;
  assign G2561 = n231 ;
  assign G2562 = n242 ;
  assign G2563 = ~n255 ;
  assign G2564 = ~n258 ;
  assign G2565 = ~n261 ;
  assign G2566 = ~n272 ;
  assign G2567 = ~n242 ;
  assign G2568 = ~n231 ;
  assign G2569 = ~n220 ;
  assign G2570 = ~n282 ;
  assign G2571 = ~n293 ;
  assign G2572 = ~n304 ;
  assign G2573 = n318 ;
  assign G2574 = n318 ;
  assign G2575 = n321 ;
  assign G2576 = n321 ;
  assign G2577 = ~n325 ;
  assign G2578 = n328 ;
  assign G2579 = n328 ;
  assign G2580 = ~n355 ;
  assign G2581 = ~n388 ;
  assign G2582 = n414 ;
  assign G2583 = n446 ;
  assign G2584 = ~n609 ;
  assign G2585 = ~n609 ;
  assign G2586 = ~n632 ;
  assign G2587 = ~n676 ;
  assign G2588 = n708 ;
  assign G2589 = n708 ;
  assign G2590 = ~n726 ;
  assign G2591 = n868 ;
  assign G2592 = 1'b0 ;
  assign G2593 = ~n873 ;
  assign G2594 = ~n873 ;
endmodule
