module top(pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 , pi8 , pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 , pi16 , pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 , po0 , po1 , po2 , po3 , po4 , po5 , po6 , po7 , po8 , po9 , po10 , po11 , po12 , po13 , po14 , po15 , po16 , po17 , po18 , po19 , po20 , po21 , po22 , po23 , po24 );
  input pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 , pi8 , pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 , pi16 , pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 ;
  output po0 , po1 , po2 , po3 , po4 , po5 , po6 , po7 , po8 , po9 , po10 , po11 , po12 , po13 , po14 , po15 , po16 , po17 , po18 , po19 , po20 , po21 , po22 , po23 , po24 ;
  wire n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674;
  assign n25 = pi5 | pi8 ;
  assign n26 = pi7 | pi10 ;
  assign n27 = pi4 | pi6 ;
  assign n28 = n26 | n27 ;
  assign n29 = n25 | n28 ;
  assign n30 = pi1 | pi2 ;
  assign n31 = pi0 | n30 ;
  assign n32 = pi3 | n31 ;
  assign n33 = pi9 | n32 ;
  assign n34 = pi11 | pi12 ;
  assign n35 = n33 | n34 ;
  assign n36 = n29 | n35 ;
  assign n37 = pi13 | n36 ;
  assign n38 = pi14 | n37 ;
  assign n39 = pi15 | n38 ;
  assign n40 = pi16 | pi17 ;
  assign n41 = n39 | n40 ;
  assign n42 = pi18 | pi19 ;
  assign n43 = pi20 | n42 ;
  assign n44 = n41 | n43 ;
  assign n45 = ~pi22 & n44 ;
  assign n46 = pi21 | pi22 ;
  assign n47 = n44 & ~n46 ;
  assign n48 = ~pi21 & pi22 ;
  assign n49 = ( pi21 & n44 ) | ( pi21 & ~n48 ) | ( n44 & ~n48 );
  assign n50 = ( ~n45 & n47 ) | ( ~n45 & n49 ) | ( n47 & n49 );
  assign n51 = ~pi22 & n38 ;
  assign n52 = ~pi15 & n51 ;
  assign n53 = pi15 | n51 ;
  assign n54 = ( ~n51 & n52 ) | ( ~n51 & n53 ) | ( n52 & n53 );
  assign n55 = ( ~pi22 & n41 ) | ( ~pi22 & n42 ) | ( n41 & n42 );
  assign n56 = ( pi20 & pi22 ) | ( pi20 & n42 ) | ( pi22 & n42 );
  assign n57 = ( pi20 & n41 ) | ( pi20 & n56 ) | ( n41 & n56 );
  assign n58 = n55 & ~n57 ;
  assign n59 = ~pi22 & n57 ;
  assign n60 = ( pi20 & n58 ) | ( pi20 & ~n59 ) | ( n58 & ~n59 );
  assign n61 = n54 | n60 ;
  assign n62 = n50 | n61 ;
  assign n63 = pi18 & ~pi22 ;
  assign n64 = ( ~pi22 & n41 ) | ( ~pi22 & n63 ) | ( n41 & n63 );
  assign n65 = pi19 & n63 ;
  assign n66 = pi19 & ~pi22 ;
  assign n67 = ( n41 & n65 ) | ( n41 & n66 ) | ( n65 & n66 );
  assign n68 = pi19 & ~n67 ;
  assign n69 = ( n64 & ~n67 ) | ( n64 & n68 ) | ( ~n67 & n68 );
  assign n70 = ~pi22 & n41 ;
  assign n71 = pi18 | pi22 ;
  assign n72 = n41 & ~n71 ;
  assign n73 = ~pi18 & n71 ;
  assign n74 = ( pi18 & n41 ) | ( pi18 & ~n73 ) | ( n41 & ~n73 );
  assign n75 = ( ~n70 & n72 ) | ( ~n70 & n74 ) | ( n72 & n74 );
  assign n76 = n69 & n75 ;
  assign n77 = pi16 & ~pi22 ;
  assign n78 = ( ~pi22 & n39 ) | ( ~pi22 & n77 ) | ( n39 & n77 );
  assign n79 = pi17 & ~n78 ;
  assign n80 = ~pi17 & n78 ;
  assign n81 = n79 | n80 ;
  assign n82 = ~pi22 & n39 ;
  assign n83 = pi16 | pi22 ;
  assign n84 = n39 & ~n83 ;
  assign n85 = pi16 | n84 ;
  assign n86 = ( ~n82 & n84 ) | ( ~n82 & n85 ) | ( n84 & n85 );
  assign n87 = n81 & ~n86 ;
  assign n88 = n76 & n87 ;
  assign n89 = ~n62 & n88 ;
  assign n90 = n81 | n86 ;
  assign n91 = n76 & ~n90 ;
  assign n92 = ~n54 & n60 ;
  assign n93 = ~n50 & n92 ;
  assign n94 = n91 & n93 ;
  assign n95 = n69 & ~n75 ;
  assign n96 = ~n90 & n95 ;
  assign n97 = n93 & n96 ;
  assign n98 = ~n50 & n60 ;
  assign n99 = n54 & n98 ;
  assign n100 = ~n69 & n75 ;
  assign n101 = ~n90 & n100 ;
  assign n102 = n99 & n101 ;
  assign n103 = n54 & ~n60 ;
  assign n104 = n50 & n103 ;
  assign n105 = ~n81 & n86 ;
  assign n106 = n95 & n105 ;
  assign n107 = n104 & n106 ;
  assign n108 = n50 & n60 ;
  assign n109 = n54 & n108 ;
  assign n110 = n87 & n95 ;
  assign n111 = n109 & n110 ;
  assign n112 = n106 & n109 ;
  assign n113 = n88 & n99 ;
  assign n114 = n100 & n105 ;
  assign n115 = n93 & n114 ;
  assign n116 = n113 | n115 ;
  assign n117 = n112 | n116 ;
  assign n118 = ~n50 & n103 ;
  assign n119 = n87 & n100 ;
  assign n120 = n118 & n119 ;
  assign n121 = ~n54 & n108 ;
  assign n122 = n106 & n121 ;
  assign n123 = n119 & n121 ;
  assign n124 = n122 | n123 ;
  assign n125 = n120 | n124 ;
  assign n126 = n117 | n125 ;
  assign n127 = n76 & n105 ;
  assign n128 = n121 & n127 ;
  assign n129 = n110 & n121 ;
  assign n130 = n81 & n86 ;
  assign n131 = n95 & n130 ;
  assign n132 = n121 & n131 ;
  assign n133 = n129 | n132 ;
  assign n134 = n128 | n133 ;
  assign n135 = n100 & n130 ;
  assign n136 = n121 & n135 ;
  assign n137 = n88 & n109 ;
  assign n138 = n136 | n137 ;
  assign n139 = n134 | n138 ;
  assign n140 = n88 & n104 ;
  assign n141 = n88 & n93 ;
  assign n142 = n140 | n141 ;
  assign n143 = n109 & n135 ;
  assign n144 = n118 & n135 ;
  assign n145 = n143 | n144 ;
  assign n146 = n142 | n145 ;
  assign n147 = n139 | n146 ;
  assign n148 = n126 | n147 ;
  assign n149 = n104 & n119 ;
  assign n150 = n69 | n75 ;
  assign n151 = n87 & ~n150 ;
  assign n152 = n99 & n151 ;
  assign n153 = n114 & n121 ;
  assign n154 = n152 | n153 ;
  assign n155 = n149 | n154 ;
  assign n156 = n148 | n155 ;
  assign n157 = n93 & n127 ;
  assign n158 = n104 & n131 ;
  assign n159 = ~n62 & n131 ;
  assign n160 = n99 & n106 ;
  assign n161 = n90 | n150 ;
  assign n162 = n99 & ~n161 ;
  assign n163 = n50 & ~n61 ;
  assign n164 = n131 & n163 ;
  assign n165 = n91 & n109 ;
  assign n166 = n109 & n127 ;
  assign n167 = n101 & n163 ;
  assign n168 = n91 & n121 ;
  assign n169 = n167 | n168 ;
  assign n170 = n166 | n169 ;
  assign n171 = n165 | n170 ;
  assign n172 = n164 | n171 ;
  assign n173 = n162 | n172 ;
  assign n174 = n160 | n173 ;
  assign n175 = n159 | n174 ;
  assign n176 = n91 & n104 ;
  assign n177 = n130 & ~n150 ;
  assign n178 = n121 & n177 ;
  assign n179 = n176 | n178 ;
  assign n180 = n93 & n131 ;
  assign n181 = n105 & ~n150 ;
  assign n182 = n109 & n181 ;
  assign n183 = n76 & n130 ;
  assign n184 = n121 & n183 ;
  assign n185 = n182 | n184 ;
  assign n186 = n101 & n104 ;
  assign n187 = n104 & n110 ;
  assign n188 = n186 | n187 ;
  assign n189 = n185 | n188 ;
  assign n190 = n180 | n189 ;
  assign n191 = n179 | n190 ;
  assign n192 = n175 | n191 ;
  assign n193 = n158 | n192 ;
  assign n194 = n157 | n193 ;
  assign n195 = n163 & n181 ;
  assign n196 = n104 & n183 ;
  assign n197 = n195 | n196 ;
  assign n198 = n194 | n197 ;
  assign n199 = n156 | n198 ;
  assign n200 = n96 & n163 ;
  assign n201 = ~n62 & n181 ;
  assign n202 = n200 | n201 ;
  assign n203 = n88 & n121 ;
  assign n204 = n114 & n118 ;
  assign n205 = n99 & n183 ;
  assign n206 = ~n161 & n163 ;
  assign n207 = n109 & ~n161 ;
  assign n208 = n109 & n119 ;
  assign n209 = n109 & n114 ;
  assign n210 = n121 & n181 ;
  assign n211 = n99 & n177 ;
  assign n212 = n88 & n118 ;
  assign n213 = n211 | n212 ;
  assign n214 = n118 & n177 ;
  assign n215 = n118 & n151 ;
  assign n216 = n214 | n215 ;
  assign n217 = n213 | n216 ;
  assign n218 = n109 & n131 ;
  assign n219 = n96 & n109 ;
  assign n220 = n218 | n219 ;
  assign n221 = n104 & n127 ;
  assign n222 = n88 & n163 ;
  assign n223 = n221 | n222 ;
  assign n224 = n220 | n223 ;
  assign n225 = n106 & n118 ;
  assign n226 = n99 & n110 ;
  assign n227 = n225 | n226 ;
  assign n228 = n224 | n227 ;
  assign n229 = n217 | n228 ;
  assign n230 = n210 | n229 ;
  assign n231 = n209 | n230 ;
  assign n232 = n208 | n231 ;
  assign n233 = n91 & n163 ;
  assign n234 = n109 & n177 ;
  assign n235 = n233 | n234 ;
  assign n236 = n232 | n235 ;
  assign n237 = n101 & n118 ;
  assign n238 = n104 & n114 ;
  assign n239 = n93 & n110 ;
  assign n240 = n238 | n239 ;
  assign n241 = n237 | n240 ;
  assign n242 = n236 | n241 ;
  assign n243 = n207 | n242 ;
  assign n244 = n206 | n243 ;
  assign n245 = n205 | n244 ;
  assign n246 = n204 | n245 ;
  assign n247 = n203 | n246 ;
  assign n248 = n202 | n247 ;
  assign n249 = n199 | n248 ;
  assign n250 = n111 | n249 ;
  assign n251 = n107 | n250 ;
  assign n252 = n102 | n251 ;
  assign n253 = n97 | n252 ;
  assign n254 = n94 | n253 ;
  assign n255 = n89 | n254 ;
  assign n256 = pi2 & pi22 ;
  assign n257 = pi0 & ~pi22 ;
  assign n258 = ( ~pi22 & n30 ) | ( ~pi22 & n257 ) | ( n30 & n257 );
  assign n259 = pi0 | pi1 ;
  assign n260 = pi2 & n259 ;
  assign n261 = n258 & ~n260 ;
  assign n262 = n256 | n261 ;
  assign n263 = ~pi22 & n36 ;
  assign n264 = pi13 & ~n263 ;
  assign n265 = ~pi13 & n263 ;
  assign n266 = n264 | n265 ;
  assign n267 = n109 & n151 ;
  assign n268 = n109 & n183 ;
  assign n269 = n267 | n268 ;
  assign n270 = n111 | n179 ;
  assign n271 = n133 | n270 ;
  assign n272 = n127 & n163 ;
  assign n273 = n221 | n234 ;
  assign n274 = n272 | n273 ;
  assign n275 = n271 | n274 ;
  assign n276 = n96 & n104 ;
  assign n277 = n200 | n276 ;
  assign n278 = n143 | n277 ;
  assign n279 = n101 & n109 ;
  assign n280 = n136 | n208 ;
  assign n281 = n106 & n163 ;
  assign n282 = n101 & n121 ;
  assign n283 = n281 | n282 ;
  assign n284 = n280 | n283 ;
  assign n285 = n279 | n284 ;
  assign n286 = n278 | n285 ;
  assign n287 = n107 | n286 ;
  assign n288 = n121 & ~n161 ;
  assign n289 = n196 | n288 ;
  assign n290 = n233 | n289 ;
  assign n291 = n287 | n290 ;
  assign n292 = n275 | n291 ;
  assign n293 = n128 | n210 ;
  assign n294 = n166 | n203 ;
  assign n295 = n293 | n294 ;
  assign n296 = n207 | n295 ;
  assign n297 = n168 | n218 ;
  assign n298 = n163 & n183 ;
  assign n299 = n165 | n298 ;
  assign n300 = n297 | n299 ;
  assign n301 = n140 | n222 ;
  assign n302 = n300 | n301 ;
  assign n303 = n137 | n302 ;
  assign n304 = n182 | n303 ;
  assign n305 = n110 & n163 ;
  assign n306 = n187 | n305 ;
  assign n307 = n104 & n135 ;
  assign n308 = n209 | n307 ;
  assign n309 = n135 & n163 ;
  assign n310 = n149 | n309 ;
  assign n311 = n96 & n121 ;
  assign n312 = n164 | n311 ;
  assign n313 = n310 | n312 ;
  assign n314 = n308 | n313 ;
  assign n315 = n124 | n314 ;
  assign n316 = n153 | n315 ;
  assign n317 = n219 | n316 ;
  assign n318 = n306 | n317 ;
  assign n319 = n158 | n318 ;
  assign n320 = n112 | n319 ;
  assign n321 = n304 | n320 ;
  assign n322 = n121 & n151 ;
  assign n323 = n184 | n322 ;
  assign n324 = n321 | n323 ;
  assign n325 = n296 | n324 ;
  assign n326 = n292 | n325 ;
  assign n327 = n269 | n326 ;
  assign n328 = n266 & n327 ;
  assign n329 = ~pi22 & n37 ;
  assign n330 = ~pi14 & n329 ;
  assign n331 = pi14 & ~n329 ;
  assign n332 = n330 | n331 ;
  assign n333 = ~n62 & n106 ;
  assign n334 = ~n62 & n110 ;
  assign n335 = n104 & ~n161 ;
  assign n336 = n99 & n131 ;
  assign n337 = n180 | n336 ;
  assign n338 = n91 & n99 ;
  assign n339 = n99 & n127 ;
  assign n340 = n338 | n339 ;
  assign n341 = n157 | n340 ;
  assign n342 = n113 | n341 ;
  assign n343 = n337 | n342 ;
  assign n344 = n163 & n177 ;
  assign n345 = n195 | n344 ;
  assign n346 = n226 | n345 ;
  assign n347 = n205 | n346 ;
  assign n348 = n141 | n347 ;
  assign n349 = n104 & n151 ;
  assign n350 = n104 & n181 ;
  assign n351 = n349 | n350 ;
  assign n352 = n93 & n183 ;
  assign n353 = n119 & n163 ;
  assign n354 = n352 | n353 ;
  assign n355 = n151 & n163 ;
  assign n356 = n104 & n177 ;
  assign n357 = n355 | n356 ;
  assign n358 = n354 | n357 ;
  assign n359 = n351 | n358 ;
  assign n360 = n348 | n359 ;
  assign n361 = n343 | n360 ;
  assign n362 = n206 | n361 ;
  assign n363 = n335 | n362 ;
  assign n364 = n94 | n363 ;
  assign n365 = n96 & n118 ;
  assign n366 = n110 & n118 ;
  assign n367 = ~n62 & n183 ;
  assign n368 = n93 & ~n161 ;
  assign n369 = n212 | n368 ;
  assign n370 = n91 & n118 ;
  assign n371 = n118 & n127 ;
  assign n372 = n370 | n371 ;
  assign n373 = n186 | n238 ;
  assign n374 = n162 | n373 ;
  assign n375 = n372 | n374 ;
  assign n376 = n114 & n163 ;
  assign n377 = n167 | n376 ;
  assign n378 = n89 | n377 ;
  assign n379 = n375 | n378 ;
  assign n380 = n369 | n379 ;
  assign n381 = n367 | n380 ;
  assign n382 = n118 & n183 ;
  assign n383 = ~n62 & n127 ;
  assign n384 = n382 | n383 ;
  assign n385 = n381 | n384 ;
  assign n386 = n118 & n131 ;
  assign n387 = ~n62 & n91 ;
  assign n388 = n159 | n387 ;
  assign n389 = n386 | n388 ;
  assign n390 = n385 | n389 ;
  assign n391 = n366 | n390 ;
  assign n392 = n365 | n391 ;
  assign n393 = n364 | n392 ;
  assign n394 = n334 | n393 ;
  assign n395 = n333 | n394 ;
  assign n396 = n225 | n395 ;
  assign n397 = n99 & n181 ;
  assign n398 = n93 & n181 ;
  assign n399 = n102 | n398 ;
  assign n400 = n397 | n399 ;
  assign n401 = n93 & n151 ;
  assign n402 = n93 & n177 ;
  assign n403 = n401 | n402 ;
  assign n404 = n400 | n403 ;
  assign n405 = n93 & n101 ;
  assign n406 = n211 | n405 ;
  assign n407 = n152 | n406 ;
  assign n408 = n404 | n407 ;
  assign n409 = n93 & n106 ;
  assign n410 = n96 & n99 ;
  assign n411 = n99 & n119 ;
  assign n412 = n93 & n119 ;
  assign n413 = n93 & n135 ;
  assign n414 = n99 & n114 ;
  assign n415 = n413 | n414 ;
  assign n416 = n412 | n415 ;
  assign n417 = n99 & n135 ;
  assign n418 = n239 | n417 ;
  assign n419 = n416 | n418 ;
  assign n420 = n411 | n419 ;
  assign n421 = n410 | n420 ;
  assign n422 = n97 | n160 ;
  assign n423 = n421 | n422 ;
  assign n424 = n409 | n423 ;
  assign n425 = n364 | n424 ;
  assign n426 = n373 | n425 ;
  assign n427 = n377 | n426 ;
  assign n428 = n408 | n427 ;
  assign n429 = n115 | n428 ;
  assign n430 = n396 & n429 ;
  assign n431 = n327 & ~n430 ;
  assign n432 = n332 | n431 ;
  assign n433 = ~n396 & n429 ;
  assign n434 = n396 & ~n429 ;
  assign n435 = n433 | n434 ;
  assign n436 = ~n431 & n435 ;
  assign n437 = n396 | n429 ;
  assign n438 = ~n327 & n437 ;
  assign n439 = n435 | n438 ;
  assign n440 = n332 & ~n439 ;
  assign n441 = n436 | n440 ;
  assign n442 = n432 & ~n441 ;
  assign n443 = ~n328 & n442 ;
  assign n444 = pi8 | pi10 ;
  assign n445 = pi4 | pi5 ;
  assign n446 = n444 | n445 ;
  assign n447 = pi6 | pi7 ;
  assign n448 = n33 | n447 ;
  assign n449 = n446 | n448 ;
  assign n450 = ~pi22 & n449 ;
  assign n451 = pi11 & ~n450 ;
  assign n452 = ~pi11 & n450 ;
  assign n453 = n451 | n452 ;
  assign n454 = n327 & n453 ;
  assign n455 = ~n62 & n96 ;
  assign n456 = n187 | n222 ;
  assign n457 = n455 | n456 ;
  assign n458 = n238 | n457 ;
  assign n459 = n239 | n458 ;
  assign n460 = n158 | n208 ;
  assign n461 = n186 | n460 ;
  assign n462 = n311 | n461 ;
  assign n463 = n356 | n462 ;
  assign n464 = n205 | n463 ;
  assign n465 = n387 | n464 ;
  assign n466 = n102 | n184 ;
  assign n467 = n97 | n466 ;
  assign n468 = n409 | n467 ;
  assign n469 = n366 | n468 ;
  assign n470 = n233 | n344 ;
  assign n471 = n376 | n470 ;
  assign n472 = n339 | n471 ;
  assign n473 = n148 | n219 ;
  assign n474 = n405 | n473 ;
  assign n475 = ~n62 & n177 ;
  assign n476 = n176 | n475 ;
  assign n477 = n474 | n476 ;
  assign n478 = n352 | n410 ;
  assign n479 = n368 | n478 ;
  assign n480 = n477 | n479 ;
  assign n481 = n472 | n480 ;
  assign n482 = n469 | n481 ;
  assign n483 = n465 | n482 ;
  assign n484 = n459 | n483 ;
  assign n485 = ~n62 & n135 ;
  assign n486 = ~n62 & n151 ;
  assign n487 = ~n62 & n119 ;
  assign n488 = n215 | n487 ;
  assign n489 = n153 | n209 ;
  assign n490 = n488 | n489 ;
  assign n491 = n367 | n490 ;
  assign n492 = n211 | n382 ;
  assign n493 = n214 | n492 ;
  assign n494 = n111 | n268 ;
  assign n495 = n218 | n494 ;
  assign n496 = n493 | n495 ;
  assign n497 = n221 | n272 ;
  assign n498 = n386 | n497 ;
  assign n499 = n496 | n498 ;
  assign n500 = n491 | n499 ;
  assign n501 = n175 | n500 ;
  assign n502 = n486 | n501 ;
  assign n503 = n203 | n353 ;
  assign n504 = n502 | n503 ;
  assign n505 = n485 | n504 ;
  assign n506 = n484 | n505 ;
  assign n507 = n206 | n383 ;
  assign n508 = n128 | n197 ;
  assign n509 = n382 | n508 ;
  assign n510 = n111 | n322 ;
  assign n511 = n355 | n510 ;
  assign n512 = n120 | n511 ;
  assign n513 = n209 | n512 ;
  assign n514 = n509 | n513 ;
  assign n515 = n234 | n514 ;
  assign n516 = n350 | n515 ;
  assign n517 = n136 | n219 ;
  assign n518 = n371 | n517 ;
  assign n519 = n169 | n518 ;
  assign n520 = n516 | n519 ;
  assign n521 = n507 | n520 ;
  assign n522 = n166 | n409 ;
  assign n523 = n288 | n298 ;
  assign n524 = n522 | n523 ;
  assign n525 = n184 | n524 ;
  assign n526 = n165 | n349 ;
  assign n527 = n525 | n526 ;
  assign n528 = n411 | n527 ;
  assign n529 = n89 | n237 ;
  assign n530 = n124 | n529 ;
  assign n531 = n112 | n208 ;
  assign n532 = n530 | n531 ;
  assign n533 = n162 | n410 ;
  assign n534 = n412 | n533 ;
  assign n535 = n532 | n534 ;
  assign n536 = n487 | n535 ;
  assign n537 = ~n62 & n114 ;
  assign n538 = n369 | n376 ;
  assign n539 = n267 | n279 ;
  assign n540 = n218 | n539 ;
  assign n541 = n538 | n540 ;
  assign n542 = n144 | n541 ;
  assign n543 = n353 | n542 ;
  assign n544 = n137 | n182 ;
  assign n545 = n133 | n544 ;
  assign n546 = n418 | n545 ;
  assign n547 = n543 | n546 ;
  assign n548 = n282 | n547 ;
  assign n549 = n178 | n548 ;
  assign n550 = n203 | n549 ;
  assign n551 = n238 | n550 ;
  assign n552 = n413 | n551 ;
  assign n553 = n537 | n552 ;
  assign n554 = n268 | n455 ;
  assign n555 = n553 | n554 ;
  assign n556 = n153 | n207 ;
  assign n557 = n143 | n160 ;
  assign n558 = n556 | n557 ;
  assign n559 = n555 | n558 ;
  assign n560 = n344 | n370 ;
  assign n561 = n210 | n311 ;
  assign n562 = n97 | n561 ;
  assign n563 = n560 | n562 ;
  assign n564 = n559 | n563 ;
  assign n565 = n536 | n564 ;
  assign n566 = n186 | n335 ;
  assign n567 = ~n62 & n101 ;
  assign n568 = n204 | n567 ;
  assign n569 = n566 | n568 ;
  assign n570 = n565 | n569 ;
  assign n571 = n528 | n570 ;
  assign n572 = n521 | n571 ;
  assign n573 = n356 | n414 ;
  assign n574 = n485 | n573 ;
  assign n575 = n367 | n574 ;
  assign n576 = n572 | n575 ;
  assign n577 = n506 & n576 ;
  assign n578 = n396 & ~n577 ;
  assign n579 = n454 & ~n578 ;
  assign n580 = ~n454 & n578 ;
  assign n581 = n579 | n580 ;
  assign n582 = pi11 & ~pi22 ;
  assign n583 = n450 | n582 ;
  assign n584 = pi12 & n583 ;
  assign n585 = pi12 | n582 ;
  assign n586 = n450 | n585 ;
  assign n587 = ~n584 & n586 ;
  assign n588 = n327 & n587 ;
  assign n589 = ~n581 & n588 ;
  assign n590 = n579 | n589 ;
  assign n591 = n328 & ~n442 ;
  assign n592 = n443 | n591 ;
  assign n593 = n590 & ~n592 ;
  assign n594 = n443 | n593 ;
  assign n595 = n506 | n576 ;
  assign n596 = ~n396 & n595 ;
  assign n597 = ~n506 & n576 ;
  assign n598 = n506 & ~n576 ;
  assign n599 = n597 | n598 ;
  assign n600 = n596 | n599 ;
  assign n601 = n332 & ~n600 ;
  assign n602 = n578 | n599 ;
  assign n603 = n332 & ~n602 ;
  assign n604 = ( n578 & ~n601 ) | ( n578 & n603 ) | ( ~n601 & n603 );
  assign n605 = ~n454 & n604 ;
  assign n606 = n454 & ~n604 ;
  assign n607 = n605 | n606 ;
  assign n608 = n431 | n435 ;
  assign n609 = n587 | n608 ;
  assign n610 = ~n439 & n586 ;
  assign n611 = ~n584 & n610 ;
  assign n612 = n609 & ~n611 ;
  assign n613 = n435 & ~n438 ;
  assign n614 = n266 & n613 ;
  assign n615 = ~n266 & n436 ;
  assign n616 = n614 | n615 ;
  assign n617 = n612 & ~n616 ;
  assign n618 = ~n607 & n617 ;
  assign n619 = n605 | n618 ;
  assign n620 = n332 & n613 ;
  assign n621 = ~n331 & n436 ;
  assign n622 = ~n330 & n621 ;
  assign n623 = n266 & ~n439 ;
  assign n624 = n266 | n608 ;
  assign n625 = ~n623 & n624 ;
  assign n626 = ~n622 & n625 ;
  assign n627 = ~n620 & n626 ;
  assign n628 = n619 & n627 ;
  assign n629 = n619 | n627 ;
  assign n630 = ~n628 & n629 ;
  assign n631 = n581 & ~n588 ;
  assign n632 = n589 | n631 ;
  assign n633 = n630 & ~n632 ;
  assign n634 = n628 | n633 ;
  assign n635 = ~n590 & n592 ;
  assign n636 = n593 | n635 ;
  assign n637 = n634 & ~n636 ;
  assign n638 = n122 | n338 ;
  assign n639 = n417 | n638 ;
  assign n640 = n107 | n158 ;
  assign n641 = n118 & n181 ;
  assign n642 = n239 | n641 ;
  assign n643 = n640 | n642 ;
  assign n644 = n374 | n643 ;
  assign n645 = n89 | n644 ;
  assign n646 = n212 | n645 ;
  assign n647 = n639 | n646 ;
  assign n648 = n409 | n412 ;
  assign n649 = n311 | n397 ;
  assign n650 = n648 | n649 ;
  assign n651 = n455 | n650 ;
  assign n652 = n152 | n215 ;
  assign n653 = n651 | n652 ;
  assign n654 = n647 | n653 ;
  assign n655 = n222 | n654 ;
  assign n656 = n221 | n349 ;
  assign n657 = n195 | n656 ;
  assign n658 = n655 | n657 ;
  assign n659 = n210 | n288 ;
  assign n660 = n234 | n659 ;
  assign n661 = n405 | n660 ;
  assign n662 = n157 | n661 ;
  assign n663 = n334 | n662 ;
  assign n664 = n118 & ~n161 ;
  assign n665 = n663 | n664 ;
  assign n666 = n387 | n665 ;
  assign n667 = n282 | n666 ;
  assign n668 = n205 | n383 ;
  assign n669 = n333 | n668 ;
  assign n670 = n115 | n410 ;
  assign n671 = n200 | n305 ;
  assign n672 = n670 | n671 ;
  assign n673 = n669 | n672 ;
  assign n674 = n485 | n673 ;
  assign n675 = n667 | n674 ;
  assign n676 = n204 | n237 ;
  assign n677 = n167 | n676 ;
  assign n678 = n178 | n677 ;
  assign n679 = n233 | n353 ;
  assign n680 = n517 | n679 ;
  assign n681 = n120 | n680 ;
  assign n682 = n678 | n681 ;
  assign n683 = n675 | n682 ;
  assign n684 = n207 | n279 ;
  assign n685 = n411 | n684 ;
  assign n686 = n143 | n307 ;
  assign n687 = n336 | n402 ;
  assign n688 = n686 | n687 ;
  assign n689 = n159 | n382 ;
  assign n690 = n688 | n689 ;
  assign n691 = n685 | n690 ;
  assign n692 = n142 | n691 ;
  assign n693 = n683 | n692 ;
  assign n694 = n658 | n693 ;
  assign n695 = n214 | n694 ;
  assign n696 = n166 | n387 ;
  assign n697 = n94 | n696 ;
  assign n698 = n112 | n168 ;
  assign n699 = n205 | n698 ;
  assign n700 = n697 | n699 ;
  assign n701 = n511 | n700 ;
  assign n702 = n160 | n176 ;
  assign n703 = n225 | n352 ;
  assign n704 = n702 | n703 ;
  assign n705 = n234 | n704 ;
  assign n706 = n701 | n705 ;
  assign n707 = n272 | n305 ;
  assign n708 = n140 | n707 ;
  assign n709 = n402 | n708 ;
  assign n710 = n89 | n709 ;
  assign n711 = n706 | n710 ;
  assign n712 = n157 | n222 ;
  assign n713 = n214 | n712 ;
  assign n714 = n371 | n713 ;
  assign n715 = n128 | n276 ;
  assign n716 = n116 | n334 ;
  assign n717 = n204 | n349 ;
  assign n718 = n350 | n475 ;
  assign n719 = n201 | n718 ;
  assign n720 = n717 | n719 ;
  assign n721 = n716 | n720 ;
  assign n722 = n152 | n721 ;
  assign n723 = n338 | n722 ;
  assign n724 = n555 | n723 ;
  assign n725 = n715 | n724 ;
  assign n726 = n107 | n165 ;
  assign n727 = n221 | n281 ;
  assign n728 = n726 | n727 ;
  assign n729 = n725 | n728 ;
  assign n730 = n714 | n729 ;
  assign n731 = n162 | n730 ;
  assign n732 = n711 | n731 ;
  assign n733 = n401 | n466 ;
  assign n734 = n641 | n733 ;
  assign n735 = n386 | n734 ;
  assign n736 = n732 | n735 ;
  assign n737 = n695 & n736 ;
  assign n738 = n506 & ~n737 ;
  assign n739 = pi4 | n32 ;
  assign n740 = pi5 | n739 ;
  assign n741 = n447 | n740 ;
  assign n742 = pi8 | n741 ;
  assign n743 = ~pi22 & n742 ;
  assign n744 = pi9 & ~n743 ;
  assign n745 = ~pi9 & n743 ;
  assign n746 = n744 | n745 ;
  assign n747 = n327 & n746 ;
  assign n748 = ~n738 & n747 ;
  assign n749 = n738 & ~n747 ;
  assign n750 = n748 | n749 ;
  assign n751 = pi9 | n742 ;
  assign n752 = ~pi22 & n751 ;
  assign n753 = ~pi10 & n752 ;
  assign n754 = pi10 & ~n752 ;
  assign n755 = n753 | n754 ;
  assign n756 = n327 & n755 ;
  assign n757 = ~n750 & n756 ;
  assign n758 = n748 | n757 ;
  assign n759 = ~n578 & n599 ;
  assign n760 = ~n332 & n759 ;
  assign n761 = ( n266 & n602 ) | ( n266 & ~n760 ) | ( n602 & ~n760 );
  assign n762 = ( n266 & ~n600 ) | ( n266 & n760 ) | ( ~n600 & n760 );
  assign n763 = n761 & ~n762 ;
  assign n764 = n436 & ~n587 ;
  assign n765 = n453 | n608 ;
  assign n766 = n587 & n613 ;
  assign n767 = ~n439 & n453 ;
  assign n768 = n766 | n767 ;
  assign n769 = n765 & ~n768 ;
  assign n770 = ~n764 & n769 ;
  assign n771 = ~n596 & n599 ;
  assign n772 = ~n332 & n770 ;
  assign n773 = ( n770 & ~n771 ) | ( n770 & n772 ) | ( ~n771 & n772 );
  assign n774 = n763 & n773 ;
  assign n775 = n695 | n736 ;
  assign n776 = ~n506 & n775 ;
  assign n777 = ~n695 & n736 ;
  assign n778 = n695 & ~n736 ;
  assign n779 = n777 | n778 ;
  assign n780 = n776 | n779 ;
  assign n781 = n332 & ~n780 ;
  assign n782 = n738 | n779 ;
  assign n783 = n332 & ~n782 ;
  assign n784 = ( n738 & ~n781 ) | ( n738 & n783 ) | ( ~n781 & n783 );
  assign n785 = ~n747 & n784 ;
  assign n786 = n266 & n771 ;
  assign n787 = ~n266 & n759 ;
  assign n788 = ( n587 & n602 ) | ( n587 & ~n787 ) | ( n602 & ~n787 );
  assign n789 = ( n587 & ~n600 ) | ( n587 & n787 ) | ( ~n600 & n787 );
  assign n790 = n788 & ~n789 ;
  assign n791 = ~n786 & n790 ;
  assign n792 = n747 & ~n784 ;
  assign n793 = n785 | n792 ;
  assign n794 = n791 & ~n793 ;
  assign n795 = n785 | n794 ;
  assign n796 = n332 & ~n770 ;
  assign n797 = n771 & n796 ;
  assign n798 = ( n763 & n770 ) | ( n763 & ~n797 ) | ( n770 & ~n797 );
  assign n799 = ~n774 & n798 ;
  assign n800 = n795 & n799 ;
  assign n801 = n774 | n800 ;
  assign n802 = n758 & n801 ;
  assign n803 = n607 & ~n617 ;
  assign n804 = n618 | n803 ;
  assign n805 = n758 | n801 ;
  assign n806 = ~n802 & n805 ;
  assign n807 = ~n804 & n806 ;
  assign n808 = n802 | n807 ;
  assign n809 = ~n630 & n632 ;
  assign n810 = n633 | n809 ;
  assign n811 = n808 & ~n810 ;
  assign n812 = ~n808 & n810 ;
  assign n813 = n811 | n812 ;
  assign n814 = n804 & ~n806 ;
  assign n815 = n807 | n814 ;
  assign n816 = n453 & n613 ;
  assign n817 = n436 & ~n453 ;
  assign n818 = n608 | n755 ;
  assign n819 = ~n439 & n755 ;
  assign n820 = n818 & ~n819 ;
  assign n821 = ~n817 & n820 ;
  assign n822 = ~n816 & n821 ;
  assign n823 = ~pi22 & n740 ;
  assign n824 = pi6 & ~pi22 ;
  assign n825 = n823 | n824 ;
  assign n826 = ~pi7 & n825 ;
  assign n827 = pi7 & ~n825 ;
  assign n828 = n826 | n827 ;
  assign n829 = n327 & n828 ;
  assign n830 = n203 | n267 ;
  assign n831 = n149 | n830 ;
  assign n832 = n97 | n402 ;
  assign n833 = n831 | n832 ;
  assign n834 = n298 | n308 ;
  assign n835 = n833 | n834 ;
  assign n836 = n205 | n835 ;
  assign n837 = n94 | n411 ;
  assign n838 = n164 | n387 ;
  assign n839 = n210 | n305 ;
  assign n840 = n838 | n839 ;
  assign n841 = n664 | n840 ;
  assign n842 = n837 | n841 ;
  assign n843 = n836 | n842 ;
  assign n844 = n128 | n141 ;
  assign n845 = n157 | n335 ;
  assign n846 = n844 | n845 ;
  assign n847 = n485 | n846 ;
  assign n848 = n215 | n386 ;
  assign n849 = n847 | n848 ;
  assign n850 = n843 | n849 ;
  assign n851 = n132 | n850 ;
  assign n852 = n176 | n184 ;
  assign n853 = n851 | n852 ;
  assign n854 = n397 | n417 ;
  assign n855 = n144 | n854 ;
  assign n856 = n853 | n855 ;
  assign n857 = n122 | n309 ;
  assign n858 = n522 | n857 ;
  assign n859 = n493 | n858 ;
  assign n860 = n111 | n278 ;
  assign n861 = n239 | n860 ;
  assign n862 = n367 | n475 ;
  assign n863 = n861 | n862 ;
  assign n864 = n859 | n863 ;
  assign n865 = n355 | n365 ;
  assign n866 = n352 | n865 ;
  assign n867 = n333 | n866 ;
  assign n868 = n864 | n867 ;
  assign n869 = n234 | n868 ;
  assign n870 = n281 | n869 ;
  assign n871 = n167 | n207 ;
  assign n872 = n187 | n233 ;
  assign n873 = n871 | n872 ;
  assign n874 = n140 | n641 ;
  assign n875 = n370 | n874 ;
  assign n876 = n873 | n875 ;
  assign n877 = n62 | n161 ;
  assign n878 = ~n107 & n877 ;
  assign n879 = n399 | n461 ;
  assign n880 = n137 | n455 ;
  assign n881 = n279 | n880 ;
  assign n882 = n879 | n881 ;
  assign n883 = n180 | n268 ;
  assign n884 = n212 | n883 ;
  assign n885 = n882 | n884 ;
  assign n886 = n878 & ~n885 ;
  assign n887 = ~n876 & n886 ;
  assign n888 = ~n115 & n887 ;
  assign n889 = ~n870 & n888 ;
  assign n890 = ~n349 & n889 ;
  assign n891 = ~n856 & n890 ;
  assign n892 = n196 | n201 ;
  assign n893 = n486 | n892 ;
  assign n894 = n891 & ~n893 ;
  assign n895 = n233 | n305 ;
  assign n896 = n211 | n895 ;
  assign n897 = n160 | n356 ;
  assign n898 = n336 | n897 ;
  assign n899 = n137 | n898 ;
  assign n900 = n896 | n899 ;
  assign n901 = n405 | n413 ;
  assign n902 = n180 | n411 ;
  assign n903 = n164 | n902 ;
  assign n904 = n186 | n903 ;
  assign n905 = n159 | n904 ;
  assign n906 = n168 | n203 ;
  assign n907 = n184 | n906 ;
  assign n908 = n339 | n907 ;
  assign n909 = n197 | n908 ;
  assign n910 = n210 | n282 ;
  assign n911 = n268 | n910 ;
  assign n912 = n219 | n272 ;
  assign n913 = n911 | n912 ;
  assign n914 = n867 | n913 ;
  assign n915 = n909 | n914 ;
  assign n916 = n166 | n322 ;
  assign n917 = n208 | n916 ;
  assign n918 = n915 | n917 ;
  assign n919 = n162 | n225 ;
  assign n920 = n712 | n919 ;
  assign n921 = n165 | n311 ;
  assign n922 = n455 | n485 ;
  assign n923 = n921 | n922 ;
  assign n924 = n920 | n923 ;
  assign n925 = n918 | n924 ;
  assign n926 = n905 | n925 ;
  assign n927 = n124 | n926 ;
  assign n928 = n140 | n200 ;
  assign n929 = n334 | n928 ;
  assign n930 = n366 | n382 ;
  assign n931 = n929 | n930 ;
  assign n932 = n128 | n931 ;
  assign n933 = n309 | n932 ;
  assign n934 = n335 | n933 ;
  assign n935 = n402 | n934 ;
  assign n936 = n927 | n935 ;
  assign n937 = n901 | n936 ;
  assign n938 = n543 | n937 ;
  assign n939 = n900 | n938 ;
  assign n940 = n281 | n409 ;
  assign n941 = n367 | n940 ;
  assign n942 = n939 | n941 ;
  assign n943 = ~n894 & n942 ;
  assign n944 = n695 & ~n943 ;
  assign n945 = n829 & ~n944 ;
  assign n946 = ~pi22 & n741 ;
  assign n947 = ~pi8 & n946 ;
  assign n948 = pi8 & ~n946 ;
  assign n949 = n947 | n948 ;
  assign n950 = ~n829 & n944 ;
  assign n951 = n945 | n950 ;
  assign n952 = n949 & ~n951 ;
  assign n953 = n327 & n952 ;
  assign n954 = n945 | n953 ;
  assign n955 = n822 & n954 ;
  assign n956 = n822 & ~n955 ;
  assign n957 = n954 & ~n955 ;
  assign n958 = n956 | n957 ;
  assign n959 = n613 & n755 ;
  assign n960 = n436 & ~n755 ;
  assign n961 = n608 | n746 ;
  assign n962 = ~n439 & n746 ;
  assign n963 = n961 & ~n962 ;
  assign n964 = ~n960 & n963 ;
  assign n965 = ~n959 & n964 ;
  assign n966 = ~n776 & n779 ;
  assign n967 = n332 & n966 ;
  assign n968 = ~n738 & n779 ;
  assign n969 = ~n332 & n968 ;
  assign n970 = ( n266 & n782 ) | ( n266 & ~n969 ) | ( n782 & ~n969 );
  assign n971 = ( n266 & ~n780 ) | ( n266 & n969 ) | ( ~n780 & n969 );
  assign n972 = n970 & ~n971 ;
  assign n973 = ~n967 & n972 ;
  assign n974 = n587 & n771 ;
  assign n975 = ~n587 & n759 ;
  assign n976 = ( n453 & n602 ) | ( n453 & ~n975 ) | ( n602 & ~n975 );
  assign n977 = ( n453 & ~n600 ) | ( n453 & n975 ) | ( ~n600 & n975 );
  assign n978 = n976 & ~n977 ;
  assign n979 = ~n974 & n978 ;
  assign n980 = ( n965 & n973 ) | ( n965 & n979 ) | ( n973 & n979 );
  assign n981 = n958 & n980 ;
  assign n982 = n955 | n981 ;
  assign n983 = n750 & ~n756 ;
  assign n984 = n757 | n983 ;
  assign n985 = n982 & ~n984 ;
  assign n986 = n795 | n799 ;
  assign n987 = ~n800 & n986 ;
  assign n988 = ~n982 & n984 ;
  assign n989 = n985 | n988 ;
  assign n990 = ~n985 & n989 ;
  assign n991 = ( n985 & n987 ) | ( n985 & ~n990 ) | ( n987 & ~n990 );
  assign n992 = ~n815 & n991 ;
  assign n993 = n815 & ~n991 ;
  assign n994 = n992 | n993 ;
  assign n995 = n958 & ~n981 ;
  assign n996 = n613 & n746 ;
  assign n997 = n436 & ~n746 ;
  assign n998 = ( n608 & n949 ) | ( n608 & ~n997 ) | ( n949 & ~n997 );
  assign n999 = ( ~n439 & n949 ) | ( ~n439 & n997 ) | ( n949 & n997 );
  assign n1000 = n998 & ~n999 ;
  assign n1001 = ~n996 & n1000 ;
  assign n1002 = n453 & n771 ;
  assign n1003 = ~n453 & n759 ;
  assign n1004 = ( n602 & n755 ) | ( n602 & ~n1003 ) | ( n755 & ~n1003 );
  assign n1005 = ( ~n600 & n755 ) | ( ~n600 & n1003 ) | ( n755 & n1003 );
  assign n1006 = n1004 & ~n1005 ;
  assign n1007 = ~n1002 & n1006 ;
  assign n1008 = n1001 & n1007 ;
  assign n1009 = n166 | n365 ;
  assign n1010 = n357 | n1009 ;
  assign n1011 = n207 | n233 ;
  assign n1012 = n417 | n1011 ;
  assign n1013 = n1010 | n1012 ;
  assign n1014 = n401 | n664 ;
  assign n1015 = n1013 | n1014 ;
  assign n1016 = n102 | n212 ;
  assign n1017 = n306 | n1016 ;
  assign n1018 = n226 | n337 ;
  assign n1019 = n1017 | n1018 ;
  assign n1020 = n225 | n567 ;
  assign n1021 = n123 | n276 ;
  assign n1022 = n1020 | n1021 ;
  assign n1023 = n539 | n1022 ;
  assign n1024 = n367 | n1023 ;
  assign n1025 = n878 & ~n1024 ;
  assign n1026 = ~n490 & n1025 ;
  assign n1027 = ~n1019 & n1026 ;
  assign n1028 = ~n1015 & n1027 ;
  assign n1029 = n338 | n410 ;
  assign n1030 = n169 | n717 ;
  assign n1031 = n837 | n1030 ;
  assign n1032 = n186 | n281 ;
  assign n1033 = n143 | n1032 ;
  assign n1034 = n1031 | n1033 ;
  assign n1035 = n1029 | n1034 ;
  assign n1036 = n386 | n1035 ;
  assign n1037 = n165 | n344 ;
  assign n1038 = n383 | n1037 ;
  assign n1039 = n409 | n1038 ;
  assign n1040 = n353 | n397 ;
  assign n1041 = n398 | n1040 ;
  assign n1042 = n1039 | n1041 ;
  assign n1043 = n222 | n335 ;
  assign n1044 = n486 | n1043 ;
  assign n1045 = n1042 | n1044 ;
  assign n1046 = n913 | n1045 ;
  assign n1047 = n116 | n1046 ;
  assign n1048 = n184 | n1047 ;
  assign n1049 = n205 | n309 ;
  assign n1050 = n1048 | n1049 ;
  assign n1051 = n366 | n1050 ;
  assign n1052 = n1036 | n1051 ;
  assign n1053 = n178 | n1052 ;
  assign n1054 = n1028 & ~n1053 ;
  assign n1055 = ~n140 & n1054 ;
  assign n1056 = ~n152 & n1055 ;
  assign n1057 = ~n157 & n1056 ;
  assign n1058 = ~n485 & n1057 ;
  assign n1059 = n523 | n838 ;
  assign n1060 = n182 | n207 ;
  assign n1061 = n353 | n1060 ;
  assign n1062 = n1059 | n1061 ;
  assign n1063 = n281 | n485 ;
  assign n1064 = n641 | n1063 ;
  assign n1065 = n1062 | n1064 ;
  assign n1066 = n386 | n929 ;
  assign n1067 = n497 | n1066 ;
  assign n1068 = n877 & ~n1067 ;
  assign n1069 = ~n373 & n1068 ;
  assign n1070 = ~n1065 & n1069 ;
  assign n1071 = ~n158 & n1070 ;
  assign n1072 = ~n276 & n1071 ;
  assign n1073 = n144 | n201 ;
  assign n1074 = n664 | n1073 ;
  assign n1075 = n237 | n1074 ;
  assign n1076 = n1072 & ~n1075 ;
  assign n1077 = n401 | n413 ;
  assign n1078 = n405 | n573 ;
  assign n1079 = n1077 | n1078 ;
  assign n1080 = n141 | n282 ;
  assign n1081 = n153 | n1080 ;
  assign n1082 = n94 | n1081 ;
  assign n1083 = n668 | n1082 ;
  assign n1084 = n341 | n1083 ;
  assign n1085 = n418 | n1084 ;
  assign n1086 = n368 | n1085 ;
  assign n1087 = n124 | n1086 ;
  assign n1088 = n1079 | n1087 ;
  assign n1089 = n1076 & ~n1088 ;
  assign n1090 = n351 | n1020 ;
  assign n1091 = n726 | n1090 ;
  assign n1092 = n208 | n1091 ;
  assign n1093 = n518 | n881 ;
  assign n1094 = n308 | n1093 ;
  assign n1095 = n1019 | n1094 ;
  assign n1096 = n1092 | n1095 ;
  assign n1097 = n268 | n1096 ;
  assign n1098 = n184 | n203 ;
  assign n1099 = n1097 | n1098 ;
  assign n1100 = n129 | n206 ;
  assign n1101 = n160 | n1100 ;
  assign n1102 = n1099 | n1101 ;
  assign n1103 = n402 | n537 ;
  assign n1104 = n1102 | n1103 ;
  assign n1105 = n1089 & ~n1104 ;
  assign n1106 = n132 | n234 ;
  assign n1107 = n398 | n1106 ;
  assign n1108 = n1105 & ~n1107 ;
  assign n1109 = n1058 | n1108 ;
  assign n1110 = ~n894 & n1109 ;
  assign n1111 = n1058 & ~n1110 ;
  assign n1112 = ~n1058 & n1110 ;
  assign n1113 = ~pi6 & n823 ;
  assign n1114 = pi6 & ~n823 ;
  assign n1115 = n1113 | n1114 ;
  assign n1116 = n327 & n1115 ;
  assign n1117 = ~n1111 & n1116 ;
  assign n1118 = ~n1112 & n1117 ;
  assign n1119 = n1111 | n1118 ;
  assign n1120 = n1001 | n1007 ;
  assign n1121 = ~n1008 & n1120 ;
  assign n1122 = n1119 & n1121 ;
  assign n1123 = n1008 | n1122 ;
  assign n1124 = n894 & ~n942 ;
  assign n1125 = n695 | n1124 ;
  assign n1126 = n894 & n942 ;
  assign n1127 = n894 | n942 ;
  assign n1128 = ~n1126 & n1127 ;
  assign n1129 = n1125 & n1128 ;
  assign n1130 = n944 | n1128 ;
  assign n1131 = ( n332 & n1129 ) | ( n332 & ~n1130 ) | ( n1129 & ~n1130 );
  assign n1132 = ( n332 & n944 ) | ( n332 & n1130 ) | ( n944 & n1130 );
  assign n1133 = ~n1131 & n1132 ;
  assign n1134 = ~n829 & n1133 ;
  assign n1135 = n829 & ~n1133 ;
  assign n1136 = n1134 | n1135 ;
  assign n1137 = n266 & n966 ;
  assign n1138 = ~n266 & n968 ;
  assign n1139 = ( n587 & n782 ) | ( n587 & ~n1138 ) | ( n782 & ~n1138 );
  assign n1140 = ( n587 & ~n780 ) | ( n587 & n1138 ) | ( ~n780 & n1138 );
  assign n1141 = n1139 & ~n1140 ;
  assign n1142 = ~n1137 & n1141 ;
  assign n1143 = ~n1136 & n1142 ;
  assign n1144 = n1134 | n1143 ;
  assign n1145 = n1123 & n1144 ;
  assign n1146 = n1123 & ~n1145 ;
  assign n1147 = n1144 & ~n1145 ;
  assign n1148 = n1146 | n1147 ;
  assign n1149 = n327 & ~n953 ;
  assign n1150 = n949 & n1149 ;
  assign n1151 = n951 | n953 ;
  assign n1152 = ~n1150 & n1151 ;
  assign n1153 = n1148 & ~n1152 ;
  assign n1154 = n1145 | n1153 ;
  assign n1155 = ~n791 & n793 ;
  assign n1156 = n794 | n1155 ;
  assign n1157 = n1154 & ~n1156 ;
  assign n1158 = ( n980 & n1154 ) | ( n980 & ~n1156 ) | ( n1154 & ~n1156 );
  assign n1159 = ( ~n958 & n1157 ) | ( ~n958 & n1158 ) | ( n1157 & n1158 );
  assign n1160 = n987 & ~n989 ;
  assign n1161 = ~n987 & n989 ;
  assign n1162 = n1160 | n1161 ;
  assign n1163 = n1159 & ~n1162 ;
  assign n1164 = ~n1154 & n1156 ;
  assign n1165 = n1162 | n1164 ;
  assign n1166 = ( n995 & n1163 ) | ( n995 & ~n1165 ) | ( n1163 & ~n1165 );
  assign n1167 = n1148 & ~n1153 ;
  assign n1168 = n1152 | n1153 ;
  assign n1169 = ~n1167 & n1168 ;
  assign n1170 = n965 & ~n1169 ;
  assign n1171 = ( ~n965 & n1169 ) | ( ~n965 & n1170 ) | ( n1169 & n1170 );
  assign n1172 = n1170 | n1171 ;
  assign n1173 = n973 & ~n979 ;
  assign n1174 = ~n973 & n979 ;
  assign n1175 = n1173 | n1174 ;
  assign n1176 = n1136 & ~n1142 ;
  assign n1177 = n1143 | n1176 ;
  assign n1178 = n613 & n949 ;
  assign n1179 = n436 & ~n949 ;
  assign n1180 = ( n608 & n828 ) | ( n608 & ~n1179 ) | ( n828 & ~n1179 );
  assign n1181 = ( ~n439 & n828 ) | ( ~n439 & n1179 ) | ( n828 & n1179 );
  assign n1182 = n1180 & ~n1181 ;
  assign n1183 = ~n1178 & n1182 ;
  assign n1184 = n602 | n746 ;
  assign n1185 = ~n600 & n746 ;
  assign n1186 = n1184 & ~n1185 ;
  assign n1187 = ( n755 & n771 ) | ( n755 & ~n1186 ) | ( n771 & ~n1186 );
  assign n1188 = ( n755 & ~n759 ) | ( n755 & n1186 ) | ( ~n759 & n1186 );
  assign n1189 = ~n1187 & n1188 ;
  assign n1190 = n1125 & ~n1128 ;
  assign n1191 = ~n944 & n1128 ;
  assign n1192 = ~n266 & n1191 ;
  assign n1193 = n266 & n1129 ;
  assign n1194 = n1192 | n1193 ;
  assign n1195 = ( n332 & n1190 ) | ( n332 & n1194 ) | ( n1190 & n1194 );
  assign n1196 = ( n332 & n1130 ) | ( n332 & ~n1194 ) | ( n1130 & ~n1194 );
  assign n1197 = ~n1195 & n1196 ;
  assign n1198 = ( n1183 & n1189 ) | ( n1183 & n1197 ) | ( n1189 & n1197 );
  assign n1199 = ~n1177 & n1198 ;
  assign n1200 = n1119 | n1121 ;
  assign n1201 = ~n1122 & n1200 ;
  assign n1202 = n1177 | n1198 ;
  assign n1203 = ( ~n1198 & n1199 ) | ( ~n1198 & n1202 ) | ( n1199 & n1202 );
  assign n1204 = n1201 & ~n1203 ;
  assign n1205 = n1199 | n1204 ;
  assign n1206 = ( ~n1172 & n1175 ) | ( ~n1172 & n1205 ) | ( n1175 & n1205 );
  assign n1207 = ( n1172 & n1175 ) | ( n1172 & n1205 ) | ( n1175 & n1205 );
  assign n1208 = ( n1172 & n1206 ) | ( n1172 & ~n1207 ) | ( n1206 & ~n1207 );
  assign n1209 = n1112 | n1119 ;
  assign n1210 = n1116 & ~n1118 ;
  assign n1211 = n1209 & ~n1210 ;
  assign n1212 = n587 & n966 ;
  assign n1213 = ~n587 & n968 ;
  assign n1214 = ( n453 & n782 ) | ( n453 & ~n1213 ) | ( n782 & ~n1213 );
  assign n1215 = ( n453 & ~n780 ) | ( n453 & n1213 ) | ( ~n780 & n1213 );
  assign n1216 = n1214 & ~n1215 ;
  assign n1217 = ~n1212 & n1216 ;
  assign n1218 = ~n1211 & n1217 ;
  assign n1219 = ~pi22 & n739 ;
  assign n1220 = pi5 & ~n1219 ;
  assign n1221 = ~pi5 & n1219 ;
  assign n1222 = n1220 | n1221 ;
  assign n1223 = n327 & n1222 ;
  assign n1224 = ~n1058 & n1223 ;
  assign n1225 = n1058 & n1108 ;
  assign n1226 = n894 & ~n1225 ;
  assign n1227 = n1058 & ~n1108 ;
  assign n1228 = ~n1058 & n1108 ;
  assign n1229 = n1227 | n1228 ;
  assign n1230 = n1226 | n1229 ;
  assign n1231 = n332 & ~n1230 ;
  assign n1232 = n1110 | n1229 ;
  assign n1233 = n332 & ~n1232 ;
  assign n1234 = ( n1110 & ~n1231 ) | ( n1110 & n1233 ) | ( ~n1231 & n1233 );
  assign n1235 = ~n1224 & n1234 ;
  assign n1236 = n1058 & ~n1223 ;
  assign n1237 = ~n1224 & n1236 ;
  assign n1238 = ( n1224 & n1235 ) | ( n1224 & ~n1237 ) | ( n1235 & ~n1237 );
  assign n1239 = n1211 & ~n1217 ;
  assign n1240 = n1218 | n1239 ;
  assign n1241 = n1238 & ~n1240 ;
  assign n1242 = n1218 | n1241 ;
  assign n1243 = n266 & n1190 ;
  assign n1244 = n266 | n1130 ;
  assign n1245 = ( n587 & ~n1191 ) | ( n587 & n1244 ) | ( ~n1191 & n1244 );
  assign n1246 = ( n587 & n1129 ) | ( n587 & ~n1244 ) | ( n1129 & ~n1244 );
  assign n1247 = n1245 & ~n1246 ;
  assign n1248 = ~n1243 & n1247 ;
  assign n1249 = n453 & n966 ;
  assign n1250 = ~n453 & n968 ;
  assign n1251 = ( n755 & n782 ) | ( n755 & ~n1250 ) | ( n782 & ~n1250 );
  assign n1252 = ( n755 & ~n780 ) | ( n755 & n1250 ) | ( ~n780 & n1250 );
  assign n1253 = n1251 & ~n1252 ;
  assign n1254 = ~n1249 & n1253 ;
  assign n1255 = n746 & n771 ;
  assign n1256 = ~n746 & n759 ;
  assign n1257 = ( n602 & n949 ) | ( n602 & ~n1256 ) | ( n949 & ~n1256 );
  assign n1258 = ( ~n600 & n949 ) | ( ~n600 & n1256 ) | ( n949 & n1256 );
  assign n1259 = n1257 & ~n1258 ;
  assign n1260 = ~n1255 & n1259 ;
  assign n1261 = ( n1248 & n1254 ) | ( n1248 & n1260 ) | ( n1254 & n1260 );
  assign n1262 = ( n1183 & ~n1189 ) | ( n1183 & n1197 ) | ( ~n1189 & n1197 );
  assign n1263 = ( ~n1183 & n1189 ) | ( ~n1183 & n1262 ) | ( n1189 & n1262 );
  assign n1264 = ( ~n1197 & n1262 ) | ( ~n1197 & n1263 ) | ( n1262 & n1263 );
  assign n1265 = n1261 & n1264 ;
  assign n1266 = n613 & n828 ;
  assign n1267 = n436 & ~n828 ;
  assign n1268 = ( n608 & n1115 ) | ( n608 & ~n1267 ) | ( n1115 & ~n1267 );
  assign n1269 = ( ~n439 & n1115 ) | ( ~n439 & n1267 ) | ( n1115 & n1267 );
  assign n1270 = n1268 & ~n1269 ;
  assign n1271 = ~n1266 & n1270 ;
  assign n1272 = ~pi22 & n32 ;
  assign n1273 = ~pi4 & n1272 ;
  assign n1274 = pi4 & ~n1272 ;
  assign n1275 = n1273 | n1274 ;
  assign n1276 = n327 & n1275 ;
  assign n1277 = ~n1058 & n1276 ;
  assign n1278 = n1058 & ~n1276 ;
  assign n1279 = n1277 | n1278 ;
  assign n1280 = ~n1226 & n1229 ;
  assign n1281 = n332 & n1280 ;
  assign n1282 = ~n1110 & n1229 ;
  assign n1283 = ~n332 & n1282 ;
  assign n1284 = ( n266 & n1232 ) | ( n266 & ~n1283 ) | ( n1232 & ~n1283 );
  assign n1285 = ( n266 & ~n1230 ) | ( n266 & n1283 ) | ( ~n1230 & n1283 );
  assign n1286 = n1284 & ~n1285 ;
  assign n1287 = ~n1281 & n1286 ;
  assign n1288 = ~n1279 & n1287 ;
  assign n1289 = n1277 | n1288 ;
  assign n1290 = n1271 & n1289 ;
  assign n1291 = n1271 | n1289 ;
  assign n1292 = ~n1290 & n1291 ;
  assign n1293 = n755 & n966 ;
  assign n1294 = ~n755 & n968 ;
  assign n1295 = ( n746 & n782 ) | ( n746 & ~n1294 ) | ( n782 & ~n1294 );
  assign n1296 = ( n746 & ~n780 ) | ( n746 & n1294 ) | ( ~n780 & n1294 );
  assign n1297 = n1295 & ~n1296 ;
  assign n1298 = ~n1293 & n1297 ;
  assign n1299 = n587 & n1190 ;
  assign n1300 = n587 | n1130 ;
  assign n1301 = ( n453 & ~n1191 ) | ( n453 & n1300 ) | ( ~n1191 & n1300 );
  assign n1302 = ( n453 & n1129 ) | ( n453 & ~n1300 ) | ( n1129 & ~n1300 );
  assign n1303 = n1301 & ~n1302 ;
  assign n1304 = ~n1299 & n1303 ;
  assign n1305 = n771 & n949 ;
  assign n1306 = n759 & ~n949 ;
  assign n1307 = ( n602 & n828 ) | ( n602 & ~n1306 ) | ( n828 & ~n1306 );
  assign n1308 = ( ~n600 & n828 ) | ( ~n600 & n1306 ) | ( n828 & n1306 );
  assign n1309 = n1307 & ~n1308 ;
  assign n1310 = ~n1305 & n1309 ;
  assign n1311 = ( n1298 & n1304 ) | ( n1298 & n1310 ) | ( n1304 & n1310 );
  assign n1312 = n1292 & n1311 ;
  assign n1313 = n1290 | n1312 ;
  assign n1314 = n1261 | n1264 ;
  assign n1315 = ~n1265 & n1314 ;
  assign n1316 = n1313 & n1315 ;
  assign n1317 = n1265 | n1316 ;
  assign n1318 = ~n1201 & n1203 ;
  assign n1319 = n1204 | n1318 ;
  assign n1320 = ( n1242 & n1317 ) | ( n1242 & ~n1319 ) | ( n1317 & ~n1319 );
  assign n1321 = n1208 & ~n1320 ;
  assign n1322 = ~n1208 & n1320 ;
  assign n1323 = n1321 | n1322 ;
  assign n1324 = ( ~n1242 & n1317 ) | ( ~n1242 & n1319 ) | ( n1317 & n1319 );
  assign n1325 = ( n1242 & ~n1319 ) | ( n1242 & n1324 ) | ( ~n1319 & n1324 );
  assign n1326 = ( ~n1317 & n1324 ) | ( ~n1317 & n1325 ) | ( n1324 & n1325 );
  assign n1327 = ~n1238 & n1240 ;
  assign n1328 = n1241 | n1327 ;
  assign n1329 = n1236 | n1238 ;
  assign n1330 = n1234 & n1236 ;
  assign n1331 = ( n1234 & ~n1235 ) | ( n1234 & n1330 ) | ( ~n1235 & n1330 );
  assign n1332 = n608 | n1222 ;
  assign n1333 = ~n439 & n1222 ;
  assign n1334 = n1332 & ~n1333 ;
  assign n1335 = ( ~n436 & n1115 ) | ( ~n436 & n1334 ) | ( n1115 & n1334 );
  assign n1336 = ( n613 & n1115 ) | ( n613 & ~n1334 ) | ( n1115 & ~n1334 );
  assign n1337 = n1335 & ~n1336 ;
  assign n1338 = pi3 & ~n258 ;
  assign n1339 = ~pi3 & n258 ;
  assign n1340 = n1338 | n1339 ;
  assign n1341 = n327 & n1340 ;
  assign n1342 = n102 | n168 ;
  assign n1343 = n153 | n485 ;
  assign n1344 = n1342 | n1343 ;
  assign n1345 = n486 | n567 ;
  assign n1346 = n201 | n414 ;
  assign n1347 = n209 | n718 ;
  assign n1348 = n164 | n1347 ;
  assign n1349 = n349 | n1348 ;
  assign n1350 = n107 | n1349 ;
  assign n1351 = n205 | n1350 ;
  assign n1352 = n352 | n1351 ;
  assign n1353 = n271 | n273 ;
  assign n1354 = ~n356 & n877 ;
  assign n1355 = n162 | n335 ;
  assign n1356 = n1354 & ~n1355 ;
  assign n1357 = n368 | n409 ;
  assign n1358 = n239 | n1357 ;
  assign n1359 = n1356 & ~n1358 ;
  assign n1360 = n507 | n928 ;
  assign n1361 = n208 | n305 ;
  assign n1362 = n402 | n1361 ;
  assign n1363 = n472 | n544 ;
  assign n1364 = n1362 | n1363 ;
  assign n1365 = n1360 | n1364 ;
  assign n1366 = n311 | n1365 ;
  assign n1367 = n207 | n1366 ;
  assign n1368 = n272 | n1367 ;
  assign n1369 = n211 | n1368 ;
  assign n1370 = n367 | n1369 ;
  assign n1371 = n144 | n370 ;
  assign n1372 = n529 | n1371 ;
  assign n1373 = n1370 | n1372 ;
  assign n1374 = n1359 & ~n1373 ;
  assign n1375 = ~n1353 & n1374 ;
  assign n1376 = ~n1352 & n1375 ;
  assign n1377 = ~n1346 & n1376 ;
  assign n1378 = ~n1345 & n1377 ;
  assign n1379 = ~n1344 & n1378 ;
  assign n1380 = ~n204 & n1379 ;
  assign n1381 = n332 & n1380 ;
  assign n1382 = n1058 | n1381 ;
  assign n1383 = n1341 & ~n1382 ;
  assign n1384 = n266 & n1280 ;
  assign n1385 = ~n266 & n1282 ;
  assign n1386 = ( n587 & n1232 ) | ( n587 & ~n1385 ) | ( n1232 & ~n1385 );
  assign n1387 = ( n587 & ~n1230 ) | ( n587 & n1385 ) | ( ~n1230 & n1385 );
  assign n1388 = n1386 & ~n1387 ;
  assign n1389 = ~n1384 & n1388 ;
  assign n1390 = ~n1341 & n1382 ;
  assign n1391 = n1383 | n1390 ;
  assign n1392 = n1389 & ~n1391 ;
  assign n1393 = n1383 | n1392 ;
  assign n1394 = n1337 & n1393 ;
  assign n1395 = n1337 | n1393 ;
  assign n1396 = ~n1394 & n1395 ;
  assign n1397 = n746 & n966 ;
  assign n1398 = ~n746 & n968 ;
  assign n1399 = ( n782 & n949 ) | ( n782 & ~n1398 ) | ( n949 & ~n1398 );
  assign n1400 = ( ~n780 & n949 ) | ( ~n780 & n1398 ) | ( n949 & n1398 );
  assign n1401 = n1399 & ~n1400 ;
  assign n1402 = ~n1397 & n1401 ;
  assign n1403 = n453 & n1190 ;
  assign n1404 = n453 | n1130 ;
  assign n1405 = ( n755 & ~n1191 ) | ( n755 & n1404 ) | ( ~n1191 & n1404 );
  assign n1406 = ( n755 & n1129 ) | ( n755 & ~n1404 ) | ( n1129 & ~n1404 );
  assign n1407 = n1405 & ~n1406 ;
  assign n1408 = ~n1403 & n1407 ;
  assign n1409 = n771 & n828 ;
  assign n1410 = n759 & ~n828 ;
  assign n1411 = ( n602 & n1115 ) | ( n602 & ~n1410 ) | ( n1115 & ~n1410 );
  assign n1412 = ( ~n600 & n1115 ) | ( ~n600 & n1410 ) | ( n1115 & n1410 );
  assign n1413 = n1411 & ~n1412 ;
  assign n1414 = ~n1409 & n1413 ;
  assign n1415 = ( n1402 & n1408 ) | ( n1402 & n1414 ) | ( n1408 & n1414 );
  assign n1416 = n1396 & n1415 ;
  assign n1417 = n1394 | n1416 ;
  assign n1418 = ( n1248 & n1260 ) | ( n1248 & ~n1261 ) | ( n1260 & ~n1261 );
  assign n1419 = ( n1254 & ~n1261 ) | ( n1254 & n1418 ) | ( ~n1261 & n1418 );
  assign n1420 = ( n1331 & n1417 ) | ( n1331 & n1419 ) | ( n1417 & n1419 );
  assign n1421 = n1417 | n1419 ;
  assign n1422 = ( ~n1329 & n1420 ) | ( ~n1329 & n1421 ) | ( n1420 & n1421 );
  assign n1423 = ~n1328 & n1422 ;
  assign n1424 = n1328 & ~n1422 ;
  assign n1425 = n1423 | n1424 ;
  assign n1426 = n1313 | n1315 ;
  assign n1427 = ~n1316 & n1426 ;
  assign n1428 = n1423 | n1427 ;
  assign n1429 = ( n1423 & ~n1425 ) | ( n1423 & n1428 ) | ( ~n1425 & n1428 );
  assign n1430 = n1326 & ~n1429 ;
  assign n1431 = n1323 | n1430 ;
  assign n1432 = ~n1159 & n1162 ;
  assign n1433 = n1162 & n1164 ;
  assign n1434 = ( ~n995 & n1432 ) | ( ~n995 & n1433 ) | ( n1432 & n1433 );
  assign n1435 = n1166 | n1434 ;
  assign n1436 = n965 | n1175 ;
  assign n1437 = n965 & n1175 ;
  assign n1438 = n1436 & ~n1437 ;
  assign n1439 = ( ~n1169 & n1205 ) | ( ~n1169 & n1438 ) | ( n1205 & n1438 );
  assign n1440 = n1157 | n1164 ;
  assign n1441 = ( n958 & n980 ) | ( n958 & ~n1440 ) | ( n980 & ~n1440 );
  assign n1442 = ( n958 & n980 ) | ( n958 & ~n1441 ) | ( n980 & ~n1441 );
  assign n1443 = ( n1440 & n1441 ) | ( n1440 & ~n1442 ) | ( n1441 & ~n1442 );
  assign n1444 = n1439 & ~n1443 ;
  assign n1445 = n1439 & n1443 ;
  assign n1446 = ( n1443 & n1444 ) | ( n1443 & ~n1445 ) | ( n1444 & ~n1445 );
  assign n1447 = n1322 | n1444 ;
  assign n1448 = ( n1444 & ~n1446 ) | ( n1444 & n1447 ) | ( ~n1446 & n1447 );
  assign n1449 = ~n1435 & n1448 ;
  assign n1450 = ~n1435 & n1444 ;
  assign n1451 = ( n1435 & n1446 ) | ( n1435 & ~n1450 ) | ( n1446 & ~n1450 );
  assign n1452 = ( n1431 & ~n1449 ) | ( n1431 & n1451 ) | ( ~n1449 & n1451 );
  assign n1453 = ~n1323 & n1429 ;
  assign n1454 = ~n1326 & n1453 ;
  assign n1455 = ( n1449 & ~n1451 ) | ( n1449 & n1454 ) | ( ~n1451 & n1454 );
  assign n1456 = ~n1425 & n1427 ;
  assign n1457 = n1425 & ~n1427 ;
  assign n1458 = n1456 | n1457 ;
  assign n1459 = n1292 | n1311 ;
  assign n1460 = ~n1312 & n1459 ;
  assign n1461 = n1279 & ~n1287 ;
  assign n1462 = n1288 | n1461 ;
  assign n1463 = n431 | n1340 ;
  assign n1464 = n608 & n1463 ;
  assign n1465 = n613 & n1340 ;
  assign n1466 = n431 & ~n1465 ;
  assign n1467 = n1464 & n1466 ;
  assign n1468 = n1058 & ~n1380 ;
  assign n1469 = n1380 | n1468 ;
  assign n1470 = n332 & ~n1469 ;
  assign n1471 = ~n332 & n1468 ;
  assign n1472 = n266 | n1058 ;
  assign n1473 = n1380 & n1472 ;
  assign n1474 = n1471 | n1473 ;
  assign n1475 = n1470 | n1474 ;
  assign n1476 = n1467 & ~n1475 ;
  assign n1477 = n608 | n1275 ;
  assign n1478 = ~n439 & n1275 ;
  assign n1479 = n1477 & ~n1478 ;
  assign n1480 = ( ~n436 & n1222 ) | ( ~n436 & n1479 ) | ( n1222 & n1479 );
  assign n1481 = ( n613 & n1222 ) | ( n613 & ~n1479 ) | ( n1222 & ~n1479 );
  assign n1482 = n1480 & ~n1481 ;
  assign n1483 = n1476 & n1482 ;
  assign n1484 = n1476 | n1482 ;
  assign n1485 = ~n1483 & n1484 ;
  assign n1486 = n755 & n1190 ;
  assign n1487 = n755 | n1130 ;
  assign n1488 = ( n746 & ~n1191 ) | ( n746 & n1487 ) | ( ~n1191 & n1487 );
  assign n1489 = ( n746 & n1129 ) | ( n746 & ~n1487 ) | ( n1129 & ~n1487 );
  assign n1490 = n1488 & ~n1489 ;
  assign n1491 = ~n1486 & n1490 ;
  assign n1492 = n949 & n966 ;
  assign n1493 = ~n949 & n968 ;
  assign n1494 = ( n782 & n828 ) | ( n782 & ~n1493 ) | ( n828 & ~n1493 );
  assign n1495 = ( ~n780 & n828 ) | ( ~n780 & n1493 ) | ( n828 & n1493 );
  assign n1496 = n1494 & ~n1495 ;
  assign n1497 = ~n1492 & n1496 ;
  assign n1498 = n771 & n1115 ;
  assign n1499 = n759 & ~n1115 ;
  assign n1500 = ( n602 & n1222 ) | ( n602 & ~n1499 ) | ( n1222 & ~n1499 );
  assign n1501 = ( ~n600 & n1222 ) | ( ~n600 & n1499 ) | ( n1222 & n1499 );
  assign n1502 = n1500 & ~n1501 ;
  assign n1503 = ~n1498 & n1502 ;
  assign n1504 = ( n1491 & n1497 ) | ( n1491 & n1503 ) | ( n1497 & n1503 );
  assign n1505 = n1483 | n1504 ;
  assign n1506 = ( n1483 & n1485 ) | ( n1483 & n1505 ) | ( n1485 & n1505 );
  assign n1507 = ( n1298 & n1310 ) | ( n1298 & ~n1311 ) | ( n1310 & ~n1311 );
  assign n1508 = ( n1304 & ~n1311 ) | ( n1304 & n1507 ) | ( ~n1311 & n1507 );
  assign n1509 = ( ~n1462 & n1506 ) | ( ~n1462 & n1508 ) | ( n1506 & n1508 );
  assign n1510 = n1460 & n1509 ;
  assign n1511 = n1329 & ~n1331 ;
  assign n1512 = ( n1331 & ~n1417 ) | ( n1331 & n1419 ) | ( ~n1417 & n1419 );
  assign n1513 = n1417 & ~n1419 ;
  assign n1514 = ( n1329 & ~n1512 ) | ( n1329 & n1513 ) | ( ~n1512 & n1513 );
  assign n1515 = ( n1417 & n1511 ) | ( n1417 & ~n1514 ) | ( n1511 & ~n1514 );
  assign n1516 = n1460 | n1509 ;
  assign n1517 = ~n1510 & n1516 ;
  assign n1518 = ~n1514 & n1517 ;
  assign n1519 = ~n1419 & n1517 ;
  assign n1520 = ( n1515 & n1518 ) | ( n1515 & n1519 ) | ( n1518 & n1519 );
  assign n1521 = n1510 | n1520 ;
  assign n1522 = ~n1458 & n1521 ;
  assign n1523 = n1458 & ~n1521 ;
  assign n1524 = n1522 | n1523 ;
  assign n1525 = n1514 & ~n1517 ;
  assign n1526 = n1419 & ~n1517 ;
  assign n1527 = ( ~n1515 & n1525 ) | ( ~n1515 & n1526 ) | ( n1525 & n1526 );
  assign n1528 = n1520 | n1527 ;
  assign n1529 = n1396 | n1415 ;
  assign n1530 = ~n1416 & n1529 ;
  assign n1531 = ~n1467 & n1475 ;
  assign n1532 = n1476 | n1531 ;
  assign n1533 = n608 | n1340 ;
  assign n1534 = ~n439 & n1340 ;
  assign n1535 = n1533 & ~n1534 ;
  assign n1536 = ( ~n436 & n1275 ) | ( ~n436 & n1535 ) | ( n1275 & n1535 );
  assign n1537 = ( n613 & n1275 ) | ( n613 & ~n1535 ) | ( n1275 & ~n1535 );
  assign n1538 = n1536 & ~n1537 ;
  assign n1539 = ~n1389 & n1391 ;
  assign n1540 = n1392 | n1539 ;
  assign n1541 = n1538 & ~n1540 ;
  assign n1542 = n587 & n1280 ;
  assign n1543 = ~n587 & n1282 ;
  assign n1544 = ( n453 & n1232 ) | ( n453 & ~n1543 ) | ( n1232 & ~n1543 );
  assign n1545 = ( n453 & ~n1230 ) | ( n453 & n1543 ) | ( ~n1230 & n1543 );
  assign n1546 = n1544 & ~n1545 ;
  assign n1547 = ~n1542 & n1546 ;
  assign n1548 = ~n1540 & n1547 ;
  assign n1549 = ( ~n1532 & n1541 ) | ( ~n1532 & n1548 ) | ( n1541 & n1548 );
  assign n1550 = ~n1538 & n1540 ;
  assign n1551 = n1540 & ~n1547 ;
  assign n1552 = ( n1532 & n1550 ) | ( n1532 & n1551 ) | ( n1550 & n1551 );
  assign n1553 = n1549 | n1552 ;
  assign n1554 = ( n1402 & n1414 ) | ( n1402 & ~n1415 ) | ( n1414 & ~n1415 );
  assign n1555 = ( n1408 & ~n1415 ) | ( n1408 & n1554 ) | ( ~n1415 & n1554 );
  assign n1556 = n1549 | n1555 ;
  assign n1557 = ( n1549 & ~n1553 ) | ( n1549 & n1556 ) | ( ~n1553 & n1556 );
  assign n1558 = n1530 & n1557 ;
  assign n1559 = n1530 | n1557 ;
  assign n1560 = ~n1558 & n1559 ;
  assign n1561 = ( n1462 & n1506 ) | ( n1462 & ~n1508 ) | ( n1506 & ~n1508 );
  assign n1562 = ( ~n1506 & n1509 ) | ( ~n1506 & n1561 ) | ( n1509 & n1561 );
  assign n1563 = n1560 & ~n1562 ;
  assign n1564 = n1558 | n1563 ;
  assign n1565 = ~n1560 & n1562 ;
  assign n1566 = n1563 | n1565 ;
  assign n1567 = n1485 & n1504 ;
  assign n1568 = n1485 | n1504 ;
  assign n1569 = ~n1567 & n1568 ;
  assign n1570 = n453 & n1280 ;
  assign n1571 = ~n453 & n1282 ;
  assign n1572 = ( n755 & n1232 ) | ( n755 & ~n1571 ) | ( n1232 & ~n1571 );
  assign n1573 = ( n755 & ~n1230 ) | ( n755 & n1571 ) | ( ~n1230 & n1571 );
  assign n1574 = n1572 & ~n1573 ;
  assign n1575 = ~n1570 & n1574 ;
  assign n1576 = n587 | n1058 ;
  assign n1577 = n1380 & n1576 ;
  assign n1578 = ( n266 & n1058 ) | ( n266 & n1380 ) | ( n1058 & n1380 );
  assign n1579 = ( n1472 & n1577 ) | ( n1472 & ~n1578 ) | ( n1577 & ~n1578 );
  assign n1580 = n771 & n1222 ;
  assign n1581 = n759 & ~n1222 ;
  assign n1582 = ( n602 & n1275 ) | ( n602 & ~n1581 ) | ( n1275 & ~n1581 );
  assign n1583 = ( ~n600 & n1275 ) | ( ~n600 & n1581 ) | ( n1275 & n1581 );
  assign n1584 = n1582 & ~n1583 ;
  assign n1585 = ~n1580 & n1584 ;
  assign n1586 = ( n1575 & ~n1579 ) | ( n1575 & n1585 ) | ( ~n1579 & n1585 );
  assign n1587 = n746 & n1190 ;
  assign n1588 = n746 | n1130 ;
  assign n1589 = ( n949 & ~n1191 ) | ( n949 & n1588 ) | ( ~n1191 & n1588 );
  assign n1590 = ( n949 & n1129 ) | ( n949 & ~n1588 ) | ( n1129 & ~n1588 );
  assign n1591 = n1589 & ~n1590 ;
  assign n1592 = ~n1587 & n1591 ;
  assign n1593 = n828 & n966 ;
  assign n1594 = ~n828 & n968 ;
  assign n1595 = ( n782 & n1115 ) | ( n782 & ~n1594 ) | ( n1115 & ~n1594 );
  assign n1596 = ( ~n780 & n1115 ) | ( ~n780 & n1594 ) | ( n1115 & n1594 );
  assign n1597 = n1595 & ~n1596 ;
  assign n1598 = ~n1593 & n1597 ;
  assign n1599 = n453 | n1058 ;
  assign n1600 = n1380 & n1599 ;
  assign n1601 = ( n587 & n1058 ) | ( n587 & n1380 ) | ( n1058 & n1380 );
  assign n1602 = ( n1576 & n1600 ) | ( n1576 & ~n1601 ) | ( n1600 & ~n1601 );
  assign n1603 = n771 & n1340 ;
  assign n1604 = n578 & ~n1603 ;
  assign n1605 = ~n1602 & n1604 ;
  assign n1606 = ( n1592 & n1598 ) | ( n1592 & n1605 ) | ( n1598 & n1605 );
  assign n1607 = ( n1491 & n1503 ) | ( n1491 & ~n1504 ) | ( n1503 & ~n1504 );
  assign n1608 = ( n1497 & ~n1504 ) | ( n1497 & n1607 ) | ( ~n1504 & n1607 );
  assign n1609 = ( n1586 & n1606 ) | ( n1586 & n1608 ) | ( n1606 & n1608 );
  assign n1610 = n1569 & n1609 ;
  assign n1611 = n1569 | n1609 ;
  assign n1612 = ~n1610 & n1611 ;
  assign n1613 = n1552 | n1556 ;
  assign n1614 = n1553 & n1555 ;
  assign n1615 = n1613 & ~n1614 ;
  assign n1616 = ~n1610 & n1615 ;
  assign n1617 = ( n1610 & n1612 ) | ( n1610 & ~n1616 ) | ( n1612 & ~n1616 );
  assign n1618 = ~n1566 & n1617 ;
  assign n1619 = n1612 & ~n1615 ;
  assign n1620 = ~n1612 & n1615 ;
  assign n1621 = n1619 | n1620 ;
  assign n1622 = n746 | n1232 ;
  assign n1623 = n746 & ~n1230 ;
  assign n1624 = n1622 & ~n1623 ;
  assign n1625 = ( n755 & n1280 ) | ( n755 & ~n1624 ) | ( n1280 & ~n1624 );
  assign n1626 = ( n755 & ~n1282 ) | ( n755 & n1624 ) | ( ~n1282 & n1624 );
  assign n1627 = ~n1625 & n1626 ;
  assign n1628 = n782 | n1222 ;
  assign n1629 = ~n780 & n1222 ;
  assign n1630 = n1628 & ~n1629 ;
  assign n1631 = ( ~n968 & n1115 ) | ( ~n968 & n1630 ) | ( n1115 & n1630 );
  assign n1632 = ( n966 & n1115 ) | ( n966 & ~n1630 ) | ( n1115 & ~n1630 );
  assign n1633 = n1631 & ~n1632 ;
  assign n1634 = ~n828 & n1191 ;
  assign n1635 = n828 & n1129 ;
  assign n1636 = n1634 | n1635 ;
  assign n1637 = ( n949 & n1130 ) | ( n949 & ~n1636 ) | ( n1130 & ~n1636 );
  assign n1638 = ( n949 & n1190 ) | ( n949 & n1636 ) | ( n1190 & n1636 );
  assign n1639 = n1637 & ~n1638 ;
  assign n1640 = ( n1627 & n1633 ) | ( n1627 & n1639 ) | ( n1633 & n1639 );
  assign n1641 = ~n1467 & n1640 ;
  assign n1642 = ~n431 & n1465 ;
  assign n1643 = ( n431 & n1464 ) | ( n431 & ~n1642 ) | ( n1464 & ~n1642 );
  assign n1644 = n1641 & n1643 ;
  assign n1645 = n1467 | n1643 ;
  assign n1646 = ( n1467 & n1641 ) | ( n1467 & n1645 ) | ( n1641 & n1645 );
  assign n1647 = n1643 & ~n1646 ;
  assign n1650 = ( n1592 & n1605 ) | ( n1592 & ~n1606 ) | ( n1605 & ~n1606 );
  assign n1651 = ( n1598 & ~n1606 ) | ( n1598 & n1650 ) | ( ~n1606 & n1650 );
  assign n1648 = n1640 & ~n1643 ;
  assign n1649 = ( n1640 & ~n1641 ) | ( n1640 & n1648 ) | ( ~n1641 & n1648 );
  assign n1652 = n1649 & n1651 ;
  assign n1653 = ( n1647 & n1651 ) | ( n1647 & n1652 ) | ( n1651 & n1652 );
  assign n1654 = n1644 | n1653 ;
  assign n1655 = ( ~n1586 & n1606 ) | ( ~n1586 & n1608 ) | ( n1606 & n1608 );
  assign n1656 = ( n1586 & ~n1606 ) | ( n1586 & n1655 ) | ( ~n1606 & n1655 );
  assign n1657 = ( ~n1608 & n1655 ) | ( ~n1608 & n1656 ) | ( n1655 & n1656 );
  assign n1658 = ( ~n1532 & n1538 ) | ( ~n1532 & n1547 ) | ( n1538 & n1547 );
  assign n1659 = ( n1532 & ~n1538 ) | ( n1532 & n1658 ) | ( ~n1538 & n1658 );
  assign n1660 = ( ~n1547 & n1658 ) | ( ~n1547 & n1659 ) | ( n1658 & n1659 );
  assign n1661 = ( n1654 & n1657 ) | ( n1654 & ~n1660 ) | ( n1657 & ~n1660 );
  assign n1662 = ~n1621 & n1661 ;
  assign n1663 = n1621 & ~n1661 ;
  assign n1664 = n1662 | n1663 ;
  assign n1665 = n1654 & n1660 ;
  assign n1666 = n1654 | n1660 ;
  assign n1667 = ~n1665 & n1666 ;
  assign n1668 = n1657 & ~n1667 ;
  assign n1672 = n1602 & ~n1604 ;
  assign n1673 = n1605 | n1672 ;
  assign n1674 = n771 & n1275 ;
  assign n1675 = n759 & ~n1275 ;
  assign n1676 = ( n602 & n1340 ) | ( n602 & ~n1675 ) | ( n1340 & ~n1675 );
  assign n1677 = ( ~n600 & n1340 ) | ( ~n600 & n1675 ) | ( n1340 & n1675 );
  assign n1678 = n1676 & ~n1677 ;
  assign n1679 = ~n1674 & n1678 ;
  assign n1680 = ~n1673 & n1679 ;
  assign n1681 = n949 | n1232 ;
  assign n1682 = n949 & ~n1230 ;
  assign n1683 = n1681 & ~n1682 ;
  assign n1684 = ( n746 & n1280 ) | ( n746 & ~n1683 ) | ( n1280 & ~n1683 );
  assign n1685 = ( n746 & ~n1282 ) | ( n746 & n1683 ) | ( ~n1282 & n1683 );
  assign n1686 = ~n1684 & n1685 ;
  assign n1687 = ~n1115 & n1191 ;
  assign n1688 = n1115 & n1129 ;
  assign n1689 = n1687 | n1688 ;
  assign n1690 = ( n828 & n1130 ) | ( n828 & ~n1689 ) | ( n1130 & ~n1689 );
  assign n1691 = ( n828 & n1190 ) | ( n828 & n1689 ) | ( n1190 & n1689 );
  assign n1692 = n1690 & ~n1691 ;
  assign n1693 = n755 | n1058 ;
  assign n1694 = n1380 & n1693 ;
  assign n1695 = ( n453 & n1058 ) | ( n453 & n1380 ) | ( n1058 & n1380 );
  assign n1696 = ( n1599 & n1694 ) | ( n1599 & ~n1695 ) | ( n1694 & ~n1695 );
  assign n1697 = ( n1686 & n1692 ) | ( n1686 & ~n1696 ) | ( n1692 & ~n1696 );
  assign n1698 = n1679 & ~n1680 ;
  assign n1699 = ( n1673 & n1680 ) | ( n1673 & ~n1698 ) | ( n1680 & ~n1698 );
  assign n1700 = n1697 & ~n1699 ;
  assign n1701 = n1680 | n1700 ;
  assign n1669 = ( n1575 & n1579 ) | ( n1575 & n1585 ) | ( n1579 & n1585 );
  assign n1670 = ( n1579 & n1585 ) | ( n1579 & ~n1669 ) | ( n1585 & ~n1669 );
  assign n1671 = ( n1575 & ~n1669 ) | ( n1575 & n1670 ) | ( ~n1669 & n1670 );
  assign n1702 = ~n1671 & n1701 ;
  assign n1703 = n1701 & ~n1702 ;
  assign n1704 = n1671 | n1702 ;
  assign n1705 = ~n1703 & n1704 ;
  assign n1706 = n1649 | n1651 ;
  assign n1707 = n1647 | n1706 ;
  assign n1708 = ~n1653 & n1707 ;
  assign n1709 = ~n1705 & n1708 ;
  assign n1710 = n1705 & ~n1708 ;
  assign n1711 = n1709 | n1710 ;
  assign n1712 = ( n1686 & n1692 ) | ( n1686 & ~n1697 ) | ( n1692 & ~n1697 );
  assign n1713 = n828 | n1232 ;
  assign n1714 = n828 & ~n1230 ;
  assign n1715 = n1713 & ~n1714 ;
  assign n1716 = ( n949 & n1280 ) | ( n949 & ~n1715 ) | ( n1280 & ~n1715 );
  assign n1717 = ( n949 & ~n1282 ) | ( n949 & n1715 ) | ( ~n1282 & n1715 );
  assign n1718 = ~n1716 & n1717 ;
  assign n1719 = n1191 & ~n1222 ;
  assign n1720 = n1129 & n1222 ;
  assign n1721 = n1719 | n1720 ;
  assign n1722 = ( n1115 & n1130 ) | ( n1115 & ~n1721 ) | ( n1130 & ~n1721 );
  assign n1723 = ( n1115 & n1190 ) | ( n1115 & n1721 ) | ( n1190 & n1721 );
  assign n1724 = n1722 & ~n1723 ;
  assign n1725 = n782 | n1340 ;
  assign n1726 = ~n780 & n1340 ;
  assign n1727 = n1725 & ~n1726 ;
  assign n1728 = ( ~n968 & n1275 ) | ( ~n968 & n1727 ) | ( n1275 & n1727 );
  assign n1729 = ( n966 & n1275 ) | ( n966 & ~n1727 ) | ( n1275 & ~n1727 );
  assign n1730 = n1728 & ~n1729 ;
  assign n1731 = ( n1718 & n1724 ) | ( n1718 & n1730 ) | ( n1724 & n1730 );
  assign n1732 = ~n1697 & n1731 ;
  assign n1733 = ~n1696 & n1731 ;
  assign n1734 = ( n1712 & n1732 ) | ( n1712 & n1733 ) | ( n1732 & n1733 );
  assign n1735 = ( n1696 & n1697 ) | ( n1696 & ~n1712 ) | ( n1697 & ~n1712 );
  assign n1736 = n1734 | n1735 ;
  assign n1737 = n782 | n1275 ;
  assign n1738 = ~n780 & n1275 ;
  assign n1739 = n1737 & ~n1738 ;
  assign n1740 = ( ~n968 & n1222 ) | ( ~n968 & n1739 ) | ( n1222 & n1739 );
  assign n1741 = ( n966 & n1222 ) | ( n966 & ~n1739 ) | ( n1222 & ~n1739 );
  assign n1742 = n1740 & ~n1741 ;
  assign n1743 = n599 & n1340 ;
  assign n1744 = n738 | n1340 ;
  assign n1745 = n782 & n1744 ;
  assign n1746 = n966 & n1340 ;
  assign n1747 = n738 & ~n1746 ;
  assign n1748 = n1745 & n1747 ;
  assign n1749 = n746 | n1058 ;
  assign n1750 = n1380 & n1749 ;
  assign n1751 = ( n755 & n1058 ) | ( n755 & n1380 ) | ( n1058 & n1380 );
  assign n1752 = ( n1693 & n1750 ) | ( n1693 & ~n1751 ) | ( n1750 & ~n1751 );
  assign n1753 = n1748 & ~n1752 ;
  assign n1754 = ( n1742 & n1743 ) | ( n1742 & ~n1753 ) | ( n1743 & ~n1753 );
  assign n1755 = ( ~n1743 & n1753 ) | ( ~n1743 & n1754 ) | ( n1753 & n1754 );
  assign n1756 = ( ~n1742 & n1754 ) | ( ~n1742 & n1755 ) | ( n1754 & n1755 );
  assign n1757 = n1697 & n1731 ;
  assign n1758 = n1696 & n1731 ;
  assign n1759 = ( ~n1712 & n1757 ) | ( ~n1712 & n1758 ) | ( n1757 & n1758 );
  assign n1760 = n1756 & n1759 ;
  assign n1761 = ( ~n1736 & n1756 ) | ( ~n1736 & n1760 ) | ( n1756 & n1760 );
  assign n1762 = n1734 | n1761 ;
  assign n1763 = ( n1627 & n1633 ) | ( n1627 & ~n1639 ) | ( n1633 & ~n1639 );
  assign n1764 = ( n1627 & n1633 ) | ( n1627 & ~n1763 ) | ( n1633 & ~n1763 );
  assign n1765 = ( n1742 & n1743 ) | ( n1742 & n1753 ) | ( n1743 & n1753 );
  assign n1766 = n1763 & n1765 ;
  assign n1767 = n1639 & n1765 ;
  assign n1768 = ( ~n1764 & n1766 ) | ( ~n1764 & n1767 ) | ( n1766 & n1767 );
  assign n1769 = n1763 | n1765 ;
  assign n1770 = n1639 | n1765 ;
  assign n1771 = ( ~n1764 & n1769 ) | ( ~n1764 & n1770 ) | ( n1769 & n1770 );
  assign n1772 = ~n1768 & n1771 ;
  assign n1773 = ~n1697 & n1699 ;
  assign n1774 = n1700 | n1773 ;
  assign n1775 = ~n1772 & n1774 ;
  assign n1776 = n1772 & ~n1774 ;
  assign n1777 = n1775 | n1776 ;
  assign n1778 = ( n1718 & n1724 ) | ( n1718 & ~n1730 ) | ( n1724 & ~n1730 );
  assign n1779 = ( n1718 & n1724 ) | ( n1718 & ~n1778 ) | ( n1724 & ~n1778 );
  assign n1780 = ( n1730 & n1778 ) | ( n1730 & ~n1779 ) | ( n1778 & ~n1779 );
  assign n1781 = n944 & ~n1191 ;
  assign n1782 = ( n1190 & n1340 ) | ( n1190 & ~n1781 ) | ( n1340 & ~n1781 );
  assign n1783 = n1781 & ~n1782 ;
  assign n1784 = n828 | n1058 ;
  assign n1785 = n1380 & n1784 ;
  assign n1786 = n949 | n1058 ;
  assign n1787 = ( n949 & n1058 ) | ( n949 & n1380 ) | ( n1058 & n1380 );
  assign n1788 = ( n1785 & n1786 ) | ( n1785 & ~n1787 ) | ( n1786 & ~n1787 );
  assign n1789 = n1783 & ~n1788 ;
  assign n1790 = ~n1783 & n1788 ;
  assign n1791 = n1789 | n1790 ;
  assign n1792 = n1222 | n1232 ;
  assign n1793 = n1222 & ~n1230 ;
  assign n1794 = n1792 & ~n1793 ;
  assign n1795 = ( n1115 & n1280 ) | ( n1115 & ~n1794 ) | ( n1280 & ~n1794 );
  assign n1796 = ( n1115 & ~n1282 ) | ( n1115 & n1794 ) | ( ~n1282 & n1794 );
  assign n1797 = ~n1795 & n1796 ;
  assign n1798 = n1191 & ~n1340 ;
  assign n1799 = n1129 & n1340 ;
  assign n1800 = n1798 | n1799 ;
  assign n1801 = ( n1130 & n1275 ) | ( n1130 & ~n1800 ) | ( n1275 & ~n1800 );
  assign n1802 = ( n1190 & n1275 ) | ( n1190 & n1800 ) | ( n1275 & n1800 );
  assign n1803 = n1801 & ~n1802 ;
  assign n1804 = ( ~n1791 & n1797 ) | ( ~n1791 & n1803 ) | ( n1797 & n1803 );
  assign n1805 = ( n1797 & n1803 ) | ( n1797 & ~n1804 ) | ( n1803 & ~n1804 );
  assign n1806 = ( n1791 & n1804 ) | ( n1791 & ~n1805 ) | ( n1804 & ~n1805 );
  assign n1807 = n1232 | n1275 ;
  assign n1808 = ~n1230 & n1275 ;
  assign n1809 = n1807 & ~n1808 ;
  assign n1810 = ( n1222 & n1280 ) | ( n1222 & ~n1809 ) | ( n1280 & ~n1809 );
  assign n1811 = ( n1222 & ~n1282 ) | ( n1222 & n1809 ) | ( ~n1282 & n1809 );
  assign n1812 = ~n1810 & n1811 ;
  assign n1813 = n1280 & n1340 ;
  assign n1814 = n1282 & n1340 ;
  assign n1815 = ( n1110 & ~n1813 ) | ( n1110 & n1814 ) | ( ~n1813 & n1814 );
  assign n1816 = n1115 & ~n1380 ;
  assign n1817 = n1222 & n1380 ;
  assign n1818 = ( n1058 & ~n1816 ) | ( n1058 & n1817 ) | ( ~n1816 & n1817 );
  assign n1819 = ~n1468 & n1816 ;
  assign n1820 = n1818 | n1819 ;
  assign n1821 = n1110 & ~n1820 ;
  assign n1822 = n1815 & n1821 ;
  assign n1823 = ~n828 & n1468 ;
  assign n1824 = n1058 | n1115 ;
  assign n1825 = n1380 & n1824 ;
  assign n1826 = n1823 | n1825 ;
  assign n1827 = n828 & ~n1380 ;
  assign n1828 = ~n1468 & n1827 ;
  assign n1829 = n1826 | n1828 ;
  assign n1830 = ( n1812 & n1822 ) | ( n1812 & ~n1829 ) | ( n1822 & ~n1829 );
  assign n1831 = ( n1812 & ~n1822 ) | ( n1812 & n1829 ) | ( ~n1822 & n1829 );
  assign n1832 = ( ~n1812 & n1830 ) | ( ~n1812 & n1831 ) | ( n1830 & n1831 );
  assign n1833 = ~n1110 & n1820 ;
  assign n1834 = ( ~n1815 & n1820 ) | ( ~n1815 & n1833 ) | ( n1820 & n1833 );
  assign n1835 = n1822 | n1834 ;
  assign n1843 = ~n1128 & n1340 ;
  assign n1836 = n1058 | n1275 ;
  assign n1837 = n1380 & n1836 ;
  assign n1838 = ( n1222 & ~n1469 ) | ( n1222 & n1837 ) | ( ~n1469 & n1837 );
  assign n1839 = ( ~n1222 & n1468 ) | ( ~n1222 & n1837 ) | ( n1468 & n1837 );
  assign n1840 = n1838 | n1839 ;
  assign n1841 = ( ~n1058 & n1227 ) | ( ~n1058 & n1340 ) | ( n1227 & n1340 );
  assign n1842 = ( n1108 & n1227 ) | ( n1108 & n1841 ) | ( n1227 & n1841 );
  assign n1844 = n1842 | n1843 ;
  assign n1845 = n1058 | n1340 ;
  assign n1846 = n1275 & ~n1380 ;
  assign n1847 = n1845 | n1846 ;
  assign n1848 = ~n1843 & n1847 ;
  assign n1849 = ( n1840 & ~n1844 ) | ( n1840 & n1848 ) | ( ~n1844 & n1848 );
  assign n1850 = ( n1835 & ~n1843 ) | ( n1835 & n1849 ) | ( ~n1843 & n1849 );
  assign n1851 = n1832 | n1850 ;
  assign n1852 = ~n1230 & n1340 ;
  assign n1853 = ( n1275 & n1280 ) | ( n1275 & n1852 ) | ( n1280 & n1852 );
  assign n1854 = ( ~n1275 & n1282 ) | ( ~n1275 & n1852 ) | ( n1282 & n1852 );
  assign n1855 = n1853 | n1854 ;
  assign n1856 = n1232 | n1340 ;
  assign n1857 = ~n1855 & n1856 ;
  assign n1858 = ( n1840 & ~n1842 ) | ( n1840 & n1847 ) | ( ~n1842 & n1847 );
  assign n1859 = n1856 & ~n1858 ;
  assign n1860 = ~n1855 & n1859 ;
  assign n1861 = ( ~n1835 & n1857 ) | ( ~n1835 & n1860 ) | ( n1857 & n1860 );
  assign n1862 = ( n1832 & n1851 ) | ( n1832 & ~n1861 ) | ( n1851 & ~n1861 );
  assign n1863 = ( n1835 & ~n1857 ) | ( n1835 & n1858 ) | ( ~n1857 & n1858 );
  assign n1864 = n1843 & ~n1863 ;
  assign n1865 = ~n1806 & n1864 ;
  assign n1866 = ( n1806 & n1862 ) | ( n1806 & ~n1865 ) | ( n1862 & ~n1865 );
  assign n1867 = ~n738 & n1746 ;
  assign n1868 = ( n738 & n1745 ) | ( n738 & ~n1867 ) | ( n1745 & ~n1867 );
  assign n1869 = ~n1748 & n1868 ;
  assign n1870 = ( n1789 & ~n1791 ) | ( n1789 & n1869 ) | ( ~n1791 & n1869 );
  assign n1871 = ( n1789 & n1803 ) | ( n1789 & n1869 ) | ( n1803 & n1869 );
  assign n1872 = ( n1797 & n1870 ) | ( n1797 & n1871 ) | ( n1870 & n1871 );
  assign n1873 = ( n1804 & n1869 ) | ( n1804 & ~n1872 ) | ( n1869 & ~n1872 );
  assign n1874 = ( n1789 & ~n1872 ) | ( n1789 & n1873 ) | ( ~n1872 & n1873 );
  assign n1875 = n1866 & ~n1874 ;
  assign n1876 = ~n746 & n1468 ;
  assign n1877 = n1380 & n1786 ;
  assign n1878 = n1876 | n1877 ;
  assign n1879 = n746 & ~n1380 ;
  assign n1880 = ~n1468 & n1879 ;
  assign n1881 = n1878 | n1880 ;
  assign n1882 = n1115 | n1232 ;
  assign n1883 = n1115 & ~n1230 ;
  assign n1884 = n1882 & ~n1883 ;
  assign n1885 = ( n828 & n1280 ) | ( n828 & ~n1884 ) | ( n1280 & ~n1884 );
  assign n1886 = ( n828 & ~n1282 ) | ( n828 & n1884 ) | ( ~n1282 & n1884 );
  assign n1887 = ~n1885 & n1886 ;
  assign n1888 = n1191 & ~n1275 ;
  assign n1889 = n1129 & n1275 ;
  assign n1890 = n1888 | n1889 ;
  assign n1891 = ( n1130 & n1222 ) | ( n1130 & ~n1890 ) | ( n1222 & ~n1890 );
  assign n1892 = ( n1190 & n1222 ) | ( n1190 & n1890 ) | ( n1222 & n1890 );
  assign n1893 = n1891 & ~n1892 ;
  assign n1894 = ( ~n1881 & n1887 ) | ( ~n1881 & n1893 ) | ( n1887 & n1893 );
  assign n1895 = ( n1887 & n1893 ) | ( n1887 & ~n1894 ) | ( n1893 & ~n1894 );
  assign n1896 = ( n1881 & n1894 ) | ( n1881 & ~n1895 ) | ( n1894 & ~n1895 );
  assign n1897 = n1806 & ~n1864 ;
  assign n1898 = n1830 & ~n1832 ;
  assign n1899 = n1830 & n1861 ;
  assign n1900 = ( ~n1851 & n1898 ) | ( ~n1851 & n1899 ) | ( n1898 & n1899 );
  assign n1901 = ( n1830 & ~n1897 ) | ( n1830 & n1900 ) | ( ~n1897 & n1900 );
  assign n1902 = ~n1896 & n1901 ;
  assign n1903 = ( n1875 & n1896 ) | ( n1875 & ~n1902 ) | ( n1896 & ~n1902 );
  assign n1904 = ~n1866 & n1874 ;
  assign n1905 = n1872 | n1901 ;
  assign n1906 = n1872 | n1874 ;
  assign n1907 = ( n1904 & n1905 ) | ( n1904 & n1906 ) | ( n1905 & n1906 );
  assign n1908 = n1903 & ~n1907 ;
  assign n1909 = ~n1748 & n1752 ;
  assign n1910 = n1753 | n1909 ;
  assign n1911 = ~n1893 & n1910 ;
  assign n1912 = n1881 & n1910 ;
  assign n1913 = ( ~n1887 & n1911 ) | ( ~n1887 & n1912 ) | ( n1911 & n1912 );
  assign n1914 = n1910 & ~n1912 ;
  assign n1915 = n1910 & ~n1911 ;
  assign n1916 = ( n1887 & n1914 ) | ( n1887 & n1915 ) | ( n1914 & n1915 );
  assign n1917 = ( n1894 & n1913 ) | ( n1894 & ~n1916 ) | ( n1913 & ~n1916 );
  assign n1918 = ( ~n1780 & n1908 ) | ( ~n1780 & n1917 ) | ( n1908 & n1917 );
  assign n1919 = n1756 | n1759 ;
  assign n1920 = n1736 & ~n1919 ;
  assign n1921 = n1761 | n1920 ;
  assign n1922 = n1872 & n1901 ;
  assign n1923 = n1872 & n1874 ;
  assign n1924 = ( n1904 & n1922 ) | ( n1904 & n1923 ) | ( n1922 & n1923 );
  assign n1925 = ( n1872 & ~n1903 ) | ( n1872 & n1924 ) | ( ~n1903 & n1924 );
  assign n1926 = ( n1778 & n1894 ) | ( n1778 & ~n1910 ) | ( n1894 & ~n1910 );
  assign n1927 = ( n1730 & n1893 ) | ( n1730 & ~n1910 ) | ( n1893 & ~n1910 );
  assign n1928 = ( ~n1730 & n1881 ) | ( ~n1730 & n1910 ) | ( n1881 & n1910 );
  assign n1929 = ( n1887 & n1927 ) | ( n1887 & ~n1928 ) | ( n1927 & ~n1928 );
  assign n1930 = ( ~n1779 & n1926 ) | ( ~n1779 & n1929 ) | ( n1926 & n1929 );
  assign n1931 = ( ~n1921 & n1925 ) | ( ~n1921 & n1930 ) | ( n1925 & n1930 );
  assign n1932 = n1780 & ~n1917 ;
  assign n1933 = ( n1921 & ~n1930 ) | ( n1921 & n1932 ) | ( ~n1930 & n1932 );
  assign n1934 = ( n1918 & ~n1931 ) | ( n1918 & n1933 ) | ( ~n1931 & n1933 );
  assign n1935 = ( ~n1762 & n1777 ) | ( ~n1762 & n1934 ) | ( n1777 & n1934 );
  assign n1936 = n1768 | n1776 ;
  assign n1937 = ~n1935 & n1936 ;
  assign n1938 = n1671 & ~n1937 ;
  assign n1939 = n1701 | n1937 ;
  assign n1940 = ( n1708 & ~n1938 ) | ( n1708 & n1939 ) | ( ~n1938 & n1939 );
  assign n1941 = n1701 | n1936 ;
  assign n1942 = n1935 & ~n1941 ;
  assign n1943 = n1671 & ~n1936 ;
  assign n1944 = n1935 & n1943 ;
  assign n1945 = ( ~n1708 & n1942 ) | ( ~n1708 & n1944 ) | ( n1942 & n1944 );
  assign n1946 = ( n1711 & ~n1940 ) | ( n1711 & n1945 ) | ( ~n1940 & n1945 );
  assign n1947 = ( ~n1657 & n1667 ) | ( ~n1657 & n1946 ) | ( n1667 & n1946 );
  assign n1948 = ~n1671 & n1936 ;
  assign n1949 = n1701 & n1936 ;
  assign n1950 = ( n1708 & n1948 ) | ( n1708 & n1949 ) | ( n1948 & n1949 );
  assign n1951 = n1671 | n1935 ;
  assign n1952 = n1701 & ~n1935 ;
  assign n1953 = ( n1708 & ~n1951 ) | ( n1708 & n1952 ) | ( ~n1951 & n1952 );
  assign n1954 = ( ~n1711 & n1950 ) | ( ~n1711 & n1953 ) | ( n1950 & n1953 );
  assign n1955 = ( n1668 & n1947 ) | ( n1668 & ~n1954 ) | ( n1947 & ~n1954 );
  assign n1956 = ~n1662 & n1955 ;
  assign n1957 = ( ~n1662 & n1664 ) | ( ~n1662 & n1956 ) | ( n1664 & n1956 );
  assign n1958 = n1566 & ~n1617 ;
  assign n1959 = n1618 | n1958 ;
  assign n1960 = ~n1618 & n1959 ;
  assign n1961 = ( ~n1618 & n1957 ) | ( ~n1618 & n1960 ) | ( n1957 & n1960 );
  assign n1962 = ( n1528 & ~n1564 ) | ( n1528 & n1961 ) | ( ~n1564 & n1961 );
  assign n1963 = ~n1522 & n1962 ;
  assign n1964 = ( ~n1522 & n1524 ) | ( ~n1522 & n1963 ) | ( n1524 & n1963 );
  assign n1965 = ( n1452 & ~n1455 ) | ( n1452 & n1964 ) | ( ~n1455 & n1964 );
  assign n1966 = ~n1166 & n1965 ;
  assign n1967 = n994 | n1966 ;
  assign n1968 = ~n992 & n1967 ;
  assign n1969 = n813 | n1968 ;
  assign n1970 = ~n811 & n1969 ;
  assign n1971 = ~n634 & n636 ;
  assign n1972 = n637 | n1971 ;
  assign n1973 = n1970 | n1972 ;
  assign n1974 = ~n637 & n1973 ;
  assign n1975 = n266 | n332 ;
  assign n1976 = n266 & n332 ;
  assign n1977 = n1975 & ~n1976 ;
  assign n1978 = n430 & ~n1977 ;
  assign n1979 = ~n430 & n1977 ;
  assign n1980 = n1978 | n1979 ;
  assign n1981 = n327 & ~n1980 ;
  assign n1982 = ~n1974 & n1981 ;
  assign n1983 = n637 | n1981 ;
  assign n1984 = n1973 & ~n1983 ;
  assign n1985 = n1982 | n1984 ;
  assign n1986 = ~n594 & n1985 ;
  assign n1987 = n594 & ~n1984 ;
  assign n1988 = ~n1982 & n1987 ;
  assign n1989 = n1986 | n1988 ;
  assign n1990 = n322 | n376 ;
  assign n1991 = n196 | n309 ;
  assign n1992 = n1990 | n1991 ;
  assign n1993 = n159 | n537 ;
  assign n1994 = n1992 | n1993 ;
  assign n1995 = n178 | n311 ;
  assign n1996 = n165 | n1995 ;
  assign n1997 = n398 | n1996 ;
  assign n1998 = n276 | n1997 ;
  assign n1999 = n129 | n664 ;
  assign n2000 = n137 | n144 ;
  assign n2001 = n368 | n1079 ;
  assign n2002 = n111 | n334 ;
  assign n2003 = n355 | n367 ;
  assign n2004 = n2002 | n2003 ;
  assign n2005 = n529 | n2004 ;
  assign n2006 = n2001 | n2005 ;
  assign n2007 = n164 | n459 ;
  assign n2008 = n140 | n2007 ;
  assign n2009 = n113 | n2008 ;
  assign n2010 = n225 | n2009 ;
  assign n2011 = n2006 | n2010 ;
  assign n2012 = n2000 | n2011 ;
  assign n2013 = n305 | n2012 ;
  assign n2014 = n354 | n2013 ;
  assign n2015 = n1999 | n2014 ;
  assign n2016 = n202 | n2015 ;
  assign n2017 = n1998 | n2016 ;
  assign n2018 = n560 | n2017 ;
  assign n2019 = n878 & ~n2018 ;
  assign n2020 = ~n1994 & n2019 ;
  assign n2021 = ~n836 & n2020 ;
  assign n2022 = n153 | n1036 ;
  assign n2023 = n112 | n2022 ;
  assign n2024 = n2021 & ~n2023 ;
  assign n2025 = n1989 & n2024 ;
  assign n2026 = n112 | n365 ;
  assign n2027 = n234 | n2026 ;
  assign n2028 = n123 | n704 ;
  assign n2029 = n281 | n2028 ;
  assign n2030 = n350 | n2029 ;
  assign n2031 = n413 | n2030 ;
  assign n2032 = n115 | n2031 ;
  assign n2033 = n486 | n2032 ;
  assign n2034 = n133 | n715 ;
  assign n2035 = n310 | n2034 ;
  assign n2036 = n2033 | n2035 ;
  assign n2037 = n690 | n2036 ;
  assign n2038 = n120 | n410 ;
  assign n2039 = n144 | n2038 ;
  assign n2040 = n288 | n556 ;
  assign n2041 = n368 | n2040 ;
  assign n2042 = n338 | n2041 ;
  assign n2043 = n374 | n488 ;
  assign n2044 = n200 | n414 ;
  assign n2045 = n142 | n2044 ;
  assign n2046 = n908 | n1041 ;
  assign n2047 = n2045 | n2046 ;
  assign n2048 = n2043 | n2047 ;
  assign n2049 = n2042 | n2048 ;
  assign n2050 = n2039 | n2049 ;
  assign n2051 = n195 | n376 ;
  assign n2052 = n401 | n537 ;
  assign n2053 = n2051 | n2052 ;
  assign n2054 = n370 | n2053 ;
  assign n2055 = n222 | n2054 ;
  assign n2056 = n668 | n2055 ;
  assign n2057 = n158 | n233 ;
  assign n2058 = n152 | n2057 ;
  assign n2059 = n2056 | n2058 ;
  assign n2060 = n180 | n475 ;
  assign n2061 = n641 | n2060 ;
  assign n2062 = n2059 | n2061 ;
  assign n2063 = n2050 | n2062 ;
  assign n2064 = n2037 | n2063 ;
  assign n2065 = n2027 | n2064 ;
  assign n2066 = n322 | n2065 ;
  assign n2067 = n219 | n2066 ;
  assign n2068 = n167 | n2067 ;
  assign n2069 = n417 | n2068 ;
  assign n2070 = n367 | n2069 ;
  assign n2071 = n237 | n2070 ;
  assign n2072 = n1970 & n1972 ;
  assign n2073 = n1973 & ~n2072 ;
  assign n2074 = n2071 & ~n2073 ;
  assign n2075 = n523 | n643 ;
  assign n2076 = n697 | n844 ;
  assign n2077 = n831 | n2076 ;
  assign n2078 = n369 | n2077 ;
  assign n2079 = n2075 | n2078 ;
  assign n2080 = n900 | n901 ;
  assign n2081 = n2079 | n2080 ;
  assign n2082 = n536 | n2081 ;
  assign n2083 = n1051 | n2082 ;
  assign n2084 = n350 | n2083 ;
  assign n2085 = n338 | n2084 ;
  assign n2086 = n401 | n2085 ;
  assign n2087 = n159 | n2086 ;
  assign n2088 = n214 | n2087 ;
  assign n2089 = n813 & n1968 ;
  assign n2090 = n1969 & ~n2089 ;
  assign n2091 = n2088 & ~n2090 ;
  assign n2092 = n994 & n1966 ;
  assign n2093 = n1967 & ~n2092 ;
  assign n2094 = n152 | n209 ;
  assign n2095 = n213 | n717 ;
  assign n2096 = n221 | n268 ;
  assign n2097 = n459 | n2096 ;
  assign n2098 = n2095 | n2097 ;
  assign n2099 = n523 | n2027 ;
  assign n2100 = n196 | n1990 ;
  assign n2101 = n2045 | n2100 ;
  assign n2102 = n2099 | n2101 ;
  assign n2103 = n2098 | n2102 ;
  assign n2104 = n2094 | n2103 ;
  assign n2105 = n382 | n412 ;
  assign n2106 = n168 | n2105 ;
  assign n2107 = n507 | n2106 ;
  assign n2108 = n372 | n2000 ;
  assign n2109 = n2107 | n2108 ;
  assign n2110 = n276 | n487 ;
  assign n2111 = n267 | n2110 ;
  assign n2112 = n195 | n845 ;
  assign n2113 = n336 | n2112 ;
  assign n2114 = n115 | n2113 ;
  assign n2115 = n94 | n2114 ;
  assign n2116 = n215 | n2115 ;
  assign n2117 = n469 | n558 ;
  assign n2118 = n2116 | n2117 ;
  assign n2119 = n218 | n2118 ;
  assign n2120 = n272 | n2119 ;
  assign n2121 = n107 | n2120 ;
  assign n2122 = n641 | n2121 ;
  assign n2123 = n2111 | n2122 ;
  assign n2124 = n307 | n333 ;
  assign n2125 = n411 | n2124 ;
  assign n2126 = n465 | n2125 ;
  assign n2127 = n2123 | n2126 ;
  assign n2128 = n2109 | n2127 ;
  assign n2129 = n2104 | n2128 ;
  assign n2130 = ~n2093 & n2129 ;
  assign n2131 = n2093 & ~n2129 ;
  assign n2132 = n2130 | n2131 ;
  assign n2133 = n336 | n485 ;
  assign n2134 = n214 | n2133 ;
  assign n2135 = n237 | n386 ;
  assign n2136 = n132 | n2135 ;
  assign n2137 = n2104 | n2136 ;
  assign n2138 = n402 | n2137 ;
  assign n2139 = n1361 | n2138 ;
  assign n2140 = n2134 | n2139 ;
  assign n2141 = n312 | n2106 ;
  assign n2142 = n341 | n2141 ;
  assign n2143 = n122 | n2142 ;
  assign n2144 = n178 | n2143 ;
  assign n2145 = n203 | n2144 ;
  assign n2146 = n405 | n2145 ;
  assign n2147 = n398 | n2146 ;
  assign n2148 = n367 | n2147 ;
  assign n2149 = n567 | n2148 ;
  assign n2150 = n878 & ~n2033 ;
  assign n2151 = ~n2149 & n2150 ;
  assign n2152 = ~n2140 & n2151 ;
  assign n2153 = n166 | n910 ;
  assign n2154 = n2152 & ~n2153 ;
  assign n2155 = ~n344 & n2154 ;
  assign n2156 = ~n158 & n2155 ;
  assign n2157 = ~n356 & n2156 ;
  assign n2158 = ~n307 & n2157 ;
  assign n2159 = ~n1444 & n1446 ;
  assign n2160 = ( n1448 & n1454 ) | ( n1448 & ~n2159 ) | ( n1454 & ~n2159 );
  assign n2161 = n1435 & ~n2160 ;
  assign n2162 = ( n1431 & ~n1448 ) | ( n1431 & n2159 ) | ( ~n1448 & n2159 );
  assign n2163 = n1435 & n2162 ;
  assign n2164 = ( n1964 & n2161 ) | ( n1964 & n2163 ) | ( n2161 & n2163 );
  assign n2165 = n1965 & ~n2164 ;
  assign n2166 = n2158 | n2165 ;
  assign n2167 = n2158 & n2165 ;
  assign n2168 = n136 | n218 ;
  assign n2169 = n107 | n2168 ;
  assign n2170 = n162 | n2169 ;
  assign n2171 = n211 | n2170 ;
  assign n2172 = n413 | n2171 ;
  assign n2173 = n239 | n2172 ;
  assign n2174 = n159 | n2173 ;
  assign n2175 = n124 | n1020 ;
  assign n2176 = n507 | n2175 ;
  assign n2177 = n2002 | n2176 ;
  assign n2178 = n876 | n2177 ;
  assign n2179 = n311 | n350 ;
  assign n2180 = n2178 | n2179 ;
  assign n2181 = n336 | n2180 ;
  assign n2182 = n352 | n2181 ;
  assign n2183 = n89 | n856 ;
  assign n2184 = n537 | n2183 ;
  assign n2185 = n219 | n238 ;
  assign n2186 = n113 | n2185 ;
  assign n2187 = n204 | n2186 ;
  assign n2188 = n366 | n2187 ;
  assign n2189 = n2184 | n2188 ;
  assign n2190 = n2182 | n2189 ;
  assign n2191 = n2174 | n2190 ;
  assign n2192 = n322 | n2191 ;
  assign n2193 = n282 | n2192 ;
  assign n2194 = n182 | n2193 ;
  assign n2195 = n234 | n2194 ;
  assign n2196 = n410 | n2195 ;
  assign n2197 = n340 | n2196 ;
  assign n2198 = n333 | n2197 ;
  assign n2199 = n1322 & ~n1446 ;
  assign n2200 = ( n1431 & n1446 ) | ( n1431 & ~n2199 ) | ( n1446 & ~n2199 );
  assign n2201 = ( ~n1446 & n1454 ) | ( ~n1446 & n2199 ) | ( n1454 & n2199 );
  assign n2202 = ( n1964 & n2200 ) | ( n1964 & ~n2201 ) | ( n2200 & ~n2201 );
  assign n2203 = ~n1322 & n1446 ;
  assign n2204 = ~n1454 & n2203 ;
  assign n2205 = n1431 & n2203 ;
  assign n2206 = ( n1964 & n2204 ) | ( n1964 & n2205 ) | ( n2204 & n2205 );
  assign n2207 = n2202 & ~n2206 ;
  assign n2208 = n2198 & ~n2207 ;
  assign n2209 = n206 | n416 ;
  assign n2210 = n641 | n664 ;
  assign n2211 = n2209 | n2210 ;
  assign n2212 = n863 | n2211 ;
  assign n2213 = n132 | n2212 ;
  assign n2214 = n918 | n920 ;
  assign n2215 = n97 | n537 ;
  assign n2216 = n837 | n857 ;
  assign n2217 = n677 | n2216 ;
  assign n2218 = n160 | n2217 ;
  assign n2219 = ( n366 & ~n2215 ) | ( n366 & n2218 ) | ( ~n2215 & n2218 );
  assign n2220 = n2215 | n2219 ;
  assign n2221 = n113 | n136 ;
  assign n2222 = n89 | n353 ;
  assign n2223 = n215 | n2222 ;
  assign n2224 = n544 | n2223 ;
  assign n2225 = n2221 | n2224 ;
  assign n2226 = n1017 | n2225 ;
  assign n2227 = n560 | n2226 ;
  assign n2228 = n308 | n2227 ;
  assign n2229 = n2220 | n2228 ;
  assign n2230 = n2214 | n2229 ;
  assign n2231 = n2213 | n2230 ;
  assign n2232 = n238 | n397 ;
  assign n2233 = n2231 | n2232 ;
  assign n2234 = ( n1431 & ~n1454 ) | ( n1431 & n1964 ) | ( ~n1454 & n1964 );
  assign n2235 = n1323 & ~n1429 ;
  assign n2236 = n1323 & n1326 ;
  assign n2237 = ( n1964 & n2235 ) | ( n1964 & n2236 ) | ( n2235 & n2236 );
  assign n2238 = n2234 & ~n2237 ;
  assign n2239 = n2233 & ~n2238 ;
  assign n2240 = ~n2233 & n2238 ;
  assign n2241 = n196 | n339 ;
  assign n2242 = n487 | n2241 ;
  assign n2243 = n182 | n214 ;
  assign n2244 = n2242 | n2243 ;
  assign n2245 = n178 | n849 ;
  assign n2246 = n2244 | n2245 ;
  assign n2247 = n309 | n353 ;
  assign n2248 = n186 | n376 ;
  assign n2249 = n2247 | n2248 ;
  assign n2250 = n409 | n2249 ;
  assign n2251 = n2246 | n2250 ;
  assign n2252 = n124 | n298 ;
  assign n2253 = n272 | n307 ;
  assign n2254 = n2252 | n2253 ;
  assign n2255 = n226 | n486 ;
  assign n2256 = n212 | n2255 ;
  assign n2257 = n2254 | n2256 ;
  assign n2258 = n337 | n2013 ;
  assign n2259 = n2038 | n2258 ;
  assign n2260 = n2257 | n2259 ;
  assign n2261 = n2251 | n2260 ;
  assign n2262 = n184 | n209 ;
  assign n2263 = n268 | n2262 ;
  assign n2264 = n158 | n2263 ;
  assign n2265 = n352 | n2264 ;
  assign n2266 = n2261 | n2265 ;
  assign n2267 = n383 | n2266 ;
  assign n2268 = ( n1326 & ~n1429 ) | ( n1326 & n1964 ) | ( ~n1429 & n1964 );
  assign n2269 = ( n1326 & n1964 ) | ( n1326 & ~n2268 ) | ( n1964 & ~n2268 );
  assign n2270 = ( n1429 & n2268 ) | ( n1429 & ~n2269 ) | ( n2268 & ~n2269 );
  assign n2271 = n2267 & ~n2270 ;
  assign n2272 = n201 | n487 ;
  assign n2273 = n370 | n2272 ;
  assign n2274 = n211 | n234 ;
  assign n2275 = n908 | n2274 ;
  assign n2276 = n116 | n2275 ;
  assign n2277 = n2273 | n2276 ;
  assign n2278 = n289 | n377 ;
  assign n2279 = n410 | n2278 ;
  assign n2280 = n102 | n2279 ;
  assign n2281 = n226 | n2280 ;
  assign n2282 = n367 | n2281 ;
  assign n2283 = n476 | n2282 ;
  assign n2284 = n845 | n2125 ;
  assign n2285 = n495 | n2284 ;
  assign n2286 = n284 | n2285 ;
  assign n2287 = n356 | n2286 ;
  assign n2288 = n2215 | n2287 ;
  assign n2289 = n225 | n2288 ;
  assign n2290 = n2283 | n2289 ;
  assign n2291 = n646 | n2290 ;
  assign n2292 = n222 | n653 ;
  assign n2293 = n276 | n639 ;
  assign n2294 = n2292 | n2293 ;
  assign n2295 = n2291 | n2294 ;
  assign n2296 = n2277 | n2295 ;
  assign n2297 = n386 | n2296 ;
  assign n2298 = n219 | n2297 ;
  assign n2299 = n1524 | n1962 ;
  assign n2300 = n1524 & n1962 ;
  assign n2301 = n2299 & ~n2300 ;
  assign n2302 = n2298 & ~n2301 ;
  assign n2303 = n417 | n455 ;
  assign n2304 = n312 | n727 ;
  assign n2305 = n2303 | n2304 ;
  assign n2306 = n2282 | n2305 ;
  assign n2307 = n878 & ~n2306 ;
  assign n2308 = ~n836 & n2307 ;
  assign n2309 = ~n913 & n2308 ;
  assign n2310 = n371 | n398 ;
  assign n2311 = n94 | n1345 ;
  assign n2312 = n2310 | n2311 ;
  assign n2313 = n339 | n386 ;
  assign n2314 = n930 | n2313 ;
  assign n2315 = n2312 | n2314 ;
  assign n2316 = n2134 | n2315 ;
  assign n2317 = n529 | n2316 ;
  assign n2318 = n867 | n2317 ;
  assign n2319 = n405 | n2318 ;
  assign n2320 = n2211 | n2319 ;
  assign n2321 = n383 | n401 ;
  assign n2322 = n225 | n2321 ;
  assign n2323 = n2320 | n2322 ;
  assign n2324 = n2309 & ~n2323 ;
  assign n2325 = ~n148 & n2324 ;
  assign n2326 = ~n322 & n2325 ;
  assign n2327 = ~n207 & n2326 ;
  assign n2328 = ~n200 & n2327 ;
  assign n2329 = ~n356 & n2328 ;
  assign n2330 = ~n215 & n2329 ;
  assign n2331 = ( ~n1528 & n1564 ) | ( ~n1528 & n1961 ) | ( n1564 & n1961 );
  assign n2332 = ( n1564 & n1961 ) | ( n1564 & ~n2331 ) | ( n1961 & ~n2331 );
  assign n2333 = ( n1528 & n2331 ) | ( n1528 & ~n2332 ) | ( n2331 & ~n2332 );
  assign n2334 = n2330 | n2333 ;
  assign n2335 = n2330 & n2333 ;
  assign n2336 = n144 | n485 ;
  assign n2337 = n197 | n2313 ;
  assign n2338 = n369 | n2337 ;
  assign n2339 = n166 | n298 ;
  assign n2340 = n355 | n2339 ;
  assign n2341 = n414 | n2340 ;
  assign n2342 = n120 | n2341 ;
  assign n2343 = n352 | n487 ;
  assign n2344 = n2342 | n2343 ;
  assign n2345 = n2338 | n2344 ;
  assign n2346 = n132 | n218 ;
  assign n2347 = n1021 | n2346 ;
  assign n2348 = n344 | n350 ;
  assign n2349 = n405 | n2348 ;
  assign n2350 = n2220 | n2349 ;
  assign n2351 = n2347 | n2350 ;
  assign n2352 = n2345 | n2351 ;
  assign n2353 = n2336 | n2352 ;
  assign n2354 = n713 | n2353 ;
  assign n2355 = n371 | n2354 ;
  assign n2356 = n153 | n311 ;
  assign n2357 = n2355 | n2356 ;
  assign n2358 = n112 | n187 ;
  assign n2359 = n107 | n2358 ;
  assign n2360 = n2357 | n2359 ;
  assign n2361 = n226 | n413 ;
  assign n2362 = n333 | n2361 ;
  assign n2363 = n2360 | n2362 ;
  assign n2364 = n1957 | n1959 ;
  assign n2365 = n1957 & n1959 ;
  assign n2366 = n2364 & ~n2365 ;
  assign n2367 = n2363 & ~n2366 ;
  assign n2368 = ~n2363 & n2366 ;
  assign n2369 = n657 | n1039 ;
  assign n2370 = n664 | n2369 ;
  assign n2371 = n529 | n2370 ;
  assign n2372 = n840 | n2371 ;
  assign n2373 = n2289 | n2372 ;
  assign n2374 = n643 | n2050 ;
  assign n2375 = n272 | n2374 ;
  assign n2376 = n2373 | n2375 ;
  assign n2377 = n187 | n401 ;
  assign n2378 = n180 | n2377 ;
  assign n2379 = n567 | n2378 ;
  assign n2380 = n2376 | n2379 ;
  assign n2381 = n1664 | n1955 ;
  assign n2382 = n1664 & ~n1955 ;
  assign n2383 = ( ~n1664 & n2381 ) | ( ~n1664 & n2382 ) | ( n2381 & n2382 );
  assign n2384 = ~n2380 & n2383 ;
  assign n2385 = n2367 | n2384 ;
  assign n2386 = n2368 | n2385 ;
  assign n2387 = ~n2367 & n2386 ;
  assign n2388 = n2334 & ~n2387 ;
  assign n2389 = ~n2335 & n2388 ;
  assign n2390 = n2334 & ~n2389 ;
  assign n2391 = ~n2298 & n2301 ;
  assign n2392 = n2302 | n2391 ;
  assign n2393 = n2390 | n2392 ;
  assign n2394 = ~n2302 & n2393 ;
  assign n2395 = ~n2267 & n2270 ;
  assign n2396 = n2271 | n2395 ;
  assign n2397 = n2394 | n2396 ;
  assign n2398 = ~n2271 & n2397 ;
  assign n2399 = n2239 | n2398 ;
  assign n2400 = n2240 | n2399 ;
  assign n2401 = ~n2239 & n2400 ;
  assign n2402 = n2198 & ~n2208 ;
  assign n2403 = n2207 | n2208 ;
  assign n2404 = ~n2402 & n2403 ;
  assign n2405 = n2401 | n2404 ;
  assign n2406 = ~n2208 & n2405 ;
  assign n2407 = n2166 & ~n2406 ;
  assign n2408 = ~n2167 & n2407 ;
  assign n2409 = n2166 & ~n2408 ;
  assign n2410 = n2132 | n2409 ;
  assign n2411 = ~n2130 & n2410 ;
  assign n2412 = ~n2088 & n2090 ;
  assign n2413 = n2091 | n2412 ;
  assign n2414 = n2411 | n2413 ;
  assign n2415 = ~n2091 & n2414 ;
  assign n2416 = ~n2071 & n2073 ;
  assign n2417 = n2074 | n2416 ;
  assign n2418 = n2415 | n2417 ;
  assign n2419 = ~n2074 & n2418 ;
  assign n2420 = n1988 | n2024 ;
  assign n2421 = n1986 | n2420 ;
  assign n2422 = ~n2419 & n2421 ;
  assign n2423 = ~n2025 & n2422 ;
  assign n2424 = n372 | n1041 ;
  assign n2425 = n2220 | n2424 ;
  assign n2426 = n1370 | n2425 ;
  assign n2427 = n178 | n218 ;
  assign n2428 = n164 | n2427 ;
  assign n2429 = n282 | n699 ;
  assign n2430 = n2428 | n2429 ;
  assign n2431 = n334 | n2430 ;
  assign n2432 = n2426 | n2431 ;
  assign n2433 = n514 | n2432 ;
  assign n2434 = n116 | n2433 ;
  assign n2435 = n281 | n2434 ;
  assign n2436 = n883 | n2435 ;
  assign n2437 = n485 | n2436 ;
  assign n2438 = n487 | n2437 ;
  assign n2439 = n225 | n2438 ;
  assign n2440 = n2421 & ~n2439 ;
  assign n2441 = ~n2423 & n2440 ;
  assign n2442 = n166 | n176 ;
  assign n2443 = n485 | n669 ;
  assign n2444 = n676 | n2443 ;
  assign n2445 = n2442 | n2444 ;
  assign n2446 = n218 | n670 ;
  assign n2447 = n200 | n2446 ;
  assign n2448 = n349 | n715 ;
  assign n2449 = n537 | n2448 ;
  assign n2450 = n2027 | n2449 ;
  assign n2451 = n190 | n2450 ;
  assign n2452 = n222 | n288 ;
  assign n2453 = n206 | n2452 ;
  assign n2454 = n2451 | n2453 ;
  assign n2455 = n355 | n2454 ;
  assign n2456 = n336 | n2455 ;
  assign n2457 = n398 | n2456 ;
  assign n2458 = n97 | n2457 ;
  assign n2459 = n401 | n2458 ;
  assign n2460 = n154 | n651 ;
  assign n2461 = n2459 | n2460 ;
  assign n2462 = n2447 | n2461 ;
  assign n2463 = n305 | n2242 ;
  assign n2464 = n120 | n167 ;
  assign n2465 = n2463 | n2464 ;
  assign n2466 = n178 | n212 ;
  assign n2467 = n141 | n233 ;
  assign n2468 = n2466 | n2467 ;
  assign n2469 = n2465 | n2468 ;
  assign n2470 = n144 | n219 ;
  assign n2471 = n136 | n353 ;
  assign n2472 = n2470 | n2471 ;
  assign n2473 = n149 | n370 ;
  assign n2474 = n89 | n137 ;
  assign n2475 = n2473 | n2474 ;
  assign n2476 = n2472 | n2475 ;
  assign n2477 = n2469 | n2476 ;
  assign n2478 = n2462 | n2477 ;
  assign n2479 = n2445 | n2478 ;
  assign n2480 = n414 | n2479 ;
  assign n2481 = n129 | n208 ;
  assign n2482 = n335 | n371 ;
  assign n2483 = n2481 | n2482 ;
  assign n2484 = n2480 | n2483 ;
  assign n2485 = n2441 & ~n2484 ;
  assign n2486 = n292 | n296 ;
  assign n2487 = n112 | n2486 ;
  assign n2488 = ~n718 & n877 ;
  assign n2489 = ~n385 & n2488 ;
  assign n2490 = ~n2487 & n2489 ;
  assign n2491 = ~n2116 & n2490 ;
  assign n2492 = ~n2211 & n2491 ;
  assign n2493 = ~n1345 & n2492 ;
  assign n2494 = ~n902 & n2493 ;
  assign n2495 = ~n417 & n2494 ;
  assign n2496 = ~n338 & n2495 ;
  assign n2497 = ~n205 & n2496 ;
  assign n2498 = ~n214 & n2497 ;
  assign n2499 = ~n201 & n2498 ;
  assign n2500 = n2485 & n2499 ;
  assign n2501 = n233 | n275 ;
  assign n2502 = n354 | n2501 ;
  assign n2503 = n310 | n1082 ;
  assign n2504 = n2502 | n2503 ;
  assign n2505 = n308 | n2504 ;
  assign n2506 = n302 | n2505 ;
  assign n2507 = n112 | n279 ;
  assign n2508 = n385 | n408 ;
  assign n2509 = n343 | n2508 ;
  assign n2510 = n2507 | n2509 ;
  assign n2511 = n123 | n2510 ;
  assign n2512 = n2506 | n2511 ;
  assign n2513 = n2500 & ~n2512 ;
  assign n2514 = n115 | n353 ;
  assign n2515 = n407 | n2514 ;
  assign n2516 = n404 | n2515 ;
  assign n2517 = n424 | n2516 ;
  assign n2518 = n287 | n385 ;
  assign n2519 = n319 | n2518 ;
  assign n2520 = n2517 | n2519 ;
  assign n2521 = n178 | n234 ;
  assign n2522 = n226 | n2521 ;
  assign n2523 = n2520 | n2522 ;
  assign n2524 = ~n2513 & n2523 ;
  assign n2525 = n2513 & ~n2523 ;
  assign n2526 = n2524 | n2525 ;
  assign n2527 = pi1 & ~n257 ;
  assign n2528 = ~pi1 & n257 ;
  assign n2529 = n2527 | n2528 ;
  assign n2530 = n262 & ~n2529 ;
  assign n2531 = ~n262 & n2529 ;
  assign n2532 = n2530 | n2531 ;
  assign n2533 = pi0 & ~n2532 ;
  assign n2534 = n2526 & n2533 ;
  assign n2535 = n2485 | n2499 ;
  assign n2536 = ~n2500 & n2535 ;
  assign n2537 = ~n259 & n2532 ;
  assign n2538 = ~n2536 & n2537 ;
  assign n2539 = n2500 | n2512 ;
  assign n2540 = n2500 & n2512 ;
  assign n2541 = n2539 & ~n2540 ;
  assign n2542 = ~pi0 & n2529 ;
  assign n2543 = n2541 & n2542 ;
  assign n2544 = n2538 | n2543 ;
  assign n2545 = n2534 | n2544 ;
  assign n2546 = n2526 | n2541 ;
  assign n2547 = n2526 & n2541 ;
  assign n2548 = n2546 & ~n2547 ;
  assign n2549 = n2536 & ~n2541 ;
  assign n2550 = n2421 & ~n2423 ;
  assign n2551 = n2439 & ~n2550 ;
  assign n2552 = n2441 | n2551 ;
  assign n2553 = ~n2025 & n2421 ;
  assign n2554 = n2419 & ~n2553 ;
  assign n2555 = n2423 | n2554 ;
  assign n2556 = n2552 & ~n2555 ;
  assign n2557 = n2415 & n2417 ;
  assign n2558 = n2418 & ~n2557 ;
  assign n2559 = ~n2555 & n2558 ;
  assign n2560 = n2555 & ~n2558 ;
  assign n2561 = n2559 | n2560 ;
  assign n2562 = n2411 & n2413 ;
  assign n2563 = n2414 & ~n2562 ;
  assign n2564 = n2558 & n2563 ;
  assign n2565 = n2132 & n2409 ;
  assign n2566 = n2410 & ~n2565 ;
  assign n2567 = n2563 & n2566 ;
  assign n2568 = n2558 | n2563 ;
  assign n2569 = ~n2564 & n2568 ;
  assign n2570 = ~n2167 & n2409 ;
  assign n2571 = n2406 | n2408 ;
  assign n2572 = ~n2570 & n2571 ;
  assign n2573 = ~n2401 & n2405 ;
  assign n2574 = ~n2404 & n2405 ;
  assign n2575 = n2573 | n2574 ;
  assign n2576 = ~n2572 & n2575 ;
  assign n2577 = ~n2398 & n2400 ;
  assign n2578 = ~n2240 & n2401 ;
  assign n2579 = n2577 | n2578 ;
  assign n2580 = n2575 & n2579 ;
  assign n2581 = n2575 | n2579 ;
  assign n2582 = ~n2580 & n2581 ;
  assign n2583 = n2394 & n2396 ;
  assign n2584 = n2397 & ~n2583 ;
  assign n2585 = n2579 & n2584 ;
  assign n2586 = n2390 & n2392 ;
  assign n2587 = n2393 & ~n2586 ;
  assign n2588 = n2584 & n2587 ;
  assign n2589 = n2387 | n2389 ;
  assign n2590 = ~n2335 & n2390 ;
  assign n2591 = n2589 & ~n2590 ;
  assign n2592 = n2587 & ~n2591 ;
  assign n2593 = ~n2587 & n2591 ;
  assign n2594 = ~n2384 & n2386 ;
  assign n2595 = ~n2368 & n2387 ;
  assign n2596 = n2594 | n2595 ;
  assign n2597 = n2380 & ~n2383 ;
  assign n2598 = n2384 | n2597 ;
  assign n2599 = n2591 & ~n2598 ;
  assign n2600 = n2596 & ~n2599 ;
  assign n2601 = ~n2593 & n2600 ;
  assign n2602 = ~n2592 & n2601 ;
  assign n2603 = n2592 | n2602 ;
  assign n2604 = n2584 | n2587 ;
  assign n2605 = n2603 & n2604 ;
  assign n2606 = ~n2588 & n2605 ;
  assign n2607 = n2588 | n2606 ;
  assign n2608 = n2579 | n2584 ;
  assign n2609 = ~n2585 & n2608 ;
  assign n2610 = n2607 & n2609 ;
  assign n2611 = n2585 | n2610 ;
  assign n2612 = n2580 | n2611 ;
  assign n2613 = ( n2580 & n2582 ) | ( n2580 & n2612 ) | ( n2582 & n2612 );
  assign n2614 = n2572 & ~n2575 ;
  assign n2615 = n2576 | n2614 ;
  assign n2616 = ~n2576 & n2615 ;
  assign n2617 = ( n2576 & n2613 ) | ( n2576 & ~n2616 ) | ( n2613 & ~n2616 );
  assign n2618 = n2563 | n2566 ;
  assign n2619 = ~n2567 & n2618 ;
  assign n2620 = n2566 & ~n2572 ;
  assign n2621 = ~n2566 & n2572 ;
  assign n2622 = n2620 | n2621 ;
  assign n2623 = ~n2620 & n2622 ;
  assign n2624 = n2619 & ~n2623 ;
  assign n2625 = n2619 & n2620 ;
  assign n2626 = ( n2617 & n2624 ) | ( n2617 & n2625 ) | ( n2624 & n2625 );
  assign n2627 = ( n2567 & n2569 ) | ( n2567 & n2626 ) | ( n2569 & n2626 );
  assign n2628 = n2564 | n2627 ;
  assign n2629 = n2559 | n2628 ;
  assign n2630 = ( n2559 & ~n2561 ) | ( n2559 & n2629 ) | ( ~n2561 & n2629 );
  assign n2631 = ~n2552 & n2555 ;
  assign n2632 = n2556 | n2631 ;
  assign n2633 = ~n2556 & n2632 ;
  assign n2634 = ( n2556 & n2630 ) | ( n2556 & ~n2633 ) | ( n2630 & ~n2633 );
  assign n2635 = n2441 | n2484 ;
  assign n2636 = n2441 & n2484 ;
  assign n2637 = n2635 & ~n2636 ;
  assign n2638 = ~n2536 & n2637 ;
  assign n2639 = n2536 & ~n2637 ;
  assign n2640 = n2638 | n2639 ;
  assign n2641 = n2552 & n2637 ;
  assign n2642 = n2552 | n2637 ;
  assign n2643 = ~n2641 & n2642 ;
  assign n2644 = n2641 | n2643 ;
  assign n2645 = ~n2640 & n2644 ;
  assign n2646 = ~n2640 & n2641 ;
  assign n2647 = ( n2634 & n2645 ) | ( n2634 & n2646 ) | ( n2645 & n2646 );
  assign n2648 = ( ~n2536 & n2541 ) | ( ~n2536 & n2638 ) | ( n2541 & n2638 );
  assign n2649 = ( ~n2549 & n2647 ) | ( ~n2549 & n2648 ) | ( n2647 & n2648 );
  assign n2650 = n2548 | n2649 ;
  assign n2651 = n2548 & n2648 ;
  assign n2652 = n2548 & ~n2549 ;
  assign n2653 = ( n2647 & n2651 ) | ( n2647 & n2652 ) | ( n2651 & n2652 );
  assign n2654 = n2650 & ~n2653 ;
  assign n2655 = pi0 & n2532 ;
  assign n2656 = n2654 & n2655 ;
  assign n2657 = n2545 | n2656 ;
  assign n2658 = n262 | n2657 ;
  assign n2659 = n262 & n2657 ;
  assign n2660 = n2658 & ~n2659 ;
  assign n2661 = ~n746 & n949 ;
  assign n2662 = n746 & ~n949 ;
  assign n2663 = n2661 | n2662 ;
  assign n2664 = n2598 & n2663 ;
  assign n2665 = n453 & ~n2664 ;
  assign n2666 = ~n746 & n755 ;
  assign n2667 = n746 & ~n755 ;
  assign n2668 = n2666 | n2667 ;
  assign n2669 = ~n2663 & n2668 ;
  assign n2670 = n2598 & n2669 ;
  assign n2671 = n453 | n755 ;
  assign n2672 = n453 & n755 ;
  assign n2673 = n2671 & ~n2672 ;
  assign n2674 = n2663 & ~n2673 ;
  assign n2675 = n2596 & n2674 ;
  assign n2676 = n2670 | n2675 ;
  assign n2677 = ~n2596 & n2598 ;
  assign n2678 = n2596 & ~n2598 ;
  assign n2679 = n2677 | n2678 ;
  assign n2680 = n2663 & n2673 ;
  assign n2681 = n2679 & n2680 ;
  assign n2682 = n2676 | n2681 ;
  assign n2683 = n453 | n2682 ;
  assign n2684 = n453 & n2682 ;
  assign n2685 = n2683 & ~n2684 ;
  assign n2686 = n2665 & n2685 ;
  assign n2687 = n2665 | n2685 ;
  assign n2688 = ~n2686 & n2687 ;
  assign n2689 = ~n828 & n949 ;
  assign n2690 = n828 & ~n949 ;
  assign n2691 = n2689 | n2690 ;
  assign n2692 = ~n828 & n1115 ;
  assign n2693 = n828 & ~n1115 ;
  assign n2694 = n2692 | n2693 ;
  assign n2695 = n1115 & ~n1222 ;
  assign n2696 = ~n1115 & n1222 ;
  assign n2697 = n2695 | n2696 ;
  assign n2698 = n2694 | n2697 ;
  assign n2699 = n2691 & ~n2698 ;
  assign n2700 = ~n2591 & n2699 ;
  assign n2701 = n2694 & ~n2697 ;
  assign n2702 = n2587 & n2701 ;
  assign n2703 = ~n2691 & n2697 ;
  assign n2704 = n2584 & n2703 ;
  assign n2705 = n2702 | n2704 ;
  assign n2706 = n2700 | n2705 ;
  assign n2707 = n2603 & ~n2606 ;
  assign n2708 = n2604 & ~n2607 ;
  assign n2709 = n2707 | n2708 ;
  assign n2710 = n2691 & n2697 ;
  assign n2711 = n2709 & n2710 ;
  assign n2712 = n2706 | n2711 ;
  assign n2713 = n949 | n2712 ;
  assign n2714 = n949 & n2712 ;
  assign n2715 = n2713 & ~n2714 ;
  assign n2716 = n2596 & n2701 ;
  assign n2717 = n2598 & ~n2698 ;
  assign n2718 = n2691 & n2717 ;
  assign n2719 = n2716 | n2718 ;
  assign n2720 = ~n2591 & n2697 ;
  assign n2721 = ~n2691 & n2720 ;
  assign n2722 = n2719 | n2721 ;
  assign n2723 = n2591 & ~n2678 ;
  assign n2724 = ~n2591 & n2678 ;
  assign n2725 = n2723 | n2724 ;
  assign n2726 = ( n2710 & n2721 ) | ( n2710 & ~n2725 ) | ( n2721 & ~n2725 );
  assign n2727 = ~n2710 & n2725 ;
  assign n2728 = ( n2719 & n2726 ) | ( n2719 & ~n2727 ) | ( n2726 & ~n2727 );
  assign n2729 = n2722 | n2728 ;
  assign n2730 = n949 | n2729 ;
  assign n2731 = n949 & n2729 ;
  assign n2732 = n2730 & ~n2731 ;
  assign n2733 = n2598 & n2701 ;
  assign n2734 = n2596 & n2697 ;
  assign n2735 = ~n2691 & n2734 ;
  assign n2736 = n2733 | n2735 ;
  assign n2737 = n2679 & n2697 ;
  assign n2738 = n2691 & n2737 ;
  assign n2739 = n949 | n2738 ;
  assign n2740 = n2736 | n2739 ;
  assign n2741 = ~n949 & n2740 ;
  assign n2742 = n2598 & n2697 ;
  assign n2743 = n949 & ~n2742 ;
  assign n2744 = n2740 & n2743 ;
  assign n2745 = n2736 | n2738 ;
  assign n2746 = n2743 & ~n2745 ;
  assign n2747 = ( n2741 & n2744 ) | ( n2741 & n2746 ) | ( n2744 & n2746 );
  assign n2748 = n2664 & n2747 ;
  assign n2749 = n2732 & n2748 ;
  assign n2750 = n2664 & ~n2749 ;
  assign n2751 = n2600 & ~n2602 ;
  assign n2752 = n2593 | n2603 ;
  assign n2753 = ~n2751 & n2752 ;
  assign n2754 = n2710 & ~n2753 ;
  assign n2755 = ~n2591 & n2701 ;
  assign n2756 = n2587 & n2703 ;
  assign n2757 = n2596 & n2699 ;
  assign n2758 = n2756 | n2757 ;
  assign n2759 = n2755 | n2758 ;
  assign n2760 = n2754 | n2759 ;
  assign n2761 = n949 & ~n2760 ;
  assign n2762 = n949 & ~n2761 ;
  assign n2763 = ( n2760 & n2761 ) | ( n2760 & ~n2762 ) | ( n2761 & ~n2762 );
  assign n2764 = ~n2749 & n2763 ;
  assign n2765 = n2732 & n2747 ;
  assign n2766 = n2763 & n2765 ;
  assign n2767 = ( n2750 & n2764 ) | ( n2750 & n2766 ) | ( n2764 & n2766 );
  assign n2768 = n2749 | n2767 ;
  assign n2769 = ( n2688 & n2715 ) | ( n2688 & n2768 ) | ( n2715 & n2768 );
  assign n2770 = n2607 | n2609 ;
  assign n2771 = ~n2610 & n2770 ;
  assign n2772 = n2710 & n2771 ;
  assign n2773 = n2579 & n2703 ;
  assign n2774 = n2587 & n2699 ;
  assign n2775 = n2584 & n2701 ;
  assign n2776 = n2774 | n2775 ;
  assign n2777 = n2773 | n2776 ;
  assign n2778 = n2772 | n2777 ;
  assign n2779 = n949 & n2778 ;
  assign n2780 = n2778 & ~n2779 ;
  assign n2781 = n949 & ~n2779 ;
  assign n2782 = n2780 | n2781 ;
  assign n2783 = ~n2591 & n2669 ;
  assign n2784 = n2587 & n2674 ;
  assign n2785 = ~n2663 & n2673 ;
  assign n2786 = ~n2668 & n2785 ;
  assign n2787 = n2596 & n2786 ;
  assign n2788 = n2784 | n2787 ;
  assign n2789 = n2783 | n2788 ;
  assign n2790 = n2680 & ~n2753 ;
  assign n2791 = n2789 | n2790 ;
  assign n2792 = n453 & n2791 ;
  assign n2793 = n453 | n2791 ;
  assign n2794 = ~n2792 & n2793 ;
  assign n2795 = ~n453 & n587 ;
  assign n2796 = n453 & ~n587 ;
  assign n2797 = n2795 | n2796 ;
  assign n2798 = n2598 & n2797 ;
  assign n2799 = ~n2591 & n2674 ;
  assign n2800 = n2598 & n2786 ;
  assign n2801 = n2596 & n2669 ;
  assign n2802 = n2800 | n2801 ;
  assign n2803 = n2799 | n2802 ;
  assign n2804 = n2680 & ~n2725 ;
  assign n2805 = n2803 | n2804 ;
  assign n2806 = n453 | n2805 ;
  assign n2807 = n453 & n2805 ;
  assign n2808 = n2806 & ~n2807 ;
  assign n2809 = n2686 & n2808 ;
  assign n2810 = ( n2794 & n2798 ) | ( n2794 & n2809 ) | ( n2798 & n2809 );
  assign n2811 = ~n266 & n587 ;
  assign n2812 = n266 & ~n587 ;
  assign n2813 = n2811 | n2812 ;
  assign n2814 = ~n2797 & n2813 ;
  assign n2815 = n2598 & n2814 ;
  assign n2816 = ~n1977 & n2797 ;
  assign n2817 = n2596 & n2816 ;
  assign n2818 = n2815 | n2817 ;
  assign n2819 = n1977 & n2797 ;
  assign n2820 = n2679 & n2819 ;
  assign n2821 = n2818 | n2820 ;
  assign n2822 = n332 & ~n2821 ;
  assign n2823 = n332 & ~n2822 ;
  assign n2824 = ( n2821 & n2822 ) | ( n2821 & ~n2823 ) | ( n2822 & ~n2823 );
  assign n2825 = n332 & n2824 ;
  assign n2826 = ~n2798 & n2825 ;
  assign n2827 = n332 | n2824 ;
  assign n2828 = ( ~n2798 & n2824 ) | ( ~n2798 & n2827 ) | ( n2824 & n2827 );
  assign n2829 = ~n2826 & n2828 ;
  assign n2830 = ~n2591 & n2786 ;
  assign n2831 = n2587 & n2669 ;
  assign n2832 = n2584 & n2674 ;
  assign n2833 = n2831 | n2832 ;
  assign n2834 = n2830 | n2833 ;
  assign n2835 = n2680 & n2709 ;
  assign n2836 = n2834 | n2835 ;
  assign n2837 = n453 | n2836 ;
  assign n2838 = n453 & n2836 ;
  assign n2839 = n2837 & ~n2838 ;
  assign n2840 = ( n2810 & n2829 ) | ( n2810 & n2839 ) | ( n2829 & n2839 );
  assign n2841 = ( n2829 & n2839 ) | ( n2829 & ~n2840 ) | ( n2839 & ~n2840 );
  assign n2842 = ( n2810 & ~n2840 ) | ( n2810 & n2841 ) | ( ~n2840 & n2841 );
  assign n2843 = n2579 & n2699 ;
  assign n2844 = n2575 & n2701 ;
  assign n2845 = n2843 | n2844 ;
  assign n2846 = ~n2572 & n2703 ;
  assign n2847 = n2845 | n2846 ;
  assign n2848 = n2613 & ~n2615 ;
  assign n2849 = ~n2613 & n2615 ;
  assign n2850 = n2848 | n2849 ;
  assign n2851 = n2710 & ~n2850 ;
  assign n2852 = n2847 | n2851 ;
  assign n2853 = n949 & n2852 ;
  assign n2854 = n2852 & ~n2853 ;
  assign n2855 = n949 & ~n2853 ;
  assign n2856 = n2854 | n2855 ;
  assign n2857 = ( n2794 & n2798 ) | ( n2794 & ~n2810 ) | ( n2798 & ~n2810 );
  assign n2858 = ( n2809 & ~n2810 ) | ( n2809 & n2857 ) | ( ~n2810 & n2857 );
  assign n2859 = n2575 & n2703 ;
  assign n2860 = n2584 & n2699 ;
  assign n2861 = n2579 & n2701 ;
  assign n2862 = n2860 | n2861 ;
  assign n2863 = n2859 | n2862 ;
  assign n2864 = n2582 & n2611 ;
  assign n2865 = n2582 | n2611 ;
  assign n2866 = ~n2864 & n2865 ;
  assign n2867 = n2710 & n2866 ;
  assign n2868 = n2863 | n2867 ;
  assign n2869 = n949 | n2868 ;
  assign n2870 = n949 & n2868 ;
  assign n2871 = n2869 & ~n2870 ;
  assign n2872 = n2858 & n2871 ;
  assign n2873 = ( n2842 & n2856 ) | ( n2842 & n2872 ) | ( n2856 & n2872 );
  assign n2874 = n2858 & ~n2871 ;
  assign n2875 = ( n2871 & ~n2872 ) | ( n2871 & n2874 ) | ( ~n2872 & n2874 );
  assign n2876 = n2842 | n2856 ;
  assign n2877 = ( n2873 & n2875 ) | ( n2873 & n2876 ) | ( n2875 & n2876 );
  assign n2878 = ( n2782 & n2873 ) | ( n2782 & n2877 ) | ( n2873 & n2877 );
  assign n2879 = n2686 | n2808 ;
  assign n2880 = ~n2809 & n2879 ;
  assign n2881 = ( n2873 & n2877 ) | ( n2873 & n2880 ) | ( n2877 & n2880 );
  assign n2882 = ( n2769 & n2878 ) | ( n2769 & n2881 ) | ( n2878 & n2881 );
  assign n2883 = n2566 & n2703 ;
  assign n2884 = ~n2572 & n2701 ;
  assign n2885 = n2575 & n2699 ;
  assign n2886 = n2884 | n2885 ;
  assign n2887 = n2883 | n2886 ;
  assign n2888 = n2617 & ~n2622 ;
  assign n2889 = ~n2617 & n2622 ;
  assign n2890 = n2888 | n2889 ;
  assign n2891 = n2710 & ~n2890 ;
  assign n2892 = n2887 | n2891 ;
  assign n2893 = n949 | n2892 ;
  assign n2894 = n949 & n2892 ;
  assign n2895 = n2893 & ~n2894 ;
  assign n2896 = ~n2591 & n2816 ;
  assign n2897 = n1977 & ~n2797 ;
  assign n2898 = ~n2813 & n2897 ;
  assign n2899 = n2598 & n2898 ;
  assign n2900 = n2596 & n2814 ;
  assign n2901 = n2899 | n2900 ;
  assign n2902 = n2896 | n2901 ;
  assign n2903 = ~n2725 & n2819 ;
  assign n2904 = n2902 | n2903 ;
  assign n2905 = n332 | n2904 ;
  assign n2906 = n332 & n2904 ;
  assign n2907 = n2905 & ~n2906 ;
  assign n2908 = n2826 & n2907 ;
  assign n2909 = n2826 | n2907 ;
  assign n2910 = ~n2908 & n2909 ;
  assign n2911 = n2680 & n2771 ;
  assign n2912 = n2579 & n2674 ;
  assign n2913 = n2587 & n2786 ;
  assign n2914 = n2584 & n2669 ;
  assign n2915 = n2913 | n2914 ;
  assign n2916 = n2912 | n2915 ;
  assign n2917 = n2911 | n2916 ;
  assign n2918 = n453 | n2917 ;
  assign n2919 = n453 & n2917 ;
  assign n2920 = n2918 & ~n2919 ;
  assign n2921 = n2910 & n2920 ;
  assign n2922 = n2910 | n2920 ;
  assign n2923 = ~n2921 & n2922 ;
  assign n2924 = n2840 | n2923 ;
  assign n2925 = n2840 & n2923 ;
  assign n2926 = n2924 & ~n2925 ;
  assign n2927 = n2895 & n2926 ;
  assign n2928 = n2895 & ~n2927 ;
  assign n2929 = ~n2895 & n2926 ;
  assign n2930 = n2928 | n2929 ;
  assign n2931 = ~n2591 & n2898 ;
  assign n2932 = n2587 & n2814 ;
  assign n2933 = n2584 & n2816 ;
  assign n2934 = n2932 | n2933 ;
  assign n2935 = n2931 | n2934 ;
  assign n2936 = n2709 & n2819 ;
  assign n2937 = n2935 | n2936 ;
  assign n2938 = n332 & n2937 ;
  assign n2939 = n332 & n2596 ;
  assign n2940 = ~n2938 & n2939 ;
  assign n2941 = n2939 & ~n2940 ;
  assign n2942 = ( n332 & n2937 ) | ( n332 & ~n2940 ) | ( n2937 & ~n2940 );
  assign n2943 = ( ~n2938 & n2941 ) | ( ~n2938 & n2942 ) | ( n2941 & n2942 );
  assign n2944 = ~n2572 & n2674 ;
  assign n2945 = n2579 & n2786 ;
  assign n2946 = n2575 & n2669 ;
  assign n2947 = n2945 | n2946 ;
  assign n2948 = n2944 | n2947 ;
  assign n2949 = n2680 & ~n2850 ;
  assign n2950 = n2948 | n2949 ;
  assign n2951 = n453 & n2950 ;
  assign n2952 = n453 | n2950 ;
  assign n2953 = ~n2951 & n2952 ;
  assign n2954 = ~n2591 & n2814 ;
  assign n2955 = n2587 & n2816 ;
  assign n2956 = n2596 & n2898 ;
  assign n2957 = n2955 | n2956 ;
  assign n2958 = n2954 | n2957 ;
  assign n2959 = ~n2753 & n2819 ;
  assign n2960 = n2958 | n2959 ;
  assign n2961 = n332 & n2960 ;
  assign n2962 = n2960 & ~n2961 ;
  assign n2963 = n332 & ~n2961 ;
  assign n2964 = n2962 | n2963 ;
  assign n2965 = n332 & n2598 ;
  assign n2966 = ( n2908 & n2964 ) | ( n2908 & n2965 ) | ( n2964 & n2965 );
  assign n2967 = ( n2943 & ~n2953 ) | ( n2943 & n2966 ) | ( ~n2953 & n2966 );
  assign n2968 = ( n2953 & ~n2966 ) | ( n2953 & n2967 ) | ( ~n2966 & n2967 );
  assign n2969 = ( ~n2943 & n2967 ) | ( ~n2943 & n2968 ) | ( n2967 & n2968 );
  assign n2970 = ( n2964 & n2965 ) | ( n2964 & ~n2966 ) | ( n2965 & ~n2966 );
  assign n2971 = n2575 & n2674 ;
  assign n2972 = n2584 & n2786 ;
  assign n2973 = n2579 & n2669 ;
  assign n2974 = n2972 | n2973 ;
  assign n2975 = n2971 | n2974 ;
  assign n2976 = n2680 & n2866 ;
  assign n2977 = n2975 | n2976 ;
  assign n2978 = n453 & n2977 ;
  assign n2979 = n453 | n2977 ;
  assign n2980 = ~n2978 & n2979 ;
  assign n2981 = ~n2966 & n2980 ;
  assign n2982 = n2907 & n2980 ;
  assign n2983 = n2826 & n2982 ;
  assign n2984 = ( n2970 & n2981 ) | ( n2970 & n2983 ) | ( n2981 & n2983 );
  assign n2985 = n2966 & ~n2980 ;
  assign n2986 = n2907 | n2980 ;
  assign n2987 = ( n2826 & n2980 ) | ( n2826 & n2986 ) | ( n2980 & n2986 );
  assign n2988 = ( n2970 & ~n2985 ) | ( n2970 & n2987 ) | ( ~n2985 & n2987 );
  assign n2989 = ~n2984 & n2988 ;
  assign n2990 = n2840 | n2921 ;
  assign n2991 = ( n2921 & n2923 ) | ( n2921 & n2990 ) | ( n2923 & n2990 );
  assign n2992 = n2989 & n2991 ;
  assign n2993 = n2984 | n2992 ;
  assign n2994 = ~n2969 & n2993 ;
  assign n2995 = n2969 & ~n2993 ;
  assign n2996 = n2994 | n2995 ;
  assign n2997 = n2558 & n2703 ;
  assign n2998 = n2563 & n2701 ;
  assign n2999 = n2566 & n2699 ;
  assign n3000 = n2998 | n2999 ;
  assign n3001 = n2997 | n3000 ;
  assign n3002 = n2567 | n2569 ;
  assign n3003 = n2626 | n3002 ;
  assign n3004 = ~n2627 & n3003 ;
  assign n3005 = n2710 & n3004 ;
  assign n3006 = n3001 | n3005 ;
  assign n3007 = n949 | n3006 ;
  assign n3008 = n949 & n3006 ;
  assign n3009 = n3007 & ~n3008 ;
  assign n3010 = n2996 & n3009 ;
  assign n3011 = n2996 | n3009 ;
  assign n3012 = ~n3010 & n3011 ;
  assign n3013 = n2989 | n2991 ;
  assign n3014 = ~n2992 & n3013 ;
  assign n3015 = n2563 & n2703 ;
  assign n3016 = n2566 & n2701 ;
  assign n3017 = ~n2572 & n2699 ;
  assign n3018 = n3016 | n3017 ;
  assign n3019 = n3015 | n3018 ;
  assign n3020 = ~n2619 & n2623 ;
  assign n3021 = n2619 | n2620 ;
  assign n3022 = ( n2617 & ~n3020 ) | ( n2617 & n3021 ) | ( ~n3020 & n3021 );
  assign n3023 = ~n2626 & n3022 ;
  assign n3024 = n2710 & n3023 ;
  assign n3025 = n3019 | n3024 ;
  assign n3026 = n949 | n3025 ;
  assign n3027 = n949 & n3025 ;
  assign n3028 = n3026 & ~n3027 ;
  assign n3029 = n3014 | n3028 ;
  assign n3030 = n3012 & n3029 ;
  assign n3031 = n3014 & n3028 ;
  assign n3032 = n3012 & n3031 ;
  assign n3033 = ( ~n2927 & n3014 ) | ( ~n2927 & n3028 ) | ( n3014 & n3028 );
  assign n3034 = n3029 & ~n3033 ;
  assign n3035 = ( n3012 & n3032 ) | ( n3012 & n3034 ) | ( n3032 & n3034 );
  assign n3036 = ( n2930 & n3030 ) | ( n2930 & n3035 ) | ( n3030 & n3035 );
  assign n3037 = n3030 & n3035 ;
  assign n3038 = ( n2882 & n3036 ) | ( n2882 & n3037 ) | ( n3036 & n3037 );
  assign n3039 = n3012 | n3029 ;
  assign n3040 = n3012 | n3031 ;
  assign n3041 = n3034 | n3040 ;
  assign n3042 = ( n2930 & n3039 ) | ( n2930 & n3041 ) | ( n3039 & n3041 );
  assign n3043 = n3039 & n3041 ;
  assign n3044 = ( n2882 & n3042 ) | ( n2882 & n3043 ) | ( n3042 & n3043 );
  assign n3045 = ~n3038 & n3044 ;
  assign n3046 = ~n1222 & n1275 ;
  assign n3047 = n1222 & ~n1275 ;
  assign n3048 = n3046 | n3047 ;
  assign n3049 = n262 & ~n1340 ;
  assign n3050 = ~n262 & n1340 ;
  assign n3051 = n3049 | n3050 ;
  assign n3052 = ~n3048 & n3051 ;
  assign n3053 = n2637 & n3052 ;
  assign n3054 = n1275 & ~n1340 ;
  assign n3055 = ~n1275 & n1340 ;
  assign n3056 = n3054 | n3055 ;
  assign n3057 = n3048 & ~n3051 ;
  assign n3058 = ~n3056 & n3057 ;
  assign n3059 = ~n2555 & n3058 ;
  assign n3060 = ~n3051 & n3056 ;
  assign n3061 = n2552 & n3060 ;
  assign n3062 = n3059 | n3061 ;
  assign n3063 = n3053 | n3062 ;
  assign n3064 = n2634 & n2643 ;
  assign n3065 = n2634 | n2643 ;
  assign n3066 = ~n3064 & n3065 ;
  assign n3067 = n3048 & n3051 ;
  assign n3068 = n3066 & n3067 ;
  assign n3069 = n3063 | n3068 ;
  assign n3070 = n1222 & n3069 ;
  assign n3071 = n1222 | n3069 ;
  assign n3072 = ~n3070 & n3071 ;
  assign n3073 = n3045 & n3072 ;
  assign n3074 = n3045 | n3072 ;
  assign n3075 = ~n3073 & n3074 ;
  assign n3076 = n2927 | n2929 ;
  assign n3077 = n2928 | n3076 ;
  assign n3078 = ( ~n3014 & n3028 ) | ( ~n3014 & n3077 ) | ( n3028 & n3077 );
  assign n3079 = ( n2927 & ~n3014 ) | ( n2927 & n3028 ) | ( ~n3014 & n3028 );
  assign n3080 = ( n2882 & n3078 ) | ( n2882 & n3079 ) | ( n3078 & n3079 );
  assign n3081 = ( n2882 & n2927 ) | ( n2882 & n3077 ) | ( n2927 & n3077 );
  assign n3082 = ( n3028 & ~n3080 ) | ( n3028 & n3081 ) | ( ~n3080 & n3081 );
  assign n3083 = n2552 & n3052 ;
  assign n3084 = n2558 & n3058 ;
  assign n3085 = ~n2555 & n3060 ;
  assign n3086 = n3084 | n3085 ;
  assign n3087 = n3083 | n3086 ;
  assign n3088 = n2630 & ~n2632 ;
  assign n3089 = ~n2630 & n2632 ;
  assign n3090 = n3088 | n3089 ;
  assign n3091 = n3067 & ~n3090 ;
  assign n3092 = n3087 | n3091 ;
  assign n3093 = n1222 & n3092 ;
  assign n3094 = n1222 | n3092 ;
  assign n3095 = ~n3093 & n3094 ;
  assign n3096 = n3080 & n3095 ;
  assign n3097 = n3014 & n3095 ;
  assign n3098 = ( ~n3082 & n3096 ) | ( ~n3082 & n3097 ) | ( n3096 & n3097 );
  assign n3099 = n3080 | n3095 ;
  assign n3100 = n3014 | n3095 ;
  assign n3101 = ( ~n3082 & n3099 ) | ( ~n3082 & n3100 ) | ( n3099 & n3100 );
  assign n3102 = ~n3098 & n3101 ;
  assign n3103 = n2882 & n2930 ;
  assign n3104 = n2882 | n2930 ;
  assign n3105 = ~n3103 & n3104 ;
  assign n3106 = ~n2842 & n2856 ;
  assign n3107 = ( ~n2856 & n2876 ) | ( ~n2856 & n3106 ) | ( n2876 & n3106 );
  assign n3108 = ( n2858 & n2871 ) | ( n2858 & n2880 ) | ( n2871 & n2880 );
  assign n3109 = ~n2769 & n3107 ;
  assign n3110 = ( n2782 & n2858 ) | ( n2782 & n2871 ) | ( n2858 & n2871 );
  assign n3111 = n3107 & ~n3110 ;
  assign n3112 = ( ~n3108 & n3109 ) | ( ~n3108 & n3111 ) | ( n3109 & n3111 );
  assign n3113 = n3107 & ~n3112 ;
  assign n3114 = n2558 & n3052 ;
  assign n3115 = n2566 & n3058 ;
  assign n3116 = n2563 & n3060 ;
  assign n3117 = n3115 | n3116 ;
  assign n3118 = n3114 | n3117 ;
  assign n3119 = n3004 & n3067 ;
  assign n3120 = n3118 | n3119 ;
  assign n3121 = n1222 | n3120 ;
  assign n3122 = n1222 & n3120 ;
  assign n3123 = n3121 & ~n3122 ;
  assign n3124 = n3112 & n3123 ;
  assign n3125 = ( n2769 & n3108 ) | ( n2769 & n3110 ) | ( n3108 & n3110 );
  assign n3126 = n3123 & n3125 ;
  assign n3127 = ( ~n3113 & n3124 ) | ( ~n3113 & n3126 ) | ( n3124 & n3126 );
  assign n3128 = n3112 | n3123 ;
  assign n3129 = n3123 | n3125 ;
  assign n3130 = ( ~n3113 & n3128 ) | ( ~n3113 & n3129 ) | ( n3128 & n3129 );
  assign n3131 = ~n3127 & n3130 ;
  assign n3132 = ( n2769 & n2782 ) | ( n2769 & n2880 ) | ( n2782 & n2880 );
  assign n3133 = n2875 & ~n3132 ;
  assign n3134 = n2875 & n3132 ;
  assign n3135 = ( n3132 & n3133 ) | ( n3132 & ~n3134 ) | ( n3133 & ~n3134 );
  assign n3136 = n2563 & n3052 ;
  assign n3137 = ~n2572 & n3058 ;
  assign n3138 = n2566 & n3060 ;
  assign n3139 = n3137 | n3138 ;
  assign n3140 = n3136 | n3139 ;
  assign n3141 = n3023 & n3067 ;
  assign n3142 = n3140 | n3141 ;
  assign n3143 = n1222 | n3142 ;
  assign n3144 = n1222 & n3142 ;
  assign n3145 = n3143 & ~n3144 ;
  assign n3146 = ~n2890 & n3067 ;
  assign n3147 = ( n2782 & n2880 ) | ( n2782 & ~n3132 ) | ( n2880 & ~n3132 );
  assign n3148 = ( n2769 & ~n3132 ) | ( n2769 & n3147 ) | ( ~n3132 & n3147 );
  assign n3149 = n2566 & n3052 ;
  assign n3150 = ~n2572 & n3060 ;
  assign n3151 = n2575 & ~n3056 ;
  assign n3152 = n3057 & n3151 ;
  assign n3153 = n3150 | n3152 ;
  assign n3154 = n3149 | n3153 ;
  assign n3155 = ( n1222 & n3148 ) | ( n1222 & n3154 ) | ( n3148 & n3154 );
  assign n3156 = n1222 | n3148 ;
  assign n3157 = ( n3146 & n3155 ) | ( n3146 & n3156 ) | ( n3155 & n3156 );
  assign n3158 = n3146 | n3154 ;
  assign n3159 = ( n3148 & ~n3157 ) | ( n3148 & n3158 ) | ( ~n3157 & n3158 );
  assign n3160 = ( n1222 & ~n3157 ) | ( n1222 & n3159 ) | ( ~n3157 & n3159 );
  assign n3161 = ( ~n2688 & n2715 ) | ( ~n2688 & n2768 ) | ( n2715 & n2768 );
  assign n3162 = ( n2688 & ~n2768 ) | ( n2688 & n3161 ) | ( ~n2768 & n3161 );
  assign n3163 = ( ~n2715 & n3161 ) | ( ~n2715 & n3162 ) | ( n3161 & n3162 );
  assign n3164 = ~n2572 & n3052 ;
  assign n3165 = n2575 & n3060 ;
  assign n3166 = n2579 & ~n3056 ;
  assign n3167 = n3057 & n3166 ;
  assign n3168 = n3165 | n3167 ;
  assign n3169 = n3164 | n3168 ;
  assign n3170 = ~n2850 & n3067 ;
  assign n3171 = n3169 | n3170 ;
  assign n3172 = n1222 & n3171 ;
  assign n3173 = n1222 | n3171 ;
  assign n3174 = ~n3172 & n3173 ;
  assign n3175 = n3163 & n3174 ;
  assign n3176 = n3160 & n3175 ;
  assign n3177 = n2579 & n3052 ;
  assign n3178 = n2587 & n3058 ;
  assign n3179 = n2584 & n3060 ;
  assign n3180 = n3178 | n3179 ;
  assign n3181 = n3177 | n3180 ;
  assign n3182 = n2771 & n3067 ;
  assign n3183 = n3181 | n3182 ;
  assign n3184 = n1222 & n3183 ;
  assign n3185 = n1222 | n3183 ;
  assign n3186 = ~n3184 & n3185 ;
  assign n3187 = n2732 | n2747 ;
  assign n3188 = ~n2765 & n3187 ;
  assign n3189 = n3186 & n3188 ;
  assign n3190 = n3186 | n3188 ;
  assign n3191 = ~n3189 & n3190 ;
  assign n3192 = n2740 | n2743 ;
  assign n3193 = ~n2743 & n2745 ;
  assign n3194 = ( n2741 & n3192 ) | ( n2741 & ~n3193 ) | ( n3192 & ~n3193 );
  assign n3195 = ~n2747 & n3194 ;
  assign n3196 = ~n2591 & n3058 ;
  assign n3197 = n2587 & n3060 ;
  assign n3198 = n2584 & n3052 ;
  assign n3199 = n3197 | n3198 ;
  assign n3200 = n3196 | n3199 ;
  assign n3201 = n2709 & n3067 ;
  assign n3202 = n3200 | n3201 ;
  assign n3203 = n1222 | n3202 ;
  assign n3204 = n1222 & n3202 ;
  assign n3205 = n3203 & ~n3204 ;
  assign n3206 = n3195 & n3205 ;
  assign n3207 = n3195 | n3205 ;
  assign n3208 = ~n3206 & n3207 ;
  assign n3209 = n2596 & n3060 ;
  assign n3210 = n2598 & ~n3056 ;
  assign n3211 = n3057 & n3210 ;
  assign n3212 = n3209 | n3211 ;
  assign n3213 = ~n2591 & n3052 ;
  assign n3214 = n3212 | n3213 ;
  assign n3215 = ( ~n2725 & n3067 ) | ( ~n2725 & n3213 ) | ( n3067 & n3213 );
  assign n3216 = n2725 & ~n3067 ;
  assign n3217 = ( n3212 & n3215 ) | ( n3212 & ~n3216 ) | ( n3215 & ~n3216 );
  assign n3218 = n3214 | n3217 ;
  assign n3219 = n1222 | n3218 ;
  assign n3220 = n1222 & n3218 ;
  assign n3221 = n3219 & ~n3220 ;
  assign n3222 = ~n2591 & n3060 ;
  assign n3223 = n2587 & n3052 ;
  assign n3224 = n2596 & n3058 ;
  assign n3225 = n3223 | n3224 ;
  assign n3226 = n3222 | n3225 ;
  assign n3227 = ~n2753 & n3067 ;
  assign n3228 = n3226 | n3227 ;
  assign n3229 = n1222 & n3228 ;
  assign n3230 = n1222 | n3228 ;
  assign n3231 = ~n3229 & n3230 ;
  assign n3232 = n2598 & n3060 ;
  assign n3233 = n2596 & n3052 ;
  assign n3234 = n3232 | n3233 ;
  assign n3235 = n2679 & n3067 ;
  assign n3236 = n1222 & ~n3235 ;
  assign n3237 = ~n3234 & n3236 ;
  assign n3238 = n1222 & ~n3237 ;
  assign n3239 = n1222 & ~n2598 ;
  assign n3240 = ( n1222 & ~n3051 ) | ( n1222 & n3239 ) | ( ~n3051 & n3239 );
  assign n3241 = n3237 & n3240 ;
  assign n3242 = n3234 | n3235 ;
  assign n3243 = n3240 & n3242 ;
  assign n3244 = ( ~n3238 & n3241 ) | ( ~n3238 & n3243 ) | ( n3241 & n3243 );
  assign n3245 = ( n2742 & n3231 ) | ( n2742 & n3244 ) | ( n3231 & n3244 );
  assign n3246 = n2742 & n3231 ;
  assign n3247 = ( n3221 & n3245 ) | ( n3221 & n3246 ) | ( n3245 & n3246 );
  assign n3248 = n3208 & n3247 ;
  assign n3249 = n3189 | n3248 ;
  assign n3250 = n3189 | n3206 ;
  assign n3251 = ( n3191 & n3249 ) | ( n3191 & n3250 ) | ( n3249 & n3250 );
  assign n3252 = n3163 | n3174 ;
  assign n3253 = ~n3175 & n3252 ;
  assign n3254 = n2749 & ~n2763 ;
  assign n3255 = n2763 | n2765 ;
  assign n3256 = ( n2750 & ~n3254 ) | ( n2750 & n3255 ) | ( ~n3254 & n3255 );
  assign n3257 = ~n2767 & n3256 ;
  assign n3258 = n3253 & n3257 ;
  assign n3259 = n2575 & n3052 ;
  assign n3260 = n2584 & n3058 ;
  assign n3261 = n2579 & n3060 ;
  assign n3262 = n3260 | n3261 ;
  assign n3263 = n3259 | n3262 ;
  assign n3264 = ( n2866 & n3067 ) | ( n2866 & n3263 ) | ( n3067 & n3263 );
  assign n3265 = ( n1222 & ~n3067 ) | ( n1222 & n3263 ) | ( ~n3067 & n3263 );
  assign n3266 = ( n1222 & ~n2866 ) | ( n1222 & n3265 ) | ( ~n2866 & n3265 );
  assign n3267 = n3264 | n3266 ;
  assign n3268 = ~n3263 & n3266 ;
  assign n3269 = ( ~n1222 & n3267 ) | ( ~n1222 & n3268 ) | ( n3267 & n3268 );
  assign n3270 = n3253 & n3269 ;
  assign n3271 = ( n3251 & n3258 ) | ( n3251 & n3270 ) | ( n3258 & n3270 );
  assign n3272 = ( n3160 & n3176 ) | ( n3160 & n3271 ) | ( n3176 & n3271 );
  assign n3273 = n1222 & n3158 ;
  assign n3274 = n3157 & ~n3273 ;
  assign n3275 = n3272 | n3274 ;
  assign n3276 = ( n3135 & n3145 ) | ( n3135 & n3275 ) | ( n3145 & n3275 );
  assign n3277 = n3127 | n3276 ;
  assign n3278 = ( n3127 & n3131 ) | ( n3127 & n3277 ) | ( n3131 & n3277 );
  assign n3279 = ~n2555 & n3052 ;
  assign n3280 = n2563 & n3058 ;
  assign n3281 = n2558 & n3060 ;
  assign n3282 = n3280 | n3281 ;
  assign n3283 = n3279 | n3282 ;
  assign n3284 = n2561 & ~n2628 ;
  assign n3285 = ~n2561 & n2628 ;
  assign n3286 = n3284 | n3285 ;
  assign n3287 = n3067 & ~n3286 ;
  assign n3288 = n3283 | n3287 ;
  assign n3289 = n1222 & n3288 ;
  assign n3290 = n1222 | n3288 ;
  assign n3291 = ~n3289 & n3290 ;
  assign n3292 = ( n3105 & n3278 ) | ( n3105 & n3291 ) | ( n3278 & n3291 );
  assign n3293 = n3102 & n3292 ;
  assign n3294 = n3098 | n3293 ;
  assign n3295 = n3075 | n3294 ;
  assign n3296 = ( n3075 & n3098 ) | ( n3075 & n3102 ) | ( n3098 & n3102 );
  assign n3297 = n3075 & n3098 ;
  assign n3298 = ( n3292 & n3296 ) | ( n3292 & n3297 ) | ( n3296 & n3297 );
  assign n3299 = n3295 & ~n3298 ;
  assign n3300 = n2660 & n3299 ;
  assign n3301 = n2660 | n3299 ;
  assign n3302 = ~n3300 & n3301 ;
  assign n3303 = n3102 | n3292 ;
  assign n3304 = ~n3293 & n3303 ;
  assign n3305 = n2533 & n2541 ;
  assign n3306 = n2537 & n2637 ;
  assign n3307 = ~n2536 & n2542 ;
  assign n3308 = n3306 | n3307 ;
  assign n3309 = n3305 | n3308 ;
  assign n3310 = ~n2536 & n2541 ;
  assign n3311 = ( n2536 & ~n2541 ) | ( n2536 & n2638 ) | ( ~n2541 & n2638 );
  assign n3312 = ( n2647 & ~n3310 ) | ( n2647 & n3311 ) | ( ~n3310 & n3311 );
  assign n3313 = n2638 | n2647 ;
  assign n3314 = ( n2536 & ~n3312 ) | ( n2536 & n3313 ) | ( ~n3312 & n3313 );
  assign n3315 = ( n2541 & n3312 ) | ( n2541 & ~n3314 ) | ( n3312 & ~n3314 );
  assign n3316 = n2655 & ~n3315 ;
  assign n3317 = n3309 | n3316 ;
  assign n3318 = n262 | n3317 ;
  assign n3319 = n262 & n3317 ;
  assign n3320 = n3318 & ~n3319 ;
  assign n3321 = n3304 & n3320 ;
  assign n3322 = ~n3304 & n3320 ;
  assign n3323 = ( n3304 & ~n3321 ) | ( n3304 & n3322 ) | ( ~n3321 & n3322 );
  assign n3324 = n2533 & ~n2536 ;
  assign n3325 = n2537 & n2552 ;
  assign n3326 = n2542 & n2637 ;
  assign n3327 = n3325 | n3326 ;
  assign n3328 = n3324 | n3327 ;
  assign n3329 = ( n2634 & n2641 ) | ( n2634 & n2644 ) | ( n2641 & n2644 );
  assign n3330 = n2640 & ~n3329 ;
  assign n3331 = n2647 | n3330 ;
  assign n3332 = n2655 & ~n3331 ;
  assign n3333 = n3328 | n3332 ;
  assign n3334 = n262 | n3333 ;
  assign n3335 = n262 & n3333 ;
  assign n3336 = n3334 & ~n3335 ;
  assign n3337 = ( n3105 & ~n3278 ) | ( n3105 & n3291 ) | ( ~n3278 & n3291 );
  assign n3338 = ( n3278 & ~n3292 ) | ( n3278 & n3337 ) | ( ~n3292 & n3337 );
  assign n3339 = ( ~n3135 & n3145 ) | ( ~n3135 & n3275 ) | ( n3145 & n3275 );
  assign n3340 = ( n3135 & ~n3276 ) | ( n3135 & n3339 ) | ( ~n3276 & n3339 );
  assign n3341 = ~n259 & n2563 ;
  assign n3342 = n2532 & n3341 ;
  assign n3343 = pi0 & ~n3286 ;
  assign n3344 = n2542 & n2558 ;
  assign n3345 = ( n2532 & n3343 ) | ( n2532 & n3344 ) | ( n3343 & n3344 );
  assign n3346 = n2532 | n3343 ;
  assign n3347 = ( n3342 & n3345 ) | ( n3342 & n3346 ) | ( n3345 & n3346 );
  assign n3348 = pi0 & ~n2555 ;
  assign n3349 = ( ~n2532 & n3344 ) | ( ~n2532 & n3348 ) | ( n3344 & n3348 );
  assign n3350 = n2532 & ~n3348 ;
  assign n3351 = ( n3342 & n3349 ) | ( n3342 & ~n3350 ) | ( n3349 & ~n3350 );
  assign n3352 = n3347 | n3351 ;
  assign n3353 = ~n262 & n3352 ;
  assign n3354 = n262 & ~n3352 ;
  assign n3355 = n3353 | n3354 ;
  assign n3356 = n3160 | n3175 ;
  assign n3357 = n3271 | n3356 ;
  assign n3358 = ~n3272 & n3357 ;
  assign n3359 = n3253 | n3257 ;
  assign n3360 = n3253 | n3269 ;
  assign n3361 = ( n3251 & n3359 ) | ( n3251 & n3360 ) | ( n3359 & n3360 );
  assign n3362 = ~n3271 & n3361 ;
  assign n3363 = ( n3355 & n3358 ) | ( n3355 & n3362 ) | ( n3358 & n3362 );
  assign n3364 = pi0 & n2530 ;
  assign n3365 = n3004 & n3364 ;
  assign n3366 = n2542 & n2563 ;
  assign n3367 = pi0 & n2558 ;
  assign n3368 = ( ~n2532 & n3366 ) | ( ~n2532 & n3367 ) | ( n3366 & n3367 );
  assign n3369 = ~n259 & n2566 ;
  assign n3370 = ( n2532 & n3366 ) | ( n2532 & n3369 ) | ( n3366 & n3369 );
  assign n3371 = n3368 | n3370 ;
  assign n3372 = n262 | n3371 ;
  assign n3373 = n2655 | n3372 ;
  assign n3374 = ( n3004 & n3372 ) | ( n3004 & n3373 ) | ( n3372 & n3373 );
  assign n3375 = ~n3365 & n3374 ;
  assign n3376 = n262 & n3371 ;
  assign n3377 = n3375 & ~n3376 ;
  assign n3378 = ( n3355 & n3358 ) | ( n3355 & n3377 ) | ( n3358 & n3377 );
  assign n3379 = n2542 & n2575 ;
  assign n3380 = pi0 & ~n2572 ;
  assign n3381 = ( ~n2532 & n3379 ) | ( ~n2532 & n3380 ) | ( n3379 & n3380 );
  assign n3382 = ~n259 & n2579 ;
  assign n3383 = ( n2532 & n3379 ) | ( n2532 & n3382 ) | ( n3379 & n3382 );
  assign n3384 = n3381 | n3383 ;
  assign n3385 = n2655 | n3384 ;
  assign n3386 = ( ~n2850 & n3384 ) | ( ~n2850 & n3385 ) | ( n3384 & n3385 );
  assign n3387 = n262 | n3386 ;
  assign n3388 = ~n262 & n3386 ;
  assign n3389 = ( ~n3386 & n3387 ) | ( ~n3386 & n3388 ) | ( n3387 & n3388 );
  assign n3390 = n2655 & n2866 ;
  assign n3391 = n2542 & n2579 ;
  assign n3392 = pi0 & n2575 ;
  assign n3393 = ( ~n2532 & n3391 ) | ( ~n2532 & n3392 ) | ( n3391 & n3392 );
  assign n3394 = ~n259 & n2584 ;
  assign n3395 = ( n2532 & n3391 ) | ( n2532 & n3394 ) | ( n3391 & n3394 );
  assign n3396 = n3393 | n3395 ;
  assign n3397 = n3390 | n3396 ;
  assign n3398 = n3221 & n3244 ;
  assign n3399 = n3221 | n3244 ;
  assign n3400 = ~n3398 & n3399 ;
  assign n3401 = n2866 & n3364 ;
  assign n3402 = n3237 | n3240 ;
  assign n3403 = n3240 | n3242 ;
  assign n3404 = ( ~n3238 & n3402 ) | ( ~n3238 & n3403 ) | ( n3402 & n3403 );
  assign n3405 = ~n3244 & n3404 ;
  assign n3406 = n2598 & n3051 ;
  assign n3407 = pi0 & ~n2753 ;
  assign n3408 = n2532 & n3407 ;
  assign n3409 = pi0 & n2587 ;
  assign n3410 = n2542 & ~n2591 ;
  assign n3411 = ( ~n2532 & n3409 ) | ( ~n2532 & n3410 ) | ( n3409 & n3410 );
  assign n3412 = n2532 & ~n3409 ;
  assign n3413 = ( n3408 & n3411 ) | ( n3408 & ~n3412 ) | ( n3411 & ~n3412 );
  assign n3414 = ~n259 & n2596 ;
  assign n3415 = ( n2532 & n3410 ) | ( n2532 & n3414 ) | ( n3410 & n3414 );
  assign n3416 = n2532 | n3414 ;
  assign n3417 = ( n3408 & n3415 ) | ( n3408 & n3416 ) | ( n3415 & n3416 );
  assign n3418 = n3413 | n3417 ;
  assign n3419 = n262 & n3418 ;
  assign n3420 = n262 | n3418 ;
  assign n3421 = ~n3419 & n3420 ;
  assign n3422 = pi0 & n2596 ;
  assign n3423 = ~n2532 & n3422 ;
  assign n3424 = n262 & ~n2598 ;
  assign n3425 = ( n262 & ~n2542 ) | ( n262 & n3424 ) | ( ~n2542 & n3424 );
  assign n3426 = ~n3423 & n3425 ;
  assign n3427 = n2533 & ~n2591 ;
  assign n3428 = n2537 & n2598 ;
  assign n3429 = n2542 & n2596 ;
  assign n3430 = n3428 | n3429 ;
  assign n3431 = n3427 | n3430 ;
  assign n3432 = n262 & n3431 ;
  assign n3433 = pi0 & n2679 ;
  assign n3434 = n2530 & n3433 ;
  assign n3435 = n3432 | n3434 ;
  assign n3436 = n2598 | n2725 ;
  assign n3437 = n2530 & ~n3436 ;
  assign n3438 = ( pi0 & n2598 ) | ( pi0 & n3437 ) | ( n2598 & n3437 );
  assign n3439 = n3435 | n3438 ;
  assign n3440 = n3426 & ~n3439 ;
  assign n3441 = ( n3406 & n3421 ) | ( n3406 & n3440 ) | ( n3421 & n3440 );
  assign n3442 = n259 | n2591 ;
  assign n3443 = n2532 & ~n3442 ;
  assign n3444 = n2542 & n2587 ;
  assign n3445 = pi0 & n2584 ;
  assign n3446 = ~n2532 & n3445 ;
  assign n3447 = n3444 | n3446 ;
  assign n3448 = ( ~n262 & n3443 ) | ( ~n262 & n3447 ) | ( n3443 & n3447 );
  assign n3449 = n262 & ~n3442 ;
  assign n3450 = n2532 & n3449 ;
  assign n3451 = pi0 & n2709 ;
  assign n3452 = n2532 & n3451 ;
  assign n3453 = ( n262 & ~n3450 ) | ( n262 & n3452 ) | ( ~n3450 & n3452 );
  assign n3454 = ~n3447 & n3453 ;
  assign n3455 = ( n3448 & ~n3450 ) | ( n3448 & n3454 ) | ( ~n3450 & n3454 );
  assign n3456 = n2530 & n3451 ;
  assign n3457 = n3455 & ~n3456 ;
  assign n3458 = ( n3405 & n3441 ) | ( n3405 & n3457 ) | ( n3441 & n3457 );
  assign n3459 = ~n3401 & n3458 ;
  assign n3460 = n2533 & n2579 ;
  assign n3461 = n2537 & n2587 ;
  assign n3462 = n2542 & n2584 ;
  assign n3463 = n3461 | n3462 ;
  assign n3464 = n3460 | n3463 ;
  assign n3465 = n2655 & n2771 ;
  assign n3466 = n3464 | n3465 ;
  assign n3467 = n262 & ~n3466 ;
  assign n3468 = ( ~n262 & n3466 ) | ( ~n262 & n3467 ) | ( n3466 & n3467 );
  assign n3469 = n3467 | n3468 ;
  assign n3470 = ~n3401 & n3469 ;
  assign n3471 = ( n3400 & n3459 ) | ( n3400 & n3470 ) | ( n3459 & n3470 );
  assign n3472 = ( n262 & n3397 ) | ( n262 & n3471 ) | ( n3397 & n3471 );
  assign n3473 = ( n262 & n3397 ) | ( n262 & ~n3401 ) | ( n3397 & ~n3401 );
  assign n3474 = ( ~n2742 & n3231 ) | ( ~n2742 & n3244 ) | ( n3231 & n3244 );
  assign n3475 = ~n2742 & n3231 ;
  assign n3476 = ( n3221 & n3474 ) | ( n3221 & n3475 ) | ( n3474 & n3475 );
  assign n3477 = ( n2742 & ~n3398 ) | ( n2742 & n3476 ) | ( ~n3398 & n3476 );
  assign n3478 = ( ~n3231 & n3476 ) | ( ~n3231 & n3477 ) | ( n3476 & n3477 );
  assign n3479 = ( n3472 & n3473 ) | ( n3472 & n3478 ) | ( n3473 & n3478 );
  assign n3480 = ( n262 & n3396 ) | ( n262 & ~n3471 ) | ( n3396 & ~n3471 );
  assign n3481 = ( n262 & n3396 ) | ( n262 & n3401 ) | ( n3396 & n3401 );
  assign n3482 = ( ~n3478 & n3480 ) | ( ~n3478 & n3481 ) | ( n3480 & n3481 );
  assign n3483 = n3479 & ~n3482 ;
  assign n3484 = n3389 & n3458 ;
  assign n3485 = n3389 & n3469 ;
  assign n3486 = ( n3400 & n3484 ) | ( n3400 & n3485 ) | ( n3484 & n3485 );
  assign n3487 = n3478 & n3486 ;
  assign n3488 = ( n3389 & n3483 ) | ( n3389 & n3487 ) | ( n3483 & n3487 );
  assign n3489 = n3208 | n3247 ;
  assign n3490 = ~n3248 & n3489 ;
  assign n3491 = n3389 | n3458 ;
  assign n3492 = n3389 | n3469 ;
  assign n3493 = ( n3400 & n3491 ) | ( n3400 & n3492 ) | ( n3491 & n3492 );
  assign n3494 = ( n3389 & n3478 ) | ( n3389 & n3493 ) | ( n3478 & n3493 );
  assign n3495 = n3490 & n3494 ;
  assign n3496 = ( n3483 & n3490 ) | ( n3483 & n3495 ) | ( n3490 & n3495 );
  assign n3497 = n3488 | n3496 ;
  assign n3498 = ( n3251 & n3257 ) | ( n3251 & n3269 ) | ( n3257 & n3269 );
  assign n3499 = ( n3251 & n3257 ) | ( n3251 & ~n3498 ) | ( n3257 & ~n3498 );
  assign n3500 = n3023 & n3364 ;
  assign n3501 = n2542 & n2566 ;
  assign n3502 = n259 | n2572 ;
  assign n3503 = ( n2532 & n3501 ) | ( n2532 & ~n3502 ) | ( n3501 & ~n3502 );
  assign n3504 = pi0 & n2563 ;
  assign n3505 = ( ~n2532 & n3501 ) | ( ~n2532 & n3504 ) | ( n3501 & n3504 );
  assign n3506 = n3503 | n3505 ;
  assign n3507 = n2655 | n3506 ;
  assign n3508 = ( n3023 & n3506 ) | ( n3023 & n3507 ) | ( n3506 & n3507 );
  assign n3509 = ( n262 & ~n3500 ) | ( n262 & n3508 ) | ( ~n3500 & n3508 );
  assign n3510 = ( n262 & n3364 ) | ( n262 & n3506 ) | ( n3364 & n3506 );
  assign n3511 = n262 & n3506 ;
  assign n3512 = ( n3023 & n3510 ) | ( n3023 & n3511 ) | ( n3510 & n3511 );
  assign n3513 = n3509 & ~n3512 ;
  assign n3514 = ( n3191 & n3206 ) | ( n3191 & n3248 ) | ( n3206 & n3248 );
  assign n3515 = n3206 | n3248 ;
  assign n3516 = n3191 | n3515 ;
  assign n3517 = ~n3514 & n3516 ;
  assign n3518 = ( ~n3498 & n3513 ) | ( ~n3498 & n3517 ) | ( n3513 & n3517 );
  assign n3519 = ( n3269 & n3513 ) | ( n3269 & n3517 ) | ( n3513 & n3517 );
  assign n3520 = ( n3499 & n3518 ) | ( n3499 & n3519 ) | ( n3518 & n3519 );
  assign n3521 = ~n2890 & n3364 ;
  assign n3522 = n2542 & ~n2572 ;
  assign n3523 = pi0 & n2566 ;
  assign n3524 = ( ~n2532 & n3522 ) | ( ~n2532 & n3523 ) | ( n3522 & n3523 );
  assign n3525 = ~n259 & n2575 ;
  assign n3526 = ( n2532 & n3522 ) | ( n2532 & n3525 ) | ( n3522 & n3525 );
  assign n3527 = n3524 | n3526 ;
  assign n3528 = n2655 | n3527 ;
  assign n3529 = ( ~n2890 & n3527 ) | ( ~n2890 & n3528 ) | ( n3527 & n3528 );
  assign n3530 = ( n262 & ~n3521 ) | ( n262 & n3529 ) | ( ~n3521 & n3529 );
  assign n3531 = ( n262 & n3364 ) | ( n262 & n3527 ) | ( n3364 & n3527 );
  assign n3532 = n262 & n3527 ;
  assign n3533 = ( ~n2890 & n3531 ) | ( ~n2890 & n3532 ) | ( n3531 & n3532 );
  assign n3534 = n3530 & ~n3533 ;
  assign n3535 = ( ~n3498 & n3513 ) | ( ~n3498 & n3534 ) | ( n3513 & n3534 );
  assign n3536 = ( n3269 & n3513 ) | ( n3269 & n3534 ) | ( n3513 & n3534 );
  assign n3537 = ( n3499 & n3535 ) | ( n3499 & n3536 ) | ( n3535 & n3536 );
  assign n3538 = ( n3497 & n3520 ) | ( n3497 & n3537 ) | ( n3520 & n3537 );
  assign n3539 = ( n3363 & n3378 ) | ( n3363 & n3538 ) | ( n3378 & n3538 );
  assign n3540 = n2655 & ~n3090 ;
  assign n3541 = n2533 & n2552 ;
  assign n3542 = n2537 & n2558 ;
  assign n3543 = n2542 & ~n2555 ;
  assign n3544 = n3542 | n3543 ;
  assign n3545 = n3541 | n3544 ;
  assign n3546 = n3540 | n3545 ;
  assign n3547 = n262 | n3546 ;
  assign n3548 = n262 & n3546 ;
  assign n3549 = n3547 & ~n3548 ;
  assign n3550 = ( n3340 & n3539 ) | ( n3340 & n3549 ) | ( n3539 & n3549 );
  assign n3551 = n3131 & n3276 ;
  assign n3552 = n3131 | n3276 ;
  assign n3553 = ~n3551 & n3552 ;
  assign n3554 = n2655 & n3066 ;
  assign n3555 = n2533 & n2637 ;
  assign n3556 = n2537 & ~n2555 ;
  assign n3557 = n2542 & n2552 ;
  assign n3558 = n3556 | n3557 ;
  assign n3559 = n3555 | n3558 ;
  assign n3560 = n3554 | n3559 ;
  assign n3561 = n262 & ~n3560 ;
  assign n3562 = ( ~n262 & n3560 ) | ( ~n262 & n3561 ) | ( n3560 & n3561 );
  assign n3563 = n3561 | n3562 ;
  assign n3564 = ( n3550 & n3553 ) | ( n3550 & n3563 ) | ( n3553 & n3563 );
  assign n3565 = ( n3336 & n3338 ) | ( n3336 & n3564 ) | ( n3338 & n3564 );
  assign n3566 = n3323 & n3565 ;
  assign n3567 = n3321 | n3566 ;
  assign n3568 = n3302 & n3567 ;
  assign n3569 = n3302 | n3567 ;
  assign n3570 = ~n3568 & n3569 ;
  assign n3571 = n255 & n3570 ;
  assign n3572 = n255 | n3570 ;
  assign n3573 = ~n3571 & n3572 ;
  assign n3574 = n195 | n370 ;
  assign n3575 = n387 | n3574 ;
  assign n3576 = n218 | n398 ;
  assign n3577 = n418 | n1092 ;
  assign n3578 = n268 | n3577 ;
  assign n3579 = n2004 | n3578 ;
  assign n3580 = n196 | n238 ;
  assign n3581 = n397 | n486 ;
  assign n3582 = n3580 | n3581 ;
  assign n3583 = n3579 | n3582 ;
  assign n3584 = n333 | n382 ;
  assign n3585 = n237 | n3584 ;
  assign n3586 = n714 | n3585 ;
  assign n3587 = n272 | n3586 ;
  assign n3588 = n3583 | n3587 ;
  assign n3589 = n410 | n3588 ;
  assign n3590 = n3576 | n3589 ;
  assign n3591 = n132 | n210 ;
  assign n3592 = n143 | n3591 ;
  assign n3593 = n3590 | n3592 ;
  assign n3594 = n97 | n412 ;
  assign n3595 = n641 | n3594 ;
  assign n3596 = n386 | n3595 ;
  assign n3597 = n144 | n3596 ;
  assign n3598 = n727 | n3597 ;
  assign n3599 = n122 | n3598 ;
  assign n3600 = n129 | n3599 ;
  assign n3601 = n176 | n3600 ;
  assign n3602 = n89 | n3601 ;
  assign n3603 = n352 | n3602 ;
  assign n3604 = n123 | n335 ;
  assign n3605 = n3603 | n3604 ;
  assign n3606 = n140 | n309 ;
  assign n3607 = n113 | n2110 ;
  assign n3608 = n3606 | n3607 ;
  assign n3609 = n307 | n405 ;
  assign n3610 = n1080 | n3609 ;
  assign n3611 = n338 | n3610 ;
  assign n3612 = n3608 | n3611 ;
  assign n3613 = n3605 | n3612 ;
  assign n3614 = n3593 | n3613 ;
  assign n3615 = n3575 | n3614 ;
  assign n3616 = n3323 | n3565 ;
  assign n3617 = ~n3566 & n3616 ;
  assign n3618 = n3336 & n3338 ;
  assign n3619 = n3336 & ~n3338 ;
  assign n3620 = ( n3338 & ~n3618 ) | ( n3338 & n3619 ) | ( ~n3618 & n3619 );
  assign n3621 = ~n3564 & n3620 ;
  assign n3622 = n310 | n2134 ;
  assign n3623 = n128 | n2174 ;
  assign n3624 = n3622 | n3623 ;
  assign n3625 = n371 | n1357 ;
  assign n3626 = n3624 | n3625 ;
  assign n3627 = n137 | n1998 ;
  assign n3628 = n143 | n3627 ;
  assign n3629 = n721 | n3628 ;
  assign n3630 = n357 | n2313 ;
  assign n3631 = n2303 | n3630 ;
  assign n3632 = n560 | n3631 ;
  assign n3633 = n3629 | n3632 ;
  assign n3634 = n3626 | n3633 ;
  assign n3635 = n2257 | n3634 ;
  assign n3636 = n288 | n3635 ;
  assign n3637 = n129 | n3636 ;
  assign n3638 = n267 | n3637 ;
  assign n3639 = n234 | n3638 ;
  assign n3640 = n164 | n3639 ;
  assign n3641 = n233 | n3640 ;
  assign n3642 = n411 | n3641 ;
  assign n3643 = ( ~n3620 & n3621 ) | ( ~n3620 & n3642 ) | ( n3621 & n3642 );
  assign n3644 = ( n3564 & n3621 ) | ( n3564 & n3643 ) | ( n3621 & n3643 );
  assign n3645 = ( n3615 & n3617 ) | ( n3615 & n3644 ) | ( n3617 & n3644 );
  assign n3646 = n3573 & n3645 ;
  assign n3647 = n3573 | n3645 ;
  assign n3648 = ~n3646 & n3647 ;
  assign n3649 = n3571 | n3646 ;
  assign n3650 = n216 | n1044 ;
  assign n3651 = n727 | n3650 ;
  assign n3652 = n1362 | n3651 ;
  assign n3653 = n2182 | n3652 ;
  assign n3654 = n528 | n3653 ;
  assign n3655 = n553 | n3654 ;
  assign n3656 = n155 | n3655 ;
  assign n3657 = n196 | n3656 ;
  assign n3658 = n115 | n3657 ;
  assign n3659 = n664 | n3658 ;
  assign n3660 = n3300 | n3568 ;
  assign n3661 = n305 | n476 ;
  assign n3662 = n216 | n3661 ;
  assign n3663 = n107 | n307 ;
  assign n3664 = n149 | n3663 ;
  assign n3665 = n3662 | n3664 ;
  assign n3666 = n333 | n366 ;
  assign n3667 = n3665 | n3666 ;
  assign n3668 = n677 | n3667 ;
  assign n3669 = n365 | n457 ;
  assign n3670 = n1994 | n3669 ;
  assign n3671 = n1074 | n3670 ;
  assign n3672 = n3668 | n3671 ;
  assign n3673 = n210 | n1345 ;
  assign n3674 = n1071 & ~n2111 ;
  assign n3675 = ~n233 & n3674 ;
  assign n3676 = ~n3673 & n3675 ;
  assign n3677 = ~n3672 & n3676 ;
  assign n3678 = ~n225 & n3677 ;
  assign n3679 = ~n120 & n3678 ;
  assign n3680 = n2525 & n3679 ;
  assign n3681 = n2525 | n3679 ;
  assign n3682 = ~n3680 & n3681 ;
  assign n3683 = ~n2526 & n3682 ;
  assign n3684 = n2526 & ~n3682 ;
  assign n3685 = n3683 | n3684 ;
  assign n3686 = n2547 | n2651 ;
  assign n3687 = n3685 | n3686 ;
  assign n3688 = n2547 | n2652 ;
  assign n3689 = n3685 | n3688 ;
  assign n3690 = ( n2647 & n3687 ) | ( n2647 & n3689 ) | ( n3687 & n3689 );
  assign n3691 = ~n3685 & n3690 ;
  assign n3692 = ( n2647 & n3686 ) | ( n2647 & n3688 ) | ( n3686 & n3688 );
  assign n3693 = ( n3690 & n3691 ) | ( n3690 & ~n3692 ) | ( n3691 & ~n3692 );
  assign n3694 = n2655 & ~n3693 ;
  assign n3695 = n2533 & ~n3682 ;
  assign n3696 = n2537 & n2541 ;
  assign n3697 = n2526 & n2542 ;
  assign n3698 = n3696 | n3697 ;
  assign n3699 = n3695 | n3698 ;
  assign n3700 = n3694 | n3699 ;
  assign n3701 = n262 & ~n3700 ;
  assign n3702 = ~n262 & n3700 ;
  assign n3703 = n3701 | n3702 ;
  assign n3704 = ~n2555 & n2703 ;
  assign n3705 = n2558 & n2701 ;
  assign n3706 = n2563 & n2699 ;
  assign n3707 = n3705 | n3706 ;
  assign n3708 = n3704 | n3707 ;
  assign n3709 = n2710 & ~n3286 ;
  assign n3710 = n3708 | n3709 ;
  assign n3711 = n949 & n3710 ;
  assign n3712 = n3710 & ~n3711 ;
  assign n3713 = n949 & ~n3711 ;
  assign n3714 = n3712 | n3713 ;
  assign n3715 = n2943 | n2966 ;
  assign n3716 = n2969 & n2984 ;
  assign n3717 = ( n2969 & n2992 ) | ( n2969 & n3716 ) | ( n2992 & n3716 );
  assign n3718 = ( ~n2967 & n3715 ) | ( ~n2967 & n3717 ) | ( n3715 & n3717 );
  assign n3719 = n2566 & n2674 ;
  assign n3720 = n2575 & n2786 ;
  assign n3721 = ~n2572 & n2669 ;
  assign n3722 = n3720 | n3721 ;
  assign n3723 = n3719 | n3722 ;
  assign n3724 = n2680 & ~n2890 ;
  assign n3725 = n3723 | n3724 ;
  assign n3726 = n453 | n3725 ;
  assign n3727 = n453 & n3725 ;
  assign n3728 = n3726 & ~n3727 ;
  assign n3729 = n2940 | n2943 ;
  assign n3730 = n332 & n2591 ;
  assign n3731 = n2579 & n2816 ;
  assign n3732 = n2587 & n2898 ;
  assign n3733 = n2584 & n2814 ;
  assign n3734 = n3732 | n3733 ;
  assign n3735 = n3731 | n3734 ;
  assign n3736 = n2771 & n2819 ;
  assign n3737 = n3735 | n3736 ;
  assign n3738 = n3730 & n3737 ;
  assign n3739 = n3730 | n3737 ;
  assign n3740 = ~n3738 & n3739 ;
  assign n3741 = n2966 & n3740 ;
  assign n3742 = n2940 & n3740 ;
  assign n3743 = ( n3729 & n3741 ) | ( n3729 & n3742 ) | ( n3741 & n3742 );
  assign n3744 = n2966 | n3740 ;
  assign n3745 = n2940 | n3740 ;
  assign n3746 = ( n3729 & n3744 ) | ( n3729 & n3745 ) | ( n3744 & n3745 );
  assign n3747 = ~n3743 & n3746 ;
  assign n3748 = ( n3715 & n3728 ) | ( n3715 & n3747 ) | ( n3728 & n3747 );
  assign n3749 = ( ~n2967 & n3728 ) | ( ~n2967 & n3747 ) | ( n3728 & n3747 );
  assign n3750 = ( n3717 & n3748 ) | ( n3717 & n3749 ) | ( n3748 & n3749 );
  assign n3751 = ( n3728 & n3747 ) | ( n3728 & ~n3750 ) | ( n3747 & ~n3750 );
  assign n3752 = ( n3718 & ~n3750 ) | ( n3718 & n3751 ) | ( ~n3750 & n3751 );
  assign n3753 = n3714 & n3752 ;
  assign n3754 = n3714 & ~n3753 ;
  assign n3755 = ~n3714 & n3752 ;
  assign n3756 = n3754 | n3755 ;
  assign n3757 = n3010 | n3032 ;
  assign n3758 = n3010 | n3012 ;
  assign n3759 = ( n3034 & n3757 ) | ( n3034 & n3758 ) | ( n3757 & n3758 );
  assign n3760 = n3756 & n3759 ;
  assign n3761 = ( n3010 & n3029 ) | ( n3010 & n3758 ) | ( n3029 & n3758 );
  assign n3762 = n3755 & n3761 ;
  assign n3763 = ( n3754 & n3761 ) | ( n3754 & n3762 ) | ( n3761 & n3762 );
  assign n3764 = ( n3103 & n3760 ) | ( n3103 & n3763 ) | ( n3760 & n3763 );
  assign n3765 = ( n2930 & n3759 ) | ( n2930 & n3761 ) | ( n3759 & n3761 );
  assign n3766 = n3759 & n3761 ;
  assign n3767 = ( n2882 & n3765 ) | ( n2882 & n3766 ) | ( n3765 & n3766 );
  assign n3768 = n3756 | n3767 ;
  assign n3769 = ~n3764 & n3768 ;
  assign n3770 = n3073 | n3298 ;
  assign n3771 = ~n2536 & n3052 ;
  assign n3772 = n2552 & n3058 ;
  assign n3773 = n2637 & n3060 ;
  assign n3774 = n3772 | n3773 ;
  assign n3775 = n3771 | n3774 ;
  assign n3776 = n3067 & ~n3331 ;
  assign n3777 = n3775 | n3776 ;
  assign n3778 = n1222 | n3777 ;
  assign n3779 = n1222 & n3777 ;
  assign n3780 = n3778 & ~n3779 ;
  assign n3781 = ( ~n3769 & n3770 ) | ( ~n3769 & n3780 ) | ( n3770 & n3780 );
  assign n3782 = ( n3770 & n3780 ) | ( n3770 & ~n3781 ) | ( n3780 & ~n3781 );
  assign n3783 = ( n3769 & n3781 ) | ( n3769 & ~n3782 ) | ( n3781 & ~n3782 );
  assign n3784 = n3703 & n3783 ;
  assign n3785 = n3703 | n3783 ;
  assign n3786 = ~n3784 & n3785 ;
  assign n3787 = n3660 & n3786 ;
  assign n3788 = n3300 | n3786 ;
  assign n3789 = n3568 | n3788 ;
  assign n3790 = ~n3787 & n3789 ;
  assign n3791 = n3659 | n3790 ;
  assign n3792 = n3659 & n3789 ;
  assign n3793 = ~n3787 & n3792 ;
  assign n3794 = n3791 & ~n3793 ;
  assign n3795 = n3649 & n3794 ;
  assign n3796 = n3649 | n3794 ;
  assign n3797 = ~n3795 & n3796 ;
  assign n3798 = n3648 & n3797 ;
  assign n3799 = n3648 | n3797 ;
  assign n3800 = ~n3798 & n3799 ;
  assign n3801 = pi22 & ~pi23 ;
  assign n3802 = ~pi22 & pi23 ;
  assign n3803 = n3801 | n3802 ;
  assign n3804 = n3800 & n3803 ;
  assign n3805 = n3793 | n3795 ;
  assign n3806 = n3784 | n3787 ;
  assign n3807 = n397 | n902 ;
  assign n3808 = n213 | n2303 ;
  assign n3809 = n348 | n3808 ;
  assign n3810 = n2038 | n3809 ;
  assign n3811 = n160 | n3810 ;
  assign n3812 = n102 | n3811 ;
  assign n3813 = n157 | n3812 ;
  assign n3814 = n488 | n832 ;
  assign n3815 = n723 | n3814 ;
  assign n3816 = n1359 & ~n1371 ;
  assign n3817 = ~n3815 & n3816 ;
  assign n3818 = ~n159 & n3817 ;
  assign n3819 = ( n2323 & ~n3813 ) | ( n2323 & n3818 ) | ( ~n3813 & n3818 );
  assign n3820 = ~n2323 & n3819 ;
  assign n3821 = ~n3807 & n3820 ;
  assign n3822 = ~n387 & n3821 ;
  assign n3823 = ~n367 & n3822 ;
  assign n3824 = ~n537 & n3823 ;
  assign n3825 = n3680 | n3824 ;
  assign n3826 = n3680 & n3824 ;
  assign n3827 = n3825 & ~n3826 ;
  assign n3828 = n2533 & ~n3827 ;
  assign n3829 = n2526 & n2537 ;
  assign n3830 = n2542 & ~n3682 ;
  assign n3831 = n3829 | n3830 ;
  assign n3832 = n3828 | n3831 ;
  assign n3833 = n3682 | n3827 ;
  assign n3834 = n3682 & n3827 ;
  assign n3835 = n3833 & ~n3834 ;
  assign n3836 = ~n3684 & n3685 ;
  assign n3837 = ( n2526 & n2547 ) | ( n2526 & ~n3682 ) | ( n2547 & ~n3682 );
  assign n3838 = ( n2652 & ~n3836 ) | ( n2652 & n3837 ) | ( ~n3836 & n3837 );
  assign n3839 = ( n2651 & ~n3836 ) | ( n2651 & n3837 ) | ( ~n3836 & n3837 );
  assign n3840 = ( n2647 & n3838 ) | ( n2647 & n3839 ) | ( n3838 & n3839 );
  assign n3841 = n3835 | n3840 ;
  assign n3842 = n3835 & n3840 ;
  assign n3843 = n3841 & ~n3842 ;
  assign n3844 = n2655 & n3843 ;
  assign n3845 = n3832 | n3844 ;
  assign n3846 = n262 & ~n3845 ;
  assign n3847 = ~n262 & n3845 ;
  assign n3848 = n3846 | n3847 ;
  assign n3849 = n2710 & ~n3090 ;
  assign n3850 = n2552 & n2703 ;
  assign n3851 = n2558 & n2699 ;
  assign n3852 = ~n2555 & n2701 ;
  assign n3853 = n3851 | n3852 ;
  assign n3854 = n3850 | n3853 ;
  assign n3855 = n3849 | n3854 ;
  assign n3856 = n949 & n3855 ;
  assign n3857 = n3855 & ~n3856 ;
  assign n3858 = n949 & ~n3856 ;
  assign n3859 = n3857 | n3858 ;
  assign n3860 = n2563 & n2674 ;
  assign n3861 = ~n2572 & n2786 ;
  assign n3862 = n2566 & n2669 ;
  assign n3863 = n3861 | n3862 ;
  assign n3864 = n3860 | n3863 ;
  assign n3865 = n2680 & n3023 ;
  assign n3866 = n3864 | n3865 ;
  assign n3867 = n453 | n3866 ;
  assign n3868 = n453 & n3866 ;
  assign n3869 = n3867 & ~n3868 ;
  assign n3870 = n2575 & n2816 ;
  assign n3871 = n2584 & n2898 ;
  assign n3872 = n2579 & n2814 ;
  assign n3873 = n3871 | n3872 ;
  assign n3874 = n3870 | n3873 ;
  assign n3875 = n2819 & n2866 ;
  assign n3876 = n3874 | n3875 ;
  assign n3877 = n332 & ~n2587 ;
  assign n3878 = n3876 & n3877 ;
  assign n3879 = n3876 | n3877 ;
  assign n3880 = ~n3878 & n3879 ;
  assign n3881 = n332 & ~n2591 ;
  assign n3882 = ~n3737 & n3881 ;
  assign n3883 = n3740 | n3882 ;
  assign n3884 = ( n2966 & n3882 ) | ( n2966 & n3883 ) | ( n3882 & n3883 );
  assign n3885 = n2940 | n3882 ;
  assign n3886 = ( n3740 & n3882 ) | ( n3740 & n3885 ) | ( n3882 & n3885 );
  assign n3887 = ( n3729 & n3884 ) | ( n3729 & n3886 ) | ( n3884 & n3886 );
  assign n3888 = ~n3880 & n3887 ;
  assign n3889 = ( n2940 & n2966 ) | ( n2940 & n3729 ) | ( n2966 & n3729 );
  assign n3890 = n3869 & n3880 ;
  assign n3891 = ~n3883 & n3890 ;
  assign n3892 = n3869 & ~n3882 ;
  assign n3893 = n3880 & n3892 ;
  assign n3894 = ( ~n3889 & n3891 ) | ( ~n3889 & n3893 ) | ( n3891 & n3893 );
  assign n3895 = ( n3869 & n3888 ) | ( n3869 & n3894 ) | ( n3888 & n3894 );
  assign n3896 = n3880 & ~n3887 ;
  assign n3897 = n3888 | n3896 ;
  assign n3898 = ~n3869 & n3897 ;
  assign n3899 = ( n3869 & ~n3895 ) | ( n3869 & n3898 ) | ( ~n3895 & n3898 );
  assign n3900 = n3750 | n3899 ;
  assign n3901 = ~n3750 & n3900 ;
  assign n3902 = ( ~n3899 & n3900 ) | ( ~n3899 & n3901 ) | ( n3900 & n3901 );
  assign n3903 = n3859 & n3902 ;
  assign n3904 = n3859 & ~n3903 ;
  assign n3905 = ~n3859 & n3902 ;
  assign n3906 = n3904 | n3905 ;
  assign n3907 = n3753 & n3905 ;
  assign n3908 = ( n3753 & n3904 ) | ( n3753 & n3907 ) | ( n3904 & n3907 );
  assign n3909 = ( n3760 & n3906 ) | ( n3760 & n3908 ) | ( n3906 & n3908 );
  assign n3910 = ( n3763 & n3906 ) | ( n3763 & n3908 ) | ( n3906 & n3908 );
  assign n3911 = ( n3103 & n3909 ) | ( n3103 & n3910 ) | ( n3909 & n3910 );
  assign n3912 = n3753 | n3905 ;
  assign n3913 = n3904 | n3912 ;
  assign n3914 = n3760 | n3913 ;
  assign n3915 = n3763 | n3913 ;
  assign n3916 = ( n3103 & n3914 ) | ( n3103 & n3915 ) | ( n3914 & n3915 );
  assign n3917 = ~n3911 & n3916 ;
  assign n3918 = n2541 & n3052 ;
  assign n3919 = n2637 & n3058 ;
  assign n3920 = ~n2536 & n3060 ;
  assign n3921 = n3919 | n3920 ;
  assign n3922 = n3918 | n3921 ;
  assign n3923 = n3067 & ~n3315 ;
  assign n3924 = n3922 | n3923 ;
  assign n3925 = n1222 | n3924 ;
  assign n3926 = n1222 & n3924 ;
  assign n3927 = n3925 & ~n3926 ;
  assign n3928 = ~n3917 & n3927 ;
  assign n3929 = n3917 & n3927 ;
  assign n3930 = n3917 & ~n3929 ;
  assign n3931 = ( n3073 & n3769 ) | ( n3073 & n3780 ) | ( n3769 & n3780 );
  assign n3932 = n3928 & n3931 ;
  assign n3933 = ( n3930 & n3931 ) | ( n3930 & n3932 ) | ( n3931 & n3932 );
  assign n3934 = n3769 | n3780 ;
  assign n3935 = n3928 & n3934 ;
  assign n3936 = ( n3930 & n3934 ) | ( n3930 & n3935 ) | ( n3934 & n3935 );
  assign n3937 = ( n3298 & n3933 ) | ( n3298 & n3936 ) | ( n3933 & n3936 );
  assign n3938 = ( n3298 & n3931 ) | ( n3298 & n3934 ) | ( n3931 & n3934 );
  assign n3939 = ( n3917 & ~n3927 ) | ( n3917 & n3938 ) | ( ~n3927 & n3938 );
  assign n3940 = ( n3928 & ~n3937 ) | ( n3928 & n3939 ) | ( ~n3937 & n3939 );
  assign n3941 = n3848 & n3940 ;
  assign n3942 = n3848 | n3940 ;
  assign n3943 = ~n3941 & n3942 ;
  assign n3944 = n3806 & n3943 ;
  assign n3945 = n3784 | n3943 ;
  assign n3946 = n3787 | n3945 ;
  assign n3947 = ~n3944 & n3946 ;
  assign n3948 = n123 | n279 ;
  assign n3949 = n1346 | n3948 ;
  assign n3950 = n523 | n2221 ;
  assign n3951 = n2149 | n3950 ;
  assign n3952 = n2038 | n3951 ;
  assign n3953 = n3949 | n3952 ;
  assign n3954 = n155 | n3953 ;
  assign n3955 = n242 | n3954 ;
  assign n3956 = n165 | n2449 ;
  assign n3957 = n3955 | n3956 ;
  assign n3958 = n137 | n3957 ;
  assign n3959 = n309 | n3958 ;
  assign n3960 = n102 | n333 ;
  assign n3961 = n186 | n3960 ;
  assign n3962 = n3959 | n3961 ;
  assign n3963 = n3947 | n3962 ;
  assign n3964 = n3946 & n3962 ;
  assign n3965 = ~n3944 & n3964 ;
  assign n3966 = n3963 & ~n3965 ;
  assign n3967 = n3805 & n3966 ;
  assign n3968 = n3805 | n3966 ;
  assign n3969 = ~n3967 & n3968 ;
  assign n3970 = n3798 & n3969 ;
  assign n3971 = n3798 | n3969 ;
  assign n3972 = ~n3970 & n3971 ;
  assign n3973 = n3804 & ~n3972 ;
  assign n3974 = ~n3804 & n3972 ;
  assign n3975 = n3973 | n3974 ;
  assign n3976 = n3800 | n3972 ;
  assign n3977 = n3803 & n3976 ;
  assign n3978 = n3965 | n3967 ;
  assign n3979 = n289 | n711 ;
  assign n3980 = n3626 | n3979 ;
  assign n3981 = n219 | n282 ;
  assign n3982 = n203 | n3981 ;
  assign n3983 = n120 | n141 ;
  assign n3984 = n1999 | n3983 ;
  assign n3985 = n3982 | n3984 ;
  assign n3986 = n562 | n3985 ;
  assign n3987 = n3980 | n3986 ;
  assign n3988 = n307 | n3987 ;
  assign n3989 = n350 | n3988 ;
  assign n3990 = n417 | n3989 ;
  assign n3991 = n410 | n3990 ;
  assign n3992 = n113 | n3991 ;
  assign n3993 = n412 | n3992 ;
  assign n3994 = n537 | n3993 ;
  assign n3995 = n2710 & n3066 ;
  assign n3996 = n2637 & n2703 ;
  assign n3997 = ~n2555 & n2699 ;
  assign n3998 = n2552 & n2701 ;
  assign n3999 = n3997 | n3998 ;
  assign n4000 = n3996 | n3999 ;
  assign n4001 = n3995 | n4000 ;
  assign n4002 = n949 & n4001 ;
  assign n4003 = n4001 & ~n4002 ;
  assign n4004 = n949 & ~n4002 ;
  assign n4005 = n4003 | n4004 ;
  assign n4006 = ~n2572 & n2816 ;
  assign n4007 = n2579 & n2898 ;
  assign n4008 = n2575 & n2814 ;
  assign n4009 = n4007 | n4008 ;
  assign n4010 = n4006 | n4009 ;
  assign n4011 = n2819 & ~n2850 ;
  assign n4012 = n4010 | n4011 ;
  assign n4013 = n332 & ~n2584 ;
  assign n4014 = n4012 & n4013 ;
  assign n4015 = n4012 | n4013 ;
  assign n4016 = ~n4014 & n4015 ;
  assign n4017 = n332 & ~n3876 ;
  assign n4018 = n2587 & n4017 ;
  assign n4019 = n3880 | n4018 ;
  assign n4020 = ( n3883 & n4018 ) | ( n3883 & n4019 ) | ( n4018 & n4019 );
  assign n4021 = n4016 & n4020 ;
  assign n4022 = n3882 | n4018 ;
  assign n4023 = ( n3880 & n4018 ) | ( n3880 & n4022 ) | ( n4018 & n4022 );
  assign n4024 = n4016 & n4023 ;
  assign n4025 = ( n3889 & n4021 ) | ( n3889 & n4024 ) | ( n4021 & n4024 );
  assign n4026 = n4016 & ~n4025 ;
  assign n4027 = n2558 & n2674 ;
  assign n4028 = n2566 & n2786 ;
  assign n4029 = n2563 & n2669 ;
  assign n4030 = n4028 | n4029 ;
  assign n4031 = n4027 | n4030 ;
  assign n4032 = n2680 & n3004 ;
  assign n4033 = n4031 | n4032 ;
  assign n4034 = n453 | n4033 ;
  assign n4035 = n453 & n4033 ;
  assign n4036 = n4034 & ~n4035 ;
  assign n4037 = ~n4025 & n4036 ;
  assign n4038 = n4020 & n4036 ;
  assign n4039 = n4023 & n4036 ;
  assign n4040 = ( n3889 & n4038 ) | ( n3889 & n4039 ) | ( n4038 & n4039 );
  assign n4041 = ( n4026 & n4037 ) | ( n4026 & n4040 ) | ( n4037 & n4040 );
  assign n4042 = n4025 & ~n4036 ;
  assign n4043 = n4020 | n4036 ;
  assign n4044 = n4023 | n4036 ;
  assign n4045 = ( n3889 & n4043 ) | ( n3889 & n4044 ) | ( n4043 & n4044 );
  assign n4046 = ( n4026 & ~n4042 ) | ( n4026 & n4045 ) | ( ~n4042 & n4045 );
  assign n4047 = ~n4041 & n4046 ;
  assign n4048 = n3869 | n3895 ;
  assign n4049 = n3898 | n4048 ;
  assign n4050 = n4047 & n4049 ;
  assign n4051 = n3895 & n4047 ;
  assign n4052 = ( n3750 & n4050 ) | ( n3750 & n4051 ) | ( n4050 & n4051 );
  assign n4053 = ( n3750 & n3895 ) | ( n3750 & n4049 ) | ( n3895 & n4049 );
  assign n4054 = n4047 | n4053 ;
  assign n4055 = ~n4052 & n4054 ;
  assign n4056 = n4005 & n4055 ;
  assign n4057 = n4005 & ~n4056 ;
  assign n4058 = ~n4005 & n4055 ;
  assign n4059 = n4057 | n4058 ;
  assign n4060 = n3903 | n3908 ;
  assign n4061 = n3903 | n3905 ;
  assign n4062 = n3904 | n4061 ;
  assign n4063 = ( n3760 & n4060 ) | ( n3760 & n4062 ) | ( n4060 & n4062 );
  assign n4064 = ( n3763 & n4060 ) | ( n3763 & n4062 ) | ( n4060 & n4062 );
  assign n4065 = ( n3103 & n4063 ) | ( n3103 & n4064 ) | ( n4063 & n4064 );
  assign n4066 = n4059 | n4065 ;
  assign n4067 = n4059 & n4065 ;
  assign n4068 = n4066 & ~n4067 ;
  assign n4069 = n2526 & n3052 ;
  assign n4070 = ~n2536 & n3058 ;
  assign n4071 = n2541 & n3060 ;
  assign n4072 = n4070 | n4071 ;
  assign n4073 = n4069 | n4072 ;
  assign n4074 = n2654 & n3067 ;
  assign n4075 = n4073 | n4074 ;
  assign n4076 = n1222 | n4075 ;
  assign n4077 = n1222 & n4075 ;
  assign n4078 = n4076 & ~n4077 ;
  assign n4079 = ~n4068 & n4078 ;
  assign n4080 = n4068 & ~n4078 ;
  assign n4081 = n4079 | n4080 ;
  assign n4082 = n3929 & ~n4081 ;
  assign n4083 = ( n3933 & ~n4081 ) | ( n3933 & n4082 ) | ( ~n4081 & n4082 );
  assign n4084 = ( n3936 & ~n4081 ) | ( n3936 & n4082 ) | ( ~n4081 & n4082 );
  assign n4085 = ( n3298 & n4083 ) | ( n3298 & n4084 ) | ( n4083 & n4084 );
  assign n4086 = n3929 | n3937 ;
  assign n4087 = n4081 | n4085 ;
  assign n4088 = ( n4085 & ~n4086 ) | ( n4085 & n4087 ) | ( ~n4086 & n4087 );
  assign n4089 = n3941 | n3944 ;
  assign n4090 = n2537 & ~n3682 ;
  assign n4091 = n2542 & ~n3827 ;
  assign n4092 = n4090 | n4091 ;
  assign n4093 = ( n3827 & n3833 ) | ( n3827 & ~n3842 ) | ( n3833 & ~n3842 );
  assign n4094 = n3827 & ~n3842 ;
  assign n4095 = n4093 & ~n4094 ;
  assign n4096 = n2655 & n4095 ;
  assign n4097 = n4092 | n4096 ;
  assign n4098 = n262 & n4097 ;
  assign n4099 = n4097 & ~n4098 ;
  assign n4100 = n262 & ~n4098 ;
  assign n4101 = n4099 | n4100 ;
  assign n4102 = ( ~n4088 & n4089 ) | ( ~n4088 & n4101 ) | ( n4089 & n4101 );
  assign n4103 = ( n4089 & n4101 ) | ( n4089 & ~n4102 ) | ( n4101 & ~n4102 );
  assign n4104 = ( n4088 & n4102 ) | ( n4088 & ~n4103 ) | ( n4102 & ~n4103 );
  assign n4105 = n3994 | n4104 ;
  assign n4106 = n3994 & n4104 ;
  assign n4107 = n4105 & ~n4106 ;
  assign n4108 = n3978 & n4107 ;
  assign n4109 = n3978 | n4107 ;
  assign n4110 = ~n4108 & n4109 ;
  assign n4111 = n3970 & n4110 ;
  assign n4112 = n3970 | n4110 ;
  assign n4113 = ~n4111 & n4112 ;
  assign n4114 = n3977 & ~n4113 ;
  assign n4115 = ~n3977 & n4113 ;
  assign n4116 = n4114 | n4115 ;
  assign n4117 = n3976 | n4113 ;
  assign n4118 = n3803 & n4117 ;
  assign n4119 = n4106 | n4108 ;
  assign n4120 = n2221 | n3597 ;
  assign n4121 = n310 | n4120 ;
  assign n4122 = n884 | n4121 ;
  assign n4123 = n2033 | n4122 ;
  assign n4124 = n1370 | n4123 ;
  assign n4125 = n666 | n4124 ;
  assign n4126 = n459 | n4125 ;
  assign n4127 = n267 | n4126 ;
  assign n4128 = n165 | n4127 ;
  assign n4129 = n355 | n4128 ;
  assign n4130 = n94 | n4129 ;
  assign n4131 = n215 | n4130 ;
  assign n4132 = n201 | n4131 ;
  assign n4133 = n2537 & ~n3827 ;
  assign n4134 = n2655 & ~n4093 ;
  assign n4135 = n4133 | n4134 ;
  assign n4136 = n262 & n4135 ;
  assign n4137 = n4135 & ~n4136 ;
  assign n4138 = n262 & ~n4136 ;
  assign n4139 = n4137 | n4138 ;
  assign n4140 = n4041 | n4052 ;
  assign n4141 = ~n2555 & n2674 ;
  assign n4142 = n2563 & n2786 ;
  assign n4143 = n2558 & n2669 ;
  assign n4144 = n4142 | n4143 ;
  assign n4145 = n4141 | n4144 ;
  assign n4146 = n2680 & ~n3286 ;
  assign n4147 = n4145 | n4146 ;
  assign n4148 = n453 | n4147 ;
  assign n4149 = n453 & n4147 ;
  assign n4150 = n4148 & ~n4149 ;
  assign n4151 = n332 & ~n4012 ;
  assign n4152 = n2584 & n4151 ;
  assign n4153 = n4016 | n4152 ;
  assign n4154 = ( n4020 & n4152 ) | ( n4020 & n4153 ) | ( n4152 & n4153 );
  assign n4155 = ( n4023 & n4152 ) | ( n4023 & n4153 ) | ( n4152 & n4153 );
  assign n4156 = ( n3889 & n4154 ) | ( n3889 & n4155 ) | ( n4154 & n4155 );
  assign n4157 = n332 & ~n2579 ;
  assign n4158 = n2566 & n2816 ;
  assign n4159 = n2575 & n2898 ;
  assign n4160 = ~n2572 & n2814 ;
  assign n4161 = n4159 | n4160 ;
  assign n4162 = n4158 | n4161 ;
  assign n4163 = n2819 & ~n2890 ;
  assign n4164 = n4162 | n4163 ;
  assign n4165 = n4157 & n4164 ;
  assign n4166 = n4157 | n4164 ;
  assign n4167 = ~n4165 & n4166 ;
  assign n4168 = n4153 & n4167 ;
  assign n4169 = n4152 & n4167 ;
  assign n4170 = ( n4020 & n4168 ) | ( n4020 & n4169 ) | ( n4168 & n4169 );
  assign n4171 = ( n4023 & n4168 ) | ( n4023 & n4169 ) | ( n4168 & n4169 );
  assign n4172 = ( n3889 & n4170 ) | ( n3889 & n4171 ) | ( n4170 & n4171 );
  assign n4173 = n4156 & ~n4172 ;
  assign n4174 = n4167 & ~n4169 ;
  assign n4175 = ~n4153 & n4167 ;
  assign n4176 = ( ~n4020 & n4174 ) | ( ~n4020 & n4175 ) | ( n4174 & n4175 );
  assign n4177 = ( ~n4023 & n4174 ) | ( ~n4023 & n4175 ) | ( n4174 & n4175 );
  assign n4178 = ( ~n3889 & n4176 ) | ( ~n3889 & n4177 ) | ( n4176 & n4177 );
  assign n4179 = n4150 & n4178 ;
  assign n4180 = ( n4150 & n4173 ) | ( n4150 & n4179 ) | ( n4173 & n4179 );
  assign n4181 = n4150 | n4178 ;
  assign n4182 = n4173 | n4181 ;
  assign n4183 = ~n4180 & n4182 ;
  assign n4184 = n4140 | n4183 ;
  assign n4185 = n4140 & n4183 ;
  assign n4186 = n4184 & ~n4185 ;
  assign n4187 = n2710 & ~n3331 ;
  assign n4188 = ~n2536 & n2703 ;
  assign n4189 = n2552 & n2699 ;
  assign n4190 = n2637 & n2701 ;
  assign n4191 = n4189 | n4190 ;
  assign n4192 = n4188 | n4191 ;
  assign n4193 = n4187 | n4192 ;
  assign n4194 = n949 & n4193 ;
  assign n4195 = n4193 & ~n4194 ;
  assign n4196 = n949 & ~n4194 ;
  assign n4197 = n4195 | n4196 ;
  assign n4198 = n4186 & ~n4197 ;
  assign n4199 = ~n4186 & n4197 ;
  assign n4200 = n4198 | n4199 ;
  assign n4201 = n4005 | n4200 ;
  assign n4202 = n4055 | n4200 ;
  assign n4203 = ( n4065 & n4201 ) | ( n4065 & n4202 ) | ( n4201 & n4202 );
  assign n4204 = n4005 & n4200 ;
  assign n4205 = n4055 & n4200 ;
  assign n4206 = ( n4065 & n4204 ) | ( n4065 & n4205 ) | ( n4204 & n4205 );
  assign n4207 = n4203 & ~n4206 ;
  assign n4208 = n3067 & ~n3690 ;
  assign n4209 = n3067 & n3692 ;
  assign n4210 = ( ~n3691 & n4208 ) | ( ~n3691 & n4209 ) | ( n4208 & n4209 );
  assign n4211 = n3052 & ~n3682 ;
  assign n4212 = n2541 & n3058 ;
  assign n4213 = n2526 & n3060 ;
  assign n4214 = n4212 | n4213 ;
  assign n4215 = n4211 | n4214 ;
  assign n4216 = n1222 | n4215 ;
  assign n4217 = n4210 | n4216 ;
  assign n4218 = n1222 & n4215 ;
  assign n4219 = ( n1222 & n4210 ) | ( n1222 & n4218 ) | ( n4210 & n4218 );
  assign n4220 = n4217 & ~n4219 ;
  assign n4221 = n4207 & n4220 ;
  assign n4222 = n4207 | n4220 ;
  assign n4223 = ~n4221 & n4222 ;
  assign n4224 = n4139 & n4223 ;
  assign n4225 = n4139 | n4223 ;
  assign n4226 = ~n4224 & n4225 ;
  assign n4227 = ( n3929 & n4068 ) | ( n3929 & n4078 ) | ( n4068 & n4078 );
  assign n4228 = n4068 | n4078 ;
  assign n4229 = ( n3937 & n4227 ) | ( n3937 & n4228 ) | ( n4227 & n4228 );
  assign n4230 = n4226 & n4229 ;
  assign n4231 = n4226 | n4229 ;
  assign n4232 = ~n4230 & n4231 ;
  assign n4233 = ( n4085 & n4089 ) | ( n4085 & n4101 ) | ( n4089 & n4101 );
  assign n4234 = ( ~n3929 & n4089 ) | ( ~n3929 & n4101 ) | ( n4089 & n4101 );
  assign n4235 = n4089 & n4101 ;
  assign n4236 = ( ~n3937 & n4234 ) | ( ~n3937 & n4235 ) | ( n4234 & n4235 );
  assign n4237 = ( n4087 & n4233 ) | ( n4087 & n4236 ) | ( n4233 & n4236 );
  assign n4238 = n4232 | n4237 ;
  assign n4239 = n4232 & n4237 ;
  assign n4240 = n4238 & ~n4239 ;
  assign n4241 = n4132 | n4240 ;
  assign n4242 = n4132 & n4240 ;
  assign n4243 = n4241 & ~n4242 ;
  assign n4244 = n4119 & n4243 ;
  assign n4245 = n4119 | n4243 ;
  assign n4246 = ~n4244 & n4245 ;
  assign n4247 = n4111 & n4246 ;
  assign n4248 = n4111 | n4246 ;
  assign n4249 = ~n4247 & n4248 ;
  assign n4250 = n4118 & ~n4249 ;
  assign n4251 = ~n4118 & n4249 ;
  assign n4252 = n4250 | n4251 ;
  assign n4253 = n4242 | n4244 ;
  assign n4254 = n204 | n399 ;
  assign n4255 = n664 | n2110 ;
  assign n4256 = n2346 | n4255 ;
  assign n4257 = n4254 | n4256 ;
  assign n4258 = n129 | n2341 ;
  assign n4259 = n352 | n4258 ;
  assign n4260 = n123 | n2336 ;
  assign n4261 = n4259 | n4260 ;
  assign n4262 = n349 | n2349 ;
  assign n4263 = n120 | n4262 ;
  assign n4264 = n4261 | n4263 ;
  assign n4265 = n4257 | n4264 ;
  assign n4266 = n507 | n4265 ;
  assign n4267 = n935 | n1345 ;
  assign n4268 = n168 | n4267 ;
  assign n4269 = n654 | n4268 ;
  assign n4270 = n4266 | n4269 ;
  assign n4271 = n182 | n4270 ;
  assign n4272 = n475 | n4271 ;
  assign n4273 = n2563 & n2816 ;
  assign n4274 = ~n2572 & n2898 ;
  assign n4275 = n2566 & n2814 ;
  assign n4276 = n4274 | n4275 ;
  assign n4277 = n4273 | n4276 ;
  assign n4278 = n2819 & n3023 ;
  assign n4279 = n4277 | n4278 ;
  assign n4280 = n332 & ~n4279 ;
  assign n4281 = n332 & ~n4280 ;
  assign n4282 = ( n4279 & n4280 ) | ( n4279 & ~n4281 ) | ( n4280 & ~n4281 );
  assign n4283 = n262 & n332 ;
  assign n4284 = n2575 & n4283 ;
  assign n4285 = n262 & ~n4284 ;
  assign n4286 = n2575 & ~n4284 ;
  assign n4287 = n332 & n4286 ;
  assign n4288 = n4285 | n4287 ;
  assign n4289 = n4282 & n4288 ;
  assign n4290 = n4282 & ~n4289 ;
  assign n4291 = n4288 & ~n4289 ;
  assign n4292 = n4290 | n4291 ;
  assign n4293 = n332 & n2579 ;
  assign n4294 = ( ~n4164 & n4172 ) | ( ~n4164 & n4293 ) | ( n4172 & n4293 );
  assign n4295 = n2552 & n2674 ;
  assign n4296 = n2558 & n2786 ;
  assign n4297 = ~n2555 & n2669 ;
  assign n4298 = n4296 | n4297 ;
  assign n4299 = n4295 | n4298 ;
  assign n4300 = n2680 & ~n3090 ;
  assign n4301 = n4299 | n4300 ;
  assign n4302 = n453 & n4301 ;
  assign n4303 = n453 | n4301 ;
  assign n4304 = ~n4302 & n4303 ;
  assign n4305 = ( n4172 & n4292 ) | ( n4172 & ~n4304 ) | ( n4292 & ~n4304 );
  assign n4306 = ~n4292 & n4304 ;
  assign n4307 = ( n4294 & n4305 ) | ( n4294 & ~n4306 ) | ( n4305 & ~n4306 );
  assign n4308 = n4172 | n4294 ;
  assign n4309 = ( n4304 & n4307 ) | ( n4304 & ~n4308 ) | ( n4307 & ~n4308 );
  assign n4310 = ( ~n4292 & n4307 ) | ( ~n4292 & n4309 ) | ( n4307 & n4309 );
  assign n4311 = n4041 | n4180 ;
  assign n4312 = ( n4180 & n4183 ) | ( n4180 & n4311 ) | ( n4183 & n4311 );
  assign n4313 = ~n4310 & n4312 ;
  assign n4314 = n4180 | n4183 ;
  assign n4315 = ~n4310 & n4314 ;
  assign n4316 = ( n4052 & n4313 ) | ( n4052 & n4315 ) | ( n4313 & n4315 );
  assign n4317 = n4310 | n4316 ;
  assign n4318 = n2541 & n2703 ;
  assign n4319 = n2637 & n2699 ;
  assign n4320 = ~n2536 & n2701 ;
  assign n4321 = n4319 | n4320 ;
  assign n4322 = n4318 | n4321 ;
  assign n4323 = n2710 & ~n3312 ;
  assign n4324 = ~n2541 & n2710 ;
  assign n4325 = ( n3314 & n4323 ) | ( n3314 & n4324 ) | ( n4323 & n4324 );
  assign n4326 = n4322 | n4325 ;
  assign n4327 = n949 & ~n4322 ;
  assign n4328 = ~n4325 & n4327 ;
  assign n4329 = n949 & ~n4327 ;
  assign n4330 = ( n949 & n4325 ) | ( n949 & n4329 ) | ( n4325 & n4329 );
  assign n4331 = ( n4326 & n4328 ) | ( n4326 & ~n4330 ) | ( n4328 & ~n4330 );
  assign n4332 = n4316 & n4331 ;
  assign n4333 = ~n4312 & n4331 ;
  assign n4334 = ~n4314 & n4331 ;
  assign n4335 = ( ~n4052 & n4333 ) | ( ~n4052 & n4334 ) | ( n4333 & n4334 );
  assign n4336 = ( n4317 & n4332 ) | ( n4317 & n4335 ) | ( n4332 & n4335 );
  assign n4337 = n4316 | n4331 ;
  assign n4338 = ( n4052 & n4312 ) | ( n4052 & n4314 ) | ( n4312 & n4314 );
  assign n4339 = ~n4331 & n4338 ;
  assign n4340 = ( n4317 & n4337 ) | ( n4317 & ~n4339 ) | ( n4337 & ~n4339 );
  assign n4341 = ~n4336 & n4340 ;
  assign n4342 = n4186 | n4341 ;
  assign n4343 = ( n4197 & n4341 ) | ( n4197 & n4342 ) | ( n4341 & n4342 );
  assign n4344 = n4205 | n4343 ;
  assign n4345 = n4204 | n4343 ;
  assign n4346 = ( n4065 & n4344 ) | ( n4065 & n4345 ) | ( n4344 & n4345 );
  assign n4347 = n4056 | n4058 ;
  assign n4348 = n4057 | n4347 ;
  assign n4349 = ( n4186 & n4197 ) | ( n4186 & n4348 ) | ( n4197 & n4348 );
  assign n4350 = n4341 & n4349 ;
  assign n4351 = ( n4056 & n4186 ) | ( n4056 & n4197 ) | ( n4186 & n4197 );
  assign n4352 = n4341 & n4351 ;
  assign n4353 = ( n4065 & n4350 ) | ( n4065 & n4352 ) | ( n4350 & n4352 );
  assign n4354 = n4346 & ~n4353 ;
  assign n4355 = n3052 & ~n3827 ;
  assign n4356 = n2526 & n3058 ;
  assign n4357 = n3060 & ~n3682 ;
  assign n4358 = n4356 | n4357 ;
  assign n4359 = n4355 | n4358 ;
  assign n4360 = n3067 & n3843 ;
  assign n4361 = n4359 | n4360 ;
  assign n4362 = n1222 & n4361 ;
  assign n4363 = n1222 | n4361 ;
  assign n4364 = ~n4362 & n4363 ;
  assign n4365 = n4354 & n4364 ;
  assign n4366 = n4354 | n4364 ;
  assign n4367 = ~n4365 & n4366 ;
  assign n4368 = n4139 | n4221 ;
  assign n4369 = ( n4221 & n4223 ) | ( n4221 & n4368 ) | ( n4223 & n4368 );
  assign n4370 = n4367 & n4369 ;
  assign n4371 = n4367 | n4369 ;
  assign n4372 = ~n4370 & n4371 ;
  assign n4373 = n4230 | n4372 ;
  assign n4374 = n4232 | n4373 ;
  assign n4375 = ( n4237 & n4373 ) | ( n4237 & n4374 ) | ( n4373 & n4374 );
  assign n4376 = ( n4230 & n4232 ) | ( n4230 & n4372 ) | ( n4232 & n4372 );
  assign n4377 = n4230 & n4372 ;
  assign n4378 = ( n4237 & n4376 ) | ( n4237 & n4377 ) | ( n4376 & n4377 );
  assign n4379 = n4375 & ~n4378 ;
  assign n4380 = n4272 | n4379 ;
  assign n4381 = n4272 & n4379 ;
  assign n4382 = n4380 & ~n4381 ;
  assign n4383 = n4253 & n4382 ;
  assign n4384 = n4253 | n4382 ;
  assign n4385 = ~n4383 & n4384 ;
  assign n4386 = n4247 | n4385 ;
  assign n4387 = n4247 & n4385 ;
  assign n4388 = n4386 & ~n4387 ;
  assign n4389 = n4117 | n4249 ;
  assign n4390 = n3803 & n4389 ;
  assign n4391 = ~n4388 & n4390 ;
  assign n4392 = n4388 & ~n4390 ;
  assign n4393 = n4391 | n4392 ;
  assign n4394 = n4381 | n4383 ;
  assign n4395 = n370 | n2459 ;
  assign n4396 = n89 | n4395 ;
  assign n4397 = n159 | n3813 ;
  assign n4398 = n179 | n726 ;
  assign n4399 = n267 | n405 ;
  assign n4400 = n383 | n4399 ;
  assign n4401 = n4398 | n4400 ;
  assign n4402 = n2188 | n4401 ;
  assign n4403 = n308 | n4402 ;
  assign n4404 = n4397 | n4403 ;
  assign n4405 = n3949 | n4404 ;
  assign n4406 = n4396 | n4405 ;
  assign n4407 = n2002 | n4406 ;
  assign n4408 = n168 | n4407 ;
  assign n4409 = n272 | n4408 ;
  assign n4410 = n281 | n4409 ;
  assign n4411 = n214 | n4410 ;
  assign n4412 = n4370 | n4378 ;
  assign n4413 = n4353 | n4365 ;
  assign n4414 = n2637 & n2674 ;
  assign n4415 = ~n2555 & n2786 ;
  assign n4416 = n2552 & n2669 ;
  assign n4417 = n4415 | n4416 ;
  assign n4418 = n4414 | n4417 ;
  assign n4419 = n2680 & n3066 ;
  assign n4420 = n4418 | n4419 ;
  assign n4421 = n453 | n4420 ;
  assign n4422 = n453 & n4420 ;
  assign n4423 = n4421 & ~n4422 ;
  assign n4424 = n4284 | n4289 ;
  assign n4425 = ~n2572 & n4283 ;
  assign n4426 = n262 & ~n4425 ;
  assign n4427 = n2572 | n4425 ;
  assign n4428 = n332 & ~n4427 ;
  assign n4429 = n4426 | n4428 ;
  assign n4430 = n4424 & n4429 ;
  assign n4431 = n4424 & ~n4430 ;
  assign n4432 = n4429 & ~n4430 ;
  assign n4433 = n4431 | n4432 ;
  assign n4434 = n2558 & n2816 ;
  assign n4435 = n2566 & n2898 ;
  assign n4436 = n2563 & n2814 ;
  assign n4437 = n4435 | n4436 ;
  assign n4438 = n4434 | n4437 ;
  assign n4439 = n2819 & n3004 ;
  assign n4440 = n4438 | n4439 ;
  assign n4441 = n332 | n4440 ;
  assign n4442 = n332 & n4440 ;
  assign n4443 = n4441 & ~n4442 ;
  assign n4444 = ( ~n4423 & n4433 ) | ( ~n4423 & n4443 ) | ( n4433 & n4443 );
  assign n4445 = ( n4423 & n4433 ) | ( n4423 & n4443 ) | ( n4433 & n4443 );
  assign n4446 = ( n4423 & n4444 ) | ( n4423 & ~n4445 ) | ( n4444 & ~n4445 );
  assign n4447 = ~n4164 & n4293 ;
  assign n4448 = n4172 | n4447 ;
  assign n4449 = ( n4292 & n4304 ) | ( n4292 & n4448 ) | ( n4304 & n4448 );
  assign n4450 = n2526 & n2703 ;
  assign n4451 = ~n2536 & n2699 ;
  assign n4452 = n2541 & n2701 ;
  assign n4453 = n4451 | n4452 ;
  assign n4454 = n4450 | n4453 ;
  assign n4455 = n2654 & n2710 ;
  assign n4456 = n4454 | n4455 ;
  assign n4457 = n949 & ~n4456 ;
  assign n4458 = n949 & ~n4457 ;
  assign n4459 = ( n4456 & n4457 ) | ( n4456 & ~n4458 ) | ( n4457 & ~n4458 );
  assign n4460 = ( n4446 & ~n4449 ) | ( n4446 & n4459 ) | ( ~n4449 & n4459 );
  assign n4461 = ( n4446 & n4449 ) | ( n4446 & ~n4459 ) | ( n4449 & ~n4459 );
  assign n4462 = ( ~n4446 & n4460 ) | ( ~n4446 & n4461 ) | ( n4460 & n4461 );
  assign n4463 = ( n4051 & n4312 ) | ( n4051 & n4314 ) | ( n4312 & n4314 );
  assign n4464 = ( n4050 & n4312 ) | ( n4050 & n4314 ) | ( n4312 & n4314 );
  assign n4465 = ( n3750 & n4463 ) | ( n3750 & n4464 ) | ( n4463 & n4464 );
  assign n4466 = n4310 & n4465 ;
  assign n4467 = n4336 | n4466 ;
  assign n4468 = n3058 & ~n3682 ;
  assign n4469 = n3060 & ~n3827 ;
  assign n4470 = n4468 | n4469 ;
  assign n4471 = n3067 & n4095 ;
  assign n4472 = n4470 | n4471 ;
  assign n4473 = n1222 | n4472 ;
  assign n4474 = n1222 & n4472 ;
  assign n4475 = n4473 & ~n4474 ;
  assign n4476 = ( n4462 & n4467 ) | ( n4462 & n4475 ) | ( n4467 & n4475 );
  assign n4477 = ( ~n4462 & n4467 ) | ( ~n4462 & n4475 ) | ( n4467 & n4475 );
  assign n4478 = ( n4462 & ~n4476 ) | ( n4462 & n4477 ) | ( ~n4476 & n4477 );
  assign n4479 = n4413 & n4478 ;
  assign n4480 = n4413 | n4478 ;
  assign n4481 = ~n4479 & n4480 ;
  assign n4482 = n4412 & n4481 ;
  assign n4483 = n4412 | n4481 ;
  assign n4484 = ~n4482 & n4483 ;
  assign n4485 = n4411 | n4484 ;
  assign n4486 = n4411 & n4484 ;
  assign n4487 = n4485 & ~n4486 ;
  assign n4488 = n4394 & n4487 ;
  assign n4489 = n4381 | n4487 ;
  assign n4490 = n4383 | n4489 ;
  assign n4491 = ~n4488 & n4490 ;
  assign n4492 = n4387 | n4491 ;
  assign n4493 = n4387 & n4491 ;
  assign n4494 = n4492 & ~n4493 ;
  assign n4495 = n4388 | n4389 ;
  assign n4496 = n3803 & n4495 ;
  assign n4497 = ~n4494 & n4496 ;
  assign n4498 = n4494 & ~n4496 ;
  assign n4499 = n4497 | n4498 ;
  assign n4500 = n4486 | n4488 ;
  assign n4501 = n832 | n1021 ;
  assign n4502 = n479 | n4501 ;
  assign n4503 = n2312 | n4502 ;
  assign n4504 = n2221 | n4503 ;
  assign n4505 = n2000 | n4504 ;
  assign n4506 = n2002 | n4505 ;
  assign n4507 = n902 | n4506 ;
  assign n4508 = n413 | n4507 ;
  assign n4509 = n930 | n2342 ;
  assign n4510 = n246 | n4509 ;
  assign n4511 = n2507 | n4510 ;
  assign n4512 = n4508 | n4511 ;
  assign n4513 = n311 | n4512 ;
  assign n4514 = n129 | n4513 ;
  assign n4515 = n162 | n4514 ;
  assign n4516 = n160 | n4515 ;
  assign n4517 = n336 | n4516 ;
  assign n4518 = n115 | n4517 ;
  assign n4519 = n3058 & ~n3827 ;
  assign n4520 = n3067 & ~n4093 ;
  assign n4521 = n4519 | n4520 ;
  assign n4522 = ~n1222 & n4521 ;
  assign n4523 = n1222 & ~n4521 ;
  assign n4524 = n4522 | n4523 ;
  assign n4525 = n4449 & n4524 ;
  assign n4526 = n4459 & n4524 ;
  assign n4527 = ( n4446 & n4525 ) | ( n4446 & n4526 ) | ( n4525 & n4526 );
  assign n4528 = n4449 | n4524 ;
  assign n4529 = n4459 | n4524 ;
  assign n4530 = ( n4446 & n4528 ) | ( n4446 & n4529 ) | ( n4528 & n4529 );
  assign n4531 = ~n4527 & n4530 ;
  assign n4532 = n2703 & ~n3682 ;
  assign n4533 = n2541 & n2699 ;
  assign n4534 = n2526 & n2701 ;
  assign n4535 = n4533 | n4534 ;
  assign n4536 = n4532 | n4535 ;
  assign n4537 = ( n2710 & ~n3693 ) | ( n2710 & n4536 ) | ( ~n3693 & n4536 );
  assign n4538 = ( n949 & n4536 ) | ( n949 & ~n4537 ) | ( n4536 & ~n4537 );
  assign n4539 = n4537 | n4538 ;
  assign n4540 = ~n4536 & n4538 ;
  assign n4541 = ( ~n949 & n4539 ) | ( ~n949 & n4540 ) | ( n4539 & n4540 );
  assign n4542 = ~n2536 & n2674 ;
  assign n4543 = n2552 & n2786 ;
  assign n4544 = n2637 & n2669 ;
  assign n4545 = n4543 | n4544 ;
  assign n4546 = n4542 | n4545 ;
  assign n4547 = n2680 & ~n3331 ;
  assign n4548 = n4546 | n4547 ;
  assign n4549 = n453 | n4548 ;
  assign n4550 = n453 & n4548 ;
  assign n4551 = n4549 & ~n4550 ;
  assign n4552 = n4425 | n4430 ;
  assign n4553 = n2566 & n4283 ;
  assign n4554 = n262 & ~n4553 ;
  assign n4555 = n2566 & ~n4553 ;
  assign n4556 = n332 & n4555 ;
  assign n4557 = n4554 | n4556 ;
  assign n4558 = n4552 & n4557 ;
  assign n4559 = n4552 & ~n4558 ;
  assign n4560 = n4557 & ~n4558 ;
  assign n4561 = n4559 | n4560 ;
  assign n4562 = ~n2555 & n2816 ;
  assign n4563 = n2563 & n2898 ;
  assign n4564 = n2558 & n2814 ;
  assign n4565 = n4563 | n4564 ;
  assign n4566 = n4562 | n4565 ;
  assign n4567 = n2819 & ~n3286 ;
  assign n4568 = n4566 | n4567 ;
  assign n4569 = n332 | n4568 ;
  assign n4570 = n332 & n4568 ;
  assign n4571 = n4569 & ~n4570 ;
  assign n4572 = ( ~n4551 & n4561 ) | ( ~n4551 & n4571 ) | ( n4561 & n4571 );
  assign n4573 = ( n4551 & n4561 ) | ( n4551 & n4571 ) | ( n4561 & n4571 );
  assign n4574 = ( n4551 & n4572 ) | ( n4551 & ~n4573 ) | ( n4572 & ~n4573 );
  assign n4575 = ( n4445 & ~n4541 ) | ( n4445 & n4574 ) | ( ~n4541 & n4574 );
  assign n4576 = ( n4541 & ~n4574 ) | ( n4541 & n4575 ) | ( ~n4574 & n4575 );
  assign n4577 = ( ~n4445 & n4575 ) | ( ~n4445 & n4576 ) | ( n4575 & n4576 );
  assign n4578 = n4531 & n4577 ;
  assign n4579 = n4531 | n4577 ;
  assign n4580 = ~n4578 & n4579 ;
  assign n4581 = n4476 & n4580 ;
  assign n4582 = n4476 | n4580 ;
  assign n4583 = ~n4581 & n4582 ;
  assign n4584 = n4412 | n4413 ;
  assign n4585 = ( n4412 & n4478 ) | ( n4412 & n4584 ) | ( n4478 & n4584 );
  assign n4586 = ( n4479 & n4481 ) | ( n4479 & n4585 ) | ( n4481 & n4585 );
  assign n4587 = n4583 & n4586 ;
  assign n4588 = n4583 | n4586 ;
  assign n4589 = ~n4587 & n4588 ;
  assign n4590 = n4518 | n4589 ;
  assign n4591 = n4518 & n4589 ;
  assign n4592 = n4590 & ~n4591 ;
  assign n4593 = n4500 & n4592 ;
  assign n4594 = n4486 | n4592 ;
  assign n4595 = n4488 | n4594 ;
  assign n4596 = ~n4593 & n4595 ;
  assign n4597 = n4493 & n4596 ;
  assign n4598 = n4493 | n4596 ;
  assign n4599 = ~n4597 & n4598 ;
  assign n4600 = n4494 | n4495 ;
  assign n4601 = n3803 & n4600 ;
  assign n4602 = ~n4599 & n4601 ;
  assign n4603 = n4599 & ~n4601 ;
  assign n4604 = n4602 | n4603 ;
  assign n4605 = n4591 | n4593 ;
  assign n4606 = n122 | n2096 ;
  assign n4607 = n386 | n4606 ;
  assign n4608 = n141 | n212 ;
  assign n4609 = n2026 | n4608 ;
  assign n4610 = n200 | n349 ;
  assign n4611 = n2100 | n4610 ;
  assign n4612 = n4609 | n4611 ;
  assign n4613 = n4607 | n4612 ;
  assign n4614 = n2094 | n3606 ;
  assign n4615 = n414 | n459 ;
  assign n4616 = n132 | n523 ;
  assign n4617 = n4615 | n4616 ;
  assign n4618 = n4614 | n4617 ;
  assign n4619 = n4613 | n4618 ;
  assign n4620 = n676 | n4619 ;
  assign n4621 = n2274 | n4620 ;
  assign n4622 = n4400 | n4621 ;
  assign n4623 = n718 | n4622 ;
  assign n4624 = n4508 | n4623 ;
  assign n4625 = n203 | n4624 ;
  assign n4626 = n182 | n4625 ;
  assign n4627 = n143 | n4626 ;
  assign n4628 = n233 | n4627 ;
  assign n4629 = n1040 | n4628 ;
  assign n4630 = n159 | n4629 ;
  assign n4631 = n333 | n4630 ;
  assign n4632 = n2703 & ~n3827 ;
  assign n4633 = n2526 & n2699 ;
  assign n4634 = n2701 & ~n3682 ;
  assign n4635 = n4633 | n4634 ;
  assign n4636 = n4632 | n4635 ;
  assign n4637 = n2710 & n3843 ;
  assign n4638 = n4636 | n4637 ;
  assign n4639 = n949 | n4638 ;
  assign n4640 = n949 & n4638 ;
  assign n4641 = n4639 & ~n4640 ;
  assign n4642 = n4541 & n4641 ;
  assign n4643 = n4443 & n4641 ;
  assign n4644 = n4433 & n4641 ;
  assign n4645 = ( n4423 & n4643 ) | ( n4423 & n4644 ) | ( n4643 & n4644 );
  assign n4646 = ( n4574 & n4642 ) | ( n4574 & n4645 ) | ( n4642 & n4645 );
  assign n4647 = n4541 | n4641 ;
  assign n4648 = n4443 | n4641 ;
  assign n4649 = n4433 | n4641 ;
  assign n4650 = ( n4423 & n4648 ) | ( n4423 & n4649 ) | ( n4648 & n4649 );
  assign n4651 = ( n4574 & n4647 ) | ( n4574 & n4650 ) | ( n4647 & n4650 );
  assign n4652 = ~n4646 & n4651 ;
  assign n4653 = n332 & n2563 ;
  assign n4654 = n262 | n1222 ;
  assign n4655 = n262 & n1222 ;
  assign n4656 = n4654 & ~n4655 ;
  assign n4657 = n4653 & n4656 ;
  assign n4658 = n4653 | n4656 ;
  assign n4659 = ~n4657 & n4658 ;
  assign n4660 = n4553 | n4558 ;
  assign n4661 = n2552 & n2816 ;
  assign n4662 = n2558 & n2898 ;
  assign n4663 = ~n2555 & n2814 ;
  assign n4664 = n4662 | n4663 ;
  assign n4665 = n4661 | n4664 ;
  assign n4666 = n2819 & ~n3090 ;
  assign n4667 = n4665 | n4666 ;
  assign n4668 = n332 & n4667 ;
  assign n4669 = n4667 & ~n4668 ;
  assign n4670 = n332 & ~n4668 ;
  assign n4671 = n4669 | n4670 ;
  assign n4672 = ( n4659 & n4660 ) | ( n4659 & n4671 ) | ( n4660 & n4671 );
  assign n4673 = ( ~n4659 & n4660 ) | ( ~n4659 & n4671 ) | ( n4660 & n4671 );
  assign n4674 = ( n4659 & ~n4672 ) | ( n4659 & n4673 ) | ( ~n4672 & n4673 );
  assign n4675 = n2541 & n2674 ;
  assign n4676 = n2637 & n2786 ;
  assign n4677 = ~n2536 & n2669 ;
  assign n4678 = n4676 | n4677 ;
  assign n4679 = n4675 | n4678 ;
  assign n4680 = n2680 & ~n3315 ;
  assign n4681 = n4679 | n4680 ;
  assign n4682 = n453 | n4681 ;
  assign n4683 = n453 & n4681 ;
  assign n4684 = n4682 & ~n4683 ;
  assign n4685 = ( n4573 & n4674 ) | ( n4573 & n4684 ) | ( n4674 & n4684 );
  assign n4686 = ( n4674 & n4684 ) | ( n4674 & ~n4685 ) | ( n4684 & ~n4685 );
  assign n4687 = ( n4573 & ~n4685 ) | ( n4573 & n4686 ) | ( ~n4685 & n4686 );
  assign n4688 = n4527 | n4531 ;
  assign n4689 = ( n4527 & n4577 ) | ( n4527 & n4688 ) | ( n4577 & n4688 );
  assign n4690 = ( n4652 & n4687 ) | ( n4652 & n4689 ) | ( n4687 & n4689 );
  assign n4691 = ( n4687 & n4689 ) | ( n4687 & ~n4690 ) | ( n4689 & ~n4690 );
  assign n4692 = ( n4652 & ~n4690 ) | ( n4652 & n4691 ) | ( ~n4690 & n4691 );
  assign n4693 = n4581 | n4587 ;
  assign n4694 = n4692 | n4693 ;
  assign n4695 = ( n4581 & n4587 ) | ( n4581 & n4692 ) | ( n4587 & n4692 );
  assign n4696 = n4694 & ~n4695 ;
  assign n4697 = n4631 & n4696 ;
  assign n4698 = n4631 | n4696 ;
  assign n4699 = ~n4697 & n4698 ;
  assign n4700 = n4605 & n4699 ;
  assign n4701 = n4605 | n4699 ;
  assign n4702 = ~n4700 & n4701 ;
  assign n4703 = n4597 & n4702 ;
  assign n4704 = n4597 | n4702 ;
  assign n4705 = ~n4703 & n4704 ;
  assign n4706 = n4599 | n4600 ;
  assign n4707 = n3803 & n4706 ;
  assign n4708 = ~n4705 & n4707 ;
  assign n4709 = n4705 & ~n4707 ;
  assign n4710 = n4708 | n4709 ;
  assign n4711 = n200 | n282 ;
  assign n4712 = n149 | n4711 ;
  assign n4713 = n414 | n4712 ;
  assign n4714 = n226 | n4713 ;
  assign n4715 = n537 | n4714 ;
  assign n4716 = n366 | n4715 ;
  assign n4717 = n148 | n2042 ;
  assign n4718 = n539 | n4717 ;
  assign n4719 = n209 | n4718 ;
  assign n4720 = n234 | n4719 ;
  assign n4721 = n158 | n4720 ;
  assign n4722 = n221 | n4721 ;
  assign n4723 = n335 | n4722 ;
  assign n4724 = n94 | n4723 ;
  assign n4725 = n204 | n4724 ;
  assign n4726 = n905 | n2223 ;
  assign n4727 = n898 | n4726 ;
  assign n4728 = ( ~n3589 & n4725 ) | ( ~n3589 & n4727 ) | ( n4725 & n4727 );
  assign n4729 = n3589 | n4728 ;
  assign n4730 = n4716 | n4729 ;
  assign n4731 = n2699 & ~n3682 ;
  assign n4732 = n2701 & ~n3827 ;
  assign n4733 = n4731 | n4732 ;
  assign n4734 = ( n2710 & n4095 ) | ( n2710 & n4733 ) | ( n4095 & n4733 );
  assign n4735 = ( n949 & n4733 ) | ( n949 & ~n4734 ) | ( n4733 & ~n4734 );
  assign n4736 = n4734 | n4735 ;
  assign n4737 = ~n4733 & n4735 ;
  assign n4738 = ( ~n949 & n4736 ) | ( ~n949 & n4737 ) | ( n4736 & n4737 );
  assign n4739 = n2637 & n2816 ;
  assign n4740 = ~n2555 & n2898 ;
  assign n4741 = n2552 & n2814 ;
  assign n4742 = n4740 | n4741 ;
  assign n4743 = n4739 | n4742 ;
  assign n4744 = n2819 & n3066 ;
  assign n4745 = n4743 | n4744 ;
  assign n4746 = n332 | n4745 ;
  assign n4747 = n332 & n4745 ;
  assign n4748 = n4746 & ~n4747 ;
  assign n4749 = n332 & n2558 ;
  assign n4750 = ~n4653 & n4654 ;
  assign n4751 = ( n4654 & ~n4656 ) | ( n4654 & n4750 ) | ( ~n4656 & n4750 );
  assign n4752 = ( ~n4748 & n4749 ) | ( ~n4748 & n4751 ) | ( n4749 & n4751 );
  assign n4753 = ( n4749 & n4751 ) | ( n4749 & ~n4752 ) | ( n4751 & ~n4752 );
  assign n4754 = ( n4748 & n4752 ) | ( n4748 & ~n4753 ) | ( n4752 & ~n4753 );
  assign n4755 = n2654 & n2680 ;
  assign n4756 = n2526 & n2674 ;
  assign n4757 = ~n2536 & n2786 ;
  assign n4758 = n2541 & n2669 ;
  assign n4759 = n4757 | n4758 ;
  assign n4760 = n4756 | n4759 ;
  assign n4761 = n4755 | n4760 ;
  assign n4762 = n453 & n4761 ;
  assign n4763 = n453 | n4761 ;
  assign n4764 = ~n4762 & n4763 ;
  assign n4765 = ( n4672 & n4754 ) | ( n4672 & n4764 ) | ( n4754 & n4764 );
  assign n4766 = ( n4672 & ~n4754 ) | ( n4672 & n4764 ) | ( ~n4754 & n4764 );
  assign n4767 = ( n4754 & ~n4765 ) | ( n4754 & n4766 ) | ( ~n4765 & n4766 );
  assign n4768 = ( n4685 & ~n4738 ) | ( n4685 & n4767 ) | ( ~n4738 & n4767 );
  assign n4769 = ( n4738 & ~n4767 ) | ( n4738 & n4768 ) | ( ~n4767 & n4768 );
  assign n4770 = n4646 | n4651 ;
  assign n4771 = ( n4646 & ~n4685 ) | ( n4646 & n4770 ) | ( ~n4685 & n4770 );
  assign n4772 = ( n4573 & n4646 ) | ( n4573 & n4770 ) | ( n4646 & n4770 );
  assign n4773 = ( n4686 & n4771 ) | ( n4686 & n4772 ) | ( n4771 & n4772 );
  assign n4774 = n4768 & n4773 ;
  assign n4775 = ~n4685 & n4773 ;
  assign n4776 = ( n4769 & n4774 ) | ( n4769 & n4775 ) | ( n4774 & n4775 );
  assign n4777 = n4768 | n4773 ;
  assign n4778 = n4685 & ~n4773 ;
  assign n4779 = ( n4769 & n4777 ) | ( n4769 & ~n4778 ) | ( n4777 & ~n4778 );
  assign n4780 = ~n4776 & n4779 ;
  assign n4781 = n4652 & ~n4685 ;
  assign n4782 = n4573 & n4652 ;
  assign n4783 = ( n4686 & n4781 ) | ( n4686 & n4782 ) | ( n4781 & n4782 );
  assign n4784 = ( n4690 & n4695 ) | ( n4690 & ~n4783 ) | ( n4695 & ~n4783 );
  assign n4785 = n4780 | n4784 ;
  assign n4786 = n4690 & n4780 ;
  assign n4787 = n4780 & ~n4783 ;
  assign n4788 = ( n4695 & n4786 ) | ( n4695 & n4787 ) | ( n4786 & n4787 );
  assign n4789 = n4785 & ~n4788 ;
  assign n4790 = n4730 | n4789 ;
  assign n4791 = n4730 & n4789 ;
  assign n4792 = n4790 & ~n4791 ;
  assign n4793 = n4605 | n4697 ;
  assign n4794 = ( n4697 & n4699 ) | ( n4697 & n4793 ) | ( n4699 & n4793 );
  assign n4795 = n4792 & n4794 ;
  assign n4796 = n4792 | n4794 ;
  assign n4797 = ~n4795 & n4796 ;
  assign n4798 = n4703 | n4797 ;
  assign n4799 = n4703 & n4797 ;
  assign n4800 = n4798 & ~n4799 ;
  assign n4801 = n4705 | n4706 ;
  assign n4802 = n3803 & n4801 ;
  assign n4803 = ~n4800 & n4802 ;
  assign n4804 = n4800 & ~n4802 ;
  assign n4805 = n4803 | n4804 ;
  assign n4818 = n4776 | n4788 ;
  assign n4819 = n4672 & ~n4754 ;
  assign n4820 = ( n4754 & n4764 ) | ( n4754 & n4819 ) | ( n4764 & n4819 );
  assign n4821 = n2699 & ~n3827 ;
  assign n4822 = n2710 & ~n4093 ;
  assign n4823 = n4821 | n4822 ;
  assign n4824 = n949 & ~n4823 ;
  assign n4825 = ~n949 & n4823 ;
  assign n4826 = n4824 | n4825 ;
  assign n4827 = n4671 & n4826 ;
  assign n4828 = n4660 & n4826 ;
  assign n4829 = ( n4659 & n4827 ) | ( n4659 & n4828 ) | ( n4827 & n4828 );
  assign n4830 = n4754 & n4829 ;
  assign n4831 = ( n4819 & n4826 ) | ( n4819 & n4830 ) | ( n4826 & n4830 );
  assign n4832 = ~n4671 & n4826 ;
  assign n4833 = ~n4660 & n4826 ;
  assign n4834 = ( ~n4659 & n4832 ) | ( ~n4659 & n4833 ) | ( n4832 & n4833 );
  assign n4835 = ( n4754 & n4826 ) | ( n4754 & n4834 ) | ( n4826 & n4834 );
  assign n4836 = ( n4820 & n4831 ) | ( n4820 & n4835 ) | ( n4831 & n4835 );
  assign n4837 = n4764 | n4826 ;
  assign n4838 = n4671 | n4826 ;
  assign n4839 = n4660 | n4826 ;
  assign n4840 = ( n4659 & n4838 ) | ( n4659 & n4839 ) | ( n4838 & n4839 );
  assign n4841 = ( n4754 & n4837 ) | ( n4754 & n4840 ) | ( n4837 & n4840 );
  assign n4842 = ~n4836 & n4841 ;
  assign n4843 = n332 & ~n2561 ;
  assign n4844 = ~n2536 & n2816 ;
  assign n4845 = n2552 & n2898 ;
  assign n4846 = n2637 & n2814 ;
  assign n4847 = n4845 | n4846 ;
  assign n4848 = n4844 | n4847 ;
  assign n4849 = n2819 & ~n3331 ;
  assign n4850 = n4848 | n4849 ;
  assign n4851 = n332 & n4850 ;
  assign n4852 = n4850 & ~n4851 ;
  assign n4853 = n332 & ~n4851 ;
  assign n4854 = n4852 | n4853 ;
  assign n4855 = n4843 | n4854 ;
  assign n4856 = n4843 & n4854 ;
  assign n4857 = n4855 & ~n4856 ;
  assign n4858 = n2674 & ~n3682 ;
  assign n4859 = n2541 & n2786 ;
  assign n4860 = n2526 & n2669 ;
  assign n4861 = n4859 | n4860 ;
  assign n4862 = n4858 | n4861 ;
  assign n4863 = n2680 & ~n3693 ;
  assign n4864 = n4862 | n4863 ;
  assign n4865 = n453 | n4864 ;
  assign n4866 = n453 & n4864 ;
  assign n4867 = n4865 & ~n4866 ;
  assign n4868 = ( n4752 & n4857 ) | ( n4752 & ~n4867 ) | ( n4857 & ~n4867 );
  assign n4869 = ( ~n4752 & n4857 ) | ( ~n4752 & n4867 ) | ( n4857 & n4867 );
  assign n4870 = ( ~n4857 & n4868 ) | ( ~n4857 & n4869 ) | ( n4868 & n4869 );
  assign n4871 = n4841 & ~n4870 ;
  assign n4872 = ~n4836 & n4871 ;
  assign n4873 = n4841 | n4870 ;
  assign n4874 = ( ~n4836 & n4870 ) | ( ~n4836 & n4873 ) | ( n4870 & n4873 );
  assign n4875 = ( ~n4842 & n4872 ) | ( ~n4842 & n4874 ) | ( n4872 & n4874 );
  assign n4876 = ( n4685 & n4738 ) | ( n4685 & n4767 ) | ( n4738 & n4767 );
  assign n4877 = ( ~n4776 & n4875 ) | ( ~n4776 & n4876 ) | ( n4875 & n4876 );
  assign n4878 = n4875 & n4876 ;
  assign n4879 = ( ~n4788 & n4877 ) | ( ~n4788 & n4878 ) | ( n4877 & n4878 );
  assign n4880 = ( n4875 & n4876 ) | ( n4875 & ~n4878 ) | ( n4876 & ~n4878 );
  assign n4881 = ( n4875 & n4876 ) | ( n4875 & ~n4877 ) | ( n4876 & ~n4877 );
  assign n4882 = ( n4788 & n4880 ) | ( n4788 & n4881 ) | ( n4880 & n4881 );
  assign n4883 = ( n4818 & n4879 ) | ( n4818 & ~n4882 ) | ( n4879 & ~n4882 );
  assign n4806 = n115 | n718 ;
  assign n4807 = n305 | n4806 ;
  assign n4808 = n680 | n4807 ;
  assign n4809 = n194 | n4808 ;
  assign n4810 = n2449 | n4809 ;
  assign n4811 = n2323 | n4810 ;
  assign n4812 = n2507 | n4811 ;
  assign n4813 = n311 | n4812 ;
  assign n4814 = n211 | n4813 ;
  assign n4815 = n221 | n4814 ;
  assign n4816 = n3606 | n4815 ;
  assign n4817 = n368 | n4816 ;
  assign n4884 = n4817 & n4883 ;
  assign n4885 = ( n239 & n4883 ) | ( n239 & n4884 ) | ( n4883 & n4884 );
  assign n4886 = n4817 | n4883 ;
  assign n4887 = n239 | n4886 ;
  assign n4888 = ~n4885 & n4887 ;
  assign n4889 = n4791 | n4792 ;
  assign n4890 = ( n4791 & n4794 ) | ( n4791 & n4889 ) | ( n4794 & n4889 );
  assign n4891 = n4888 & n4890 ;
  assign n4892 = n4888 | n4890 ;
  assign n4893 = ~n4891 & n4892 ;
  assign n4894 = n4799 | n4893 ;
  assign n4895 = n4799 & n4893 ;
  assign n4896 = n4894 & ~n4895 ;
  assign n4897 = n4800 | n4801 ;
  assign n4898 = n3803 & n4897 ;
  assign n4899 = ~n4896 & n4898 ;
  assign n4900 = n4896 & ~n4898 ;
  assign n4901 = n4899 | n4900 ;
  assign n4914 = n332 & ~n2555 ;
  assign n4915 = ~n4749 & n4914 ;
  assign n4916 = n4843 & ~n4915 ;
  assign n4917 = ( n4854 & n4915 ) | ( n4854 & ~n4916 ) | ( n4915 & ~n4916 );
  assign n4918 = n332 & n2552 ;
  assign n4919 = ( ~n949 & n4749 ) | ( ~n949 & n4918 ) | ( n4749 & n4918 );
  assign n4920 = ( n949 & ~n4918 ) | ( n949 & n4919 ) | ( ~n4918 & n4919 );
  assign n4921 = ( ~n4749 & n4919 ) | ( ~n4749 & n4920 ) | ( n4919 & n4920 );
  assign n4922 = n4917 & ~n4921 ;
  assign n4923 = ~n4917 & n4921 ;
  assign n4924 = n4922 | n4923 ;
  assign n4925 = n2541 & n2816 ;
  assign n4926 = n2637 & n2898 ;
  assign n4927 = ~n2536 & n2814 ;
  assign n4928 = n4926 | n4927 ;
  assign n4929 = n4925 | n4928 ;
  assign n4930 = n2819 & ~n3315 ;
  assign n4931 = n4929 | n4930 ;
  assign n4932 = n332 & n4931 ;
  assign n4933 = n332 & ~n4932 ;
  assign n4934 = n4931 & ~n4932 ;
  assign n4935 = n4933 | n4934 ;
  assign n4936 = ~n4924 & n4935 ;
  assign n4937 = n4924 & n4935 ;
  assign n4938 = ( n4924 & n4936 ) | ( n4924 & ~n4937 ) | ( n4936 & ~n4937 );
  assign n4939 = n2674 & ~n3827 ;
  assign n4940 = n2526 & n2786 ;
  assign n4941 = n2669 & ~n3682 ;
  assign n4942 = n4940 | n4941 ;
  assign n4943 = n4939 | n4942 ;
  assign n4944 = n2680 & n3843 ;
  assign n4945 = n4943 | n4944 ;
  assign n4946 = n453 | n4945 ;
  assign n4947 = n453 & n4945 ;
  assign n4948 = n4946 & ~n4947 ;
  assign n4949 = n4867 & n4948 ;
  assign n4950 = n4748 & n4948 ;
  assign n4951 = ~n4749 & n4948 ;
  assign n4952 = ( ~n4751 & n4950 ) | ( ~n4751 & n4951 ) | ( n4950 & n4951 );
  assign n4953 = ( ~n4857 & n4949 ) | ( ~n4857 & n4952 ) | ( n4949 & n4952 );
  assign n4954 = n4868 | n4953 ;
  assign n4955 = ~n4867 & n4948 ;
  assign n4956 = ~n4748 & n4948 ;
  assign n4957 = n4749 & n4948 ;
  assign n4958 = ( n4751 & n4956 ) | ( n4751 & n4957 ) | ( n4956 & n4957 );
  assign n4959 = ( n4857 & n4955 ) | ( n4857 & n4958 ) | ( n4955 & n4958 );
  assign n4960 = n4954 & ~n4959 ;
  assign n4961 = n4938 & n4960 ;
  assign n4962 = n4938 | n4960 ;
  assign n4963 = ~n4961 & n4962 ;
  assign n4964 = n4836 | n4963 ;
  assign n4965 = n4841 & n4870 ;
  assign n4966 = ~n4836 & n4965 ;
  assign n4967 = n4964 | n4966 ;
  assign n4968 = ( n4836 & n4963 ) | ( n4836 & n4966 ) | ( n4963 & n4966 );
  assign n4969 = n4967 & ~n4968 ;
  assign n4970 = n4875 | n4876 ;
  assign n4971 = ( n4776 & n4875 ) | ( n4776 & n4876 ) | ( n4875 & n4876 );
  assign n4972 = ( n4788 & n4970 ) | ( n4788 & n4971 ) | ( n4970 & n4971 );
  assign n4973 = n4969 | n4972 ;
  assign n4974 = n4969 & n4971 ;
  assign n4975 = n4969 & n4970 ;
  assign n4976 = ( n4788 & n4974 ) | ( n4788 & n4975 ) | ( n4974 & n4975 );
  assign n4977 = n4973 & ~n4976 ;
  assign n4902 = n202 | n516 ;
  assign n4903 = n374 | n418 ;
  assign n4904 = n4902 | n4903 ;
  assign n4905 = n3602 | n3609 ;
  assign n4906 = n142 | n4905 ;
  assign n4907 = n155 | n4906 ;
  assign n4908 = n1051 | n4907 ;
  assign n4909 = n2507 | n4908 ;
  assign n4910 = n4904 | n4909 ;
  assign n4911 = n298 | n903 ;
  assign n4912 = n187 | n4911 ;
  assign n4913 = n4910 | n4912 ;
  assign n4978 = n4913 & n4977 ;
  assign n4979 = ( n402 & n4977 ) | ( n402 & n4978 ) | ( n4977 & n4978 );
  assign n4980 = n4913 | n4977 ;
  assign n4981 = n402 | n4980 ;
  assign n4982 = ~n4979 & n4981 ;
  assign n4983 = n4884 | n4890 ;
  assign n4984 = n4883 | n4890 ;
  assign n4985 = ( n239 & n4983 ) | ( n239 & n4984 ) | ( n4983 & n4984 );
  assign n4986 = ( n4885 & n4888 ) | ( n4885 & n4985 ) | ( n4888 & n4985 );
  assign n4987 = n4982 & n4986 ;
  assign n4988 = n4982 | n4986 ;
  assign n4989 = ~n4987 & n4988 ;
  assign n4990 = n4895 | n4989 ;
  assign n4991 = n4895 & n4989 ;
  assign n4992 = n4990 & ~n4991 ;
  assign n4993 = n4896 | n4897 ;
  assign n4994 = n3803 & n4993 ;
  assign n4995 = ~n4992 & n4994 ;
  assign n4996 = n4992 & ~n4994 ;
  assign n4997 = n4995 | n4996 ;
  assign n4998 = n276 | n343 ;
  assign n4999 = n404 | n929 ;
  assign n5000 = n838 | n4999 ;
  assign n5001 = n3666 | n5000 ;
  assign n5002 = ( ~n569 & n3665 ) | ( ~n569 & n5001 ) | ( n3665 & n5001 );
  assign n5003 = n3665 & n5001 ;
  assign n5004 = ( ~n565 & n5002 ) | ( ~n565 & n5003 ) | ( n5002 & n5003 );
  assign n5005 = n570 | n5004 ;
  assign n5006 = n4998 | n5005 ;
  assign n5007 = n2526 & n2816 ;
  assign n5008 = ~n2536 & n2898 ;
  assign n5009 = n2541 & n2814 ;
  assign n5010 = n5008 | n5009 ;
  assign n5011 = n5007 | n5010 ;
  assign n5012 = n2654 & n2819 ;
  assign n5013 = n5011 | n5012 ;
  assign n5014 = n332 | n5013 ;
  assign n5015 = n332 & n5013 ;
  assign n5016 = n5014 & ~n5015 ;
  assign n5017 = n332 & n2637 ;
  assign n5018 = ( ~n4919 & n5016 ) | ( ~n4919 & n5017 ) | ( n5016 & n5017 );
  assign n5019 = ( n4919 & ~n5017 ) | ( n4919 & n5018 ) | ( ~n5017 & n5018 );
  assign n5020 = ( ~n5016 & n5018 ) | ( ~n5016 & n5019 ) | ( n5018 & n5019 );
  assign n5021 = n4922 | n4935 ;
  assign n5022 = ( n4922 & ~n4924 ) | ( n4922 & n5021 ) | ( ~n4924 & n5021 );
  assign n5023 = ~n5020 & n5022 ;
  assign n5024 = n2786 & ~n3682 ;
  assign n5025 = n2669 & ~n3827 ;
  assign n5026 = n5024 | n5025 ;
  assign n5027 = n2680 & n4095 ;
  assign n5028 = n5026 | n5027 ;
  assign n5029 = n453 & n5028 ;
  assign n5030 = n453 | n5028 ;
  assign n5031 = ~n5029 & n5030 ;
  assign n5032 = ( ~n5020 & n5022 ) | ( ~n5020 & n5031 ) | ( n5022 & n5031 );
  assign n5033 = ~n5023 & n5032 ;
  assign n5034 = n5018 & ~n5031 ;
  assign n5035 = n5016 | n5031 ;
  assign n5036 = ( n5019 & n5034 ) | ( n5019 & ~n5035 ) | ( n5034 & ~n5035 );
  assign n5037 = ( n5022 & ~n5031 ) | ( n5022 & n5036 ) | ( ~n5031 & n5036 );
  assign n5038 = ( ~n5022 & n5023 ) | ( ~n5022 & n5037 ) | ( n5023 & n5037 );
  assign n5039 = n5033 | n5038 ;
  assign n5040 = ~n4953 & n4962 ;
  assign n5041 = n4968 | n4971 ;
  assign n5042 = ( n4968 & n4969 ) | ( n4968 & n5041 ) | ( n4969 & n5041 );
  assign n5043 = ( n5039 & n5040 ) | ( n5039 & ~n5042 ) | ( n5040 & ~n5042 );
  assign n5044 = n4968 | n4970 ;
  assign n5045 = ( n4968 & n4969 ) | ( n4968 & n5044 ) | ( n4969 & n5044 );
  assign n5046 = ( n5039 & n5040 ) | ( n5039 & ~n5045 ) | ( n5040 & ~n5045 );
  assign n5047 = ( ~n4788 & n5043 ) | ( ~n4788 & n5046 ) | ( n5043 & n5046 );
  assign n5048 = ( n4788 & n5042 ) | ( n4788 & n5045 ) | ( n5042 & n5045 );
  assign n5049 = ( ~n5040 & n5047 ) | ( ~n5040 & n5048 ) | ( n5047 & n5048 );
  assign n5050 = ( ~n5039 & n5047 ) | ( ~n5039 & n5049 ) | ( n5047 & n5049 );
  assign n5051 = n5006 | n5050 ;
  assign n5052 = n5006 & n5050 ;
  assign n5053 = n5051 & ~n5052 ;
  assign n5054 = n4979 | n4982 ;
  assign n5055 = ( n4979 & n4986 ) | ( n4979 & n5054 ) | ( n4986 & n5054 );
  assign n5056 = n5053 & n5055 ;
  assign n5057 = n5053 | n5055 ;
  assign n5058 = ~n5056 & n5057 ;
  assign n5059 = n4991 | n5058 ;
  assign n5060 = n4991 & n5058 ;
  assign n5061 = n5059 & ~n5060 ;
  assign n5062 = n4992 | n4993 ;
  assign n5063 = n3803 & n5062 ;
  assign n5064 = ~n5061 & n5063 ;
  assign n5065 = n5061 & ~n5063 ;
  assign n5066 = n5064 | n5065 ;
  assign n5067 = n2122 | n3985 ;
  assign n5068 = n167 | n398 ;
  assign n5069 = n176 | n5068 ;
  assign n5070 = n149 | n5069 ;
  assign n5071 = n211 | n5070 ;
  assign n5072 = n2243 | n5071 ;
  assign n5073 = n884 | n5072 ;
  assign n5074 = n5067 | n5073 ;
  assign n5075 = n122 | n5074 ;
  assign n5076 = n112 | n5075 ;
  assign n5077 = n204 | n5076 ;
  assign n5078 = n2011 | n5077 ;
  assign n5079 = n332 & ~n2536 ;
  assign n5080 = ~n5017 & n5079 ;
  assign n5081 = n5017 & ~n5079 ;
  assign n5082 = n5080 | n5081 ;
  assign n5083 = ( n4919 & n5016 ) | ( n4919 & ~n5017 ) | ( n5016 & ~n5017 );
  assign n5084 = n5082 | n5083 ;
  assign n5085 = n5082 & n5083 ;
  assign n5086 = n5084 & ~n5085 ;
  assign n5087 = n2786 & ~n3827 ;
  assign n5088 = n2680 & ~n4093 ;
  assign n5089 = n5087 | n5088 ;
  assign n5090 = n453 | n5089 ;
  assign n5091 = n453 & n5089 ;
  assign n5092 = n5090 & ~n5091 ;
  assign n5093 = n2816 & ~n3682 ;
  assign n5094 = n2541 & n2898 ;
  assign n5095 = n2526 & n2814 ;
  assign n5096 = n5094 | n5095 ;
  assign n5097 = n5093 | n5096 ;
  assign n5098 = n2819 & ~n3693 ;
  assign n5099 = n5097 | n5098 ;
  assign n5100 = n332 & n5099 ;
  assign n5101 = n332 & ~n5100 ;
  assign n5102 = n5099 & ~n5100 ;
  assign n5103 = n5101 | n5102 ;
  assign n5104 = n5092 & n5103 ;
  assign n5105 = n5103 & ~n5104 ;
  assign n5106 = ( n5092 & ~n5104 ) | ( n5092 & n5105 ) | ( ~n5104 & n5105 );
  assign n5107 = n5086 & ~n5106 ;
  assign n5108 = n5106 | n5107 ;
  assign n5109 = ( ~n5086 & n5107 ) | ( ~n5086 & n5108 ) | ( n5107 & n5108 );
  assign n5110 = ~n5023 & n5109 ;
  assign n5111 = ~n5033 & n5110 ;
  assign n5112 = n5032 & ~n5109 ;
  assign n5113 = n5111 | n5112 ;
  assign n5114 = n5047 & n5113 ;
  assign n5115 = n5039 | n5040 ;
  assign n5116 = n5039 & n5040 ;
  assign n5117 = n5115 & ~n5116 ;
  assign n5118 = n4968 & n5117 ;
  assign n5119 = n5113 | n5115 ;
  assign n5120 = ( n5113 & ~n5118 ) | ( n5113 & n5119 ) | ( ~n5118 & n5119 );
  assign n5121 = ( n5113 & ~n5117 ) | ( n5113 & n5119 ) | ( ~n5117 & n5119 );
  assign n5122 = ( ~n4974 & n5120 ) | ( ~n4974 & n5121 ) | ( n5120 & n5121 );
  assign n5123 = ( ~n4975 & n5120 ) | ( ~n4975 & n5121 ) | ( n5120 & n5121 );
  assign n5124 = ( ~n4788 & n5122 ) | ( ~n4788 & n5123 ) | ( n5122 & n5123 );
  assign n5125 = ~n5114 & n5124 ;
  assign n5126 = ( n5052 & n5078 ) | ( n5052 & n5125 ) | ( n5078 & n5125 );
  assign n5127 = ( n5051 & n5078 ) | ( n5051 & n5125 ) | ( n5078 & n5125 );
  assign n5128 = ( n5055 & n5126 ) | ( n5055 & n5127 ) | ( n5126 & n5127 );
  assign n5129 = ( ~n5052 & n5078 ) | ( ~n5052 & n5125 ) | ( n5078 & n5125 );
  assign n5130 = ( ~n5051 & n5078 ) | ( ~n5051 & n5125 ) | ( n5078 & n5125 );
  assign n5131 = ( ~n5055 & n5129 ) | ( ~n5055 & n5130 ) | ( n5129 & n5130 );
  assign n5132 = n5052 | n5053 ;
  assign n5133 = ( n5052 & n5055 ) | ( n5052 & n5132 ) | ( n5055 & n5132 );
  assign n5134 = ( ~n5128 & n5131 ) | ( ~n5128 & n5133 ) | ( n5131 & n5133 );
  assign n5135 = n5060 | n5134 ;
  assign n5136 = n5060 & n5134 ;
  assign n5137 = n5135 & ~n5136 ;
  assign n5138 = n5061 | n5062 ;
  assign n5139 = n3803 & n5138 ;
  assign n5140 = ~n5137 & n5139 ;
  assign n5141 = n5137 & ~n5139 ;
  assign n5142 = n5140 | n5141 ;
  assign n5143 = n182 | n268 ;
  assign n5144 = n196 | n356 ;
  assign n5145 = n5143 | n5144 ;
  assign n5146 = n102 | n2000 ;
  assign n5147 = n3949 | n5146 ;
  assign n5148 = n5145 | n5147 ;
  assign n5149 = n1036 | n2062 ;
  assign n5150 = n910 | n5149 ;
  assign n5151 = n5148 | n5150 ;
  assign n5152 = n184 | n5151 ;
  assign n5153 = n3626 | n5152 ;
  assign n5154 = n200 | n344 ;
  assign n5155 = n160 | n5154 ;
  assign n5156 = n141 | n5155 ;
  assign n5157 = n387 | n5156 ;
  assign n5158 = n455 | n5157 ;
  assign n5159 = n5153 | n5158 ;
  assign n5160 = n2816 & ~n3827 ;
  assign n5161 = n2526 & n2898 ;
  assign n5162 = n2814 & ~n3682 ;
  assign n5163 = n5161 | n5162 ;
  assign n5164 = n5160 | n5163 ;
  assign n5165 = n2819 & n3843 ;
  assign n5166 = n5164 | n5165 ;
  assign n5167 = n332 & n5166 ;
  assign n5168 = n5166 & ~n5167 ;
  assign n5169 = n332 & ~n5167 ;
  assign n5170 = n5168 | n5169 ;
  assign n5171 = ~n5081 & n5082 ;
  assign n5172 = n332 & n2541 ;
  assign n5173 = ~n453 & n5079 ;
  assign n5174 = n453 & ~n5079 ;
  assign n5175 = n5173 | n5174 ;
  assign n5176 = n5172 & ~n5175 ;
  assign n5177 = ~n5172 & n5175 ;
  assign n5178 = n5176 | n5177 ;
  assign n5179 = ( n5083 & n5170 ) | ( n5083 & ~n5178 ) | ( n5170 & ~n5178 );
  assign n5180 = ( n5081 & n5170 ) | ( n5081 & ~n5178 ) | ( n5170 & ~n5178 );
  assign n5181 = ( ~n5171 & n5179 ) | ( ~n5171 & n5180 ) | ( n5179 & n5180 );
  assign n5182 = ( n5081 & n5083 ) | ( n5081 & ~n5171 ) | ( n5083 & ~n5171 );
  assign n5183 = ( n5178 & n5181 ) | ( n5178 & ~n5182 ) | ( n5181 & ~n5182 );
  assign n5184 = ( ~n5170 & n5181 ) | ( ~n5170 & n5183 ) | ( n5181 & n5183 );
  assign n5185 = ~n5086 & n5106 ;
  assign n5186 = n5104 & ~n5181 ;
  assign n5187 = n5104 & n5170 ;
  assign n5188 = ( ~n5183 & n5186 ) | ( ~n5183 & n5187 ) | ( n5186 & n5187 );
  assign n5189 = ( ~n5184 & n5185 ) | ( ~n5184 & n5188 ) | ( n5185 & n5188 );
  assign n5190 = ~n5104 & n5181 ;
  assign n5191 = n5104 | n5170 ;
  assign n5192 = ( n5183 & n5190 ) | ( n5183 & ~n5191 ) | ( n5190 & ~n5191 );
  assign n5193 = ~n5185 & n5192 ;
  assign n5194 = n5189 | n5193 ;
  assign n5195 = n5112 & ~n5194 ;
  assign n5196 = ( n5124 & n5194 ) | ( n5124 & ~n5195 ) | ( n5194 & ~n5195 );
  assign n5197 = ~n5112 & n5194 ;
  assign n5198 = n5124 & n5197 ;
  assign n5199 = n5196 & ~n5198 ;
  assign n5200 = n5159 & n5199 ;
  assign n5201 = n5159 | n5199 ;
  assign n5202 = ~n5200 & n5201 ;
  assign n5203 = n5127 & ~n5202 ;
  assign n5204 = n5126 & ~n5202 ;
  assign n5205 = ( n5055 & n5203 ) | ( n5055 & n5204 ) | ( n5203 & n5204 );
  assign n5206 = ~n5127 & n5202 ;
  assign n5207 = ~n5126 & n5202 ;
  assign n5208 = ( ~n5055 & n5206 ) | ( ~n5055 & n5207 ) | ( n5206 & n5207 );
  assign n5209 = n5205 | n5208 ;
  assign n5210 = n5134 & n5209 ;
  assign n5211 = n5060 & n5210 ;
  assign n5212 = n5134 | n5209 ;
  assign n5213 = ( n5060 & n5209 ) | ( n5060 & n5212 ) | ( n5209 & n5212 );
  assign n5214 = ~n5211 & n5213 ;
  assign n5215 = n5137 | n5138 ;
  assign n5216 = n3803 & n5215 ;
  assign n5217 = ~n5214 & n5216 ;
  assign n5218 = n5214 & ~n5216 ;
  assign n5219 = n5217 | n5218 ;
  assign n5220 = n5200 | n5202 ;
  assign n5221 = n377 | n2044 ;
  assign n5222 = n368 | n2043 ;
  assign n5223 = n2080 | n5222 ;
  assign n5224 = n5221 | n5223 ;
  assign n5225 = n272 | n1352 ;
  assign n5226 = n268 | n5225 ;
  assign n5227 = n2040 | n5226 ;
  assign n5228 = n410 | n486 ;
  assign n5229 = n210 | n5228 ;
  assign n5230 = n2243 | n2303 ;
  assign n5231 = n5229 | n5230 ;
  assign n5232 = n5227 | n5231 ;
  assign n5233 = n2336 | n3981 ;
  assign n5234 = n120 | n338 ;
  assign n5235 = n142 | n5234 ;
  assign n5236 = n5233 | n5235 ;
  assign n5237 = n5232 | n5236 ;
  assign n5238 = n2046 | n5237 ;
  assign n5239 = n136 | n2507 ;
  assign n5240 = n5238 | n5239 ;
  assign n5241 = n5224 | n5240 ;
  assign n5242 = n111 | n166 ;
  assign n5243 = n5241 | n5242 ;
  assign n5244 = n344 | n5243 ;
  assign n5245 = n355 | n5244 ;
  assign n5246 = n276 | n5245 ;
  assign n5247 = n412 | n5246 ;
  assign n5248 = n332 & n2526 ;
  assign n5249 = n5172 | n5173 ;
  assign n5250 = ( n5173 & ~n5175 ) | ( n5173 & n5249 ) | ( ~n5175 & n5249 );
  assign n5251 = n2814 & ~n3827 ;
  assign n5252 = n2813 | n3682 ;
  assign n5253 = n2897 & ~n5252 ;
  assign n5254 = n5251 | n5253 ;
  assign n5255 = n2819 & n4095 ;
  assign n5256 = n332 & ~n5255 ;
  assign n5257 = ~n5254 & n5256 ;
  assign n5258 = n332 & ~n5257 ;
  assign n5259 = ( n5248 & n5250 ) | ( n5248 & n5257 ) | ( n5250 & n5257 );
  assign n5260 = n5254 | n5255 ;
  assign n5261 = ( n5248 & n5250 ) | ( n5248 & n5260 ) | ( n5250 & n5260 );
  assign n5262 = ( ~n5258 & n5259 ) | ( ~n5258 & n5261 ) | ( n5259 & n5261 );
  assign n5263 = ( n5248 & n5250 ) | ( n5248 & ~n5262 ) | ( n5250 & ~n5262 );
  assign n5264 = n5181 & n5262 ;
  assign n5265 = ( n5257 & ~n5258 ) | ( n5257 & n5260 ) | ( ~n5258 & n5260 );
  assign n5266 = n5181 & ~n5265 ;
  assign n5267 = ( ~n5263 & n5264 ) | ( ~n5263 & n5266 ) | ( n5264 & n5266 );
  assign n5268 = n5181 | n5262 ;
  assign n5269 = ~n5181 & n5265 ;
  assign n5270 = ( n5263 & ~n5268 ) | ( n5263 & n5269 ) | ( ~n5268 & n5269 );
  assign n5271 = n5267 | n5270 ;
  assign n5272 = n5189 | n5195 ;
  assign n5273 = ~n5189 & n5194 ;
  assign n5274 = ( n5124 & ~n5272 ) | ( n5124 & n5273 ) | ( ~n5272 & n5273 );
  assign n5275 = n5271 | n5274 ;
  assign n5276 = n5271 & n5274 ;
  assign n5277 = n5275 & ~n5276 ;
  assign n5278 = n5247 | n5277 ;
  assign n5279 = n5247 & n5277 ;
  assign n5280 = n5278 & ~n5279 ;
  assign n5281 = n5126 & n5280 ;
  assign n5282 = n5200 & n5280 ;
  assign n5283 = ( n5220 & n5281 ) | ( n5220 & n5282 ) | ( n5281 & n5282 );
  assign n5284 = ( n5200 & n5202 ) | ( n5200 & n5280 ) | ( n5202 & n5280 );
  assign n5285 = ( n5127 & n5282 ) | ( n5127 & n5284 ) | ( n5282 & n5284 );
  assign n5286 = ( n5055 & n5283 ) | ( n5055 & n5285 ) | ( n5283 & n5285 );
  assign n5287 = n5220 | n5280 ;
  assign n5288 = n5200 | n5280 ;
  assign n5289 = ( n5127 & n5287 ) | ( n5127 & n5288 ) | ( n5287 & n5288 );
  assign n5290 = n5126 | n5280 ;
  assign n5291 = ( n5220 & n5288 ) | ( n5220 & n5290 ) | ( n5288 & n5290 );
  assign n5292 = ( n5055 & n5289 ) | ( n5055 & n5291 ) | ( n5289 & n5291 );
  assign n5293 = ~n5286 & n5292 ;
  assign n5294 = n5209 & n5293 ;
  assign n5295 = n5136 & n5294 ;
  assign n5296 = n5211 | n5293 ;
  assign n5297 = ~n5295 & n5296 ;
  assign n5298 = n5214 | n5215 ;
  assign n5299 = n3803 & n5298 ;
  assign n5300 = ~n5297 & n5299 ;
  assign n5301 = n5297 & ~n5299 ;
  assign n5302 = n5300 | n5301 ;
  assign n5303 = n311 | n1103 ;
  assign n5304 = n322 | n5303 ;
  assign n5305 = n1102 | n5304 ;
  assign n5306 = n195 | n5305 ;
  assign n5307 = n930 | n5306 ;
  assign n5308 = n560 | n5071 ;
  assign n5309 = ( ~n2250 & n5307 ) | ( ~n2250 & n5308 ) | ( n5307 & n5308 );
  assign n5310 = n5307 & n5308 ;
  assign n5311 = ( ~n2246 & n5309 ) | ( ~n2246 & n5310 ) | ( n5309 & n5310 );
  assign n5312 = n2251 | n5311 ;
  assign n5313 = n222 | n238 ;
  assign n5314 = n368 | n412 ;
  assign n5315 = n5313 | n5314 ;
  assign n5316 = n641 | n5315 ;
  assign n5317 = n111 | n1014 ;
  assign n5318 = n1013 | n5317 ;
  assign n5319 = n5316 | n5318 ;
  assign n5320 = n5312 | n5319 ;
  assign n5321 = n332 & ~n3685 ;
  assign n5322 = n2819 & ~n4093 ;
  assign n5323 = n2813 | n3827 ;
  assign n5324 = n2897 & ~n5323 ;
  assign n5325 = n5322 | n5324 ;
  assign n5326 = n332 & ~n5325 ;
  assign n5327 = ~n332 & n5325 ;
  assign n5328 = n5326 | n5327 ;
  assign n5329 = ~n5321 & n5328 ;
  assign n5330 = n5321 & ~n5328 ;
  assign n5331 = n5329 | n5330 ;
  assign n5332 = ( ~n5248 & n5250 ) | ( ~n5248 & n5257 ) | ( n5250 & n5257 );
  assign n5333 = ( ~n5248 & n5250 ) | ( ~n5248 & n5260 ) | ( n5250 & n5260 );
  assign n5334 = ( ~n5258 & n5332 ) | ( ~n5258 & n5333 ) | ( n5332 & n5333 );
  assign n5335 = n5331 & ~n5334 ;
  assign n5336 = ~n5331 & n5334 ;
  assign n5337 = n5335 | n5336 ;
  assign n5338 = ~n5267 & n5274 ;
  assign n5339 = ( ~n5267 & n5271 ) | ( ~n5267 & n5338 ) | ( n5271 & n5338 );
  assign n5340 = n5337 & n5339 ;
  assign n5341 = n5337 | n5339 ;
  assign n5342 = ~n5340 & n5341 ;
  assign n5343 = n5320 & n5342 ;
  assign n5344 = n5320 | n5342 ;
  assign n5345 = ~n5343 & n5344 ;
  assign n5346 = n5279 & ~n5343 ;
  assign n5347 = ( n5283 & n5345 ) | ( n5283 & n5346 ) | ( n5345 & n5346 );
  assign n5348 = n5279 & n5345 ;
  assign n5349 = ( n5284 & n5345 ) | ( n5284 & n5348 ) | ( n5345 & n5348 );
  assign n5350 = ( n5282 & n5345 ) | ( n5282 & n5348 ) | ( n5345 & n5348 );
  assign n5351 = ( n5127 & n5349 ) | ( n5127 & n5350 ) | ( n5349 & n5350 );
  assign n5352 = ( n5055 & n5347 ) | ( n5055 & n5351 ) | ( n5347 & n5351 );
  assign n5353 = n5279 | n5345 ;
  assign n5354 = n5285 | n5353 ;
  assign n5355 = n5283 | n5353 ;
  assign n5356 = ( n5055 & n5354 ) | ( n5055 & n5355 ) | ( n5354 & n5355 );
  assign n5357 = ~n5352 & n5356 ;
  assign n5358 = n5294 & n5357 ;
  assign n5359 = n5136 & n5358 ;
  assign n5360 = n5294 | n5357 ;
  assign n5361 = ( n5136 & n5357 ) | ( n5136 & n5360 ) | ( n5357 & n5360 );
  assign n5362 = ~n5359 & n5361 ;
  assign n5363 = n5297 | n5298 ;
  assign n5364 = n3803 & n5363 ;
  assign n5365 = ~n5362 & n5364 ;
  assign n5366 = n5362 & ~n5364 ;
  assign n5367 = n5365 | n5366 ;
  assign n5368 = n102 | n5145 ;
  assign n5369 = n522 | n2106 ;
  assign n5370 = n2184 | n5369 ;
  assign n5371 = n5368 | n5370 ;
  assign n5372 = n228 | n373 ;
  assign n5373 = n5371 | n5372 ;
  assign n5374 = n153 | n3629 ;
  assign n5375 = n336 | n5374 ;
  assign n5376 = n371 | n5375 ;
  assign n5377 = n5373 | n5376 ;
  assign n5378 = ~n2526 & n3827 ;
  assign n5379 = ( n332 & n2526 ) | ( n332 & n5378 ) | ( n2526 & n5378 );
  assign n5380 = ( ~n3827 & n5378 ) | ( ~n3827 & n5379 ) | ( n5378 & n5379 );
  assign n5381 = n332 & ~n3682 ;
  assign n5382 = ~n5248 & n5381 ;
  assign n5383 = n5321 & ~n5382 ;
  assign n5384 = ( n5328 & n5382 ) | ( n5328 & ~n5383 ) | ( n5382 & ~n5383 );
  assign n5385 = ( n5334 & ~n5380 ) | ( n5334 & n5384 ) | ( ~n5380 & n5384 );
  assign n5386 = ~n5380 & n5384 ;
  assign n5387 = ( ~n5331 & n5385 ) | ( ~n5331 & n5386 ) | ( n5385 & n5386 );
  assign n5388 = n5380 & ~n5384 ;
  assign n5389 = ( n5337 & ~n5387 ) | ( n5337 & n5388 ) | ( ~n5387 & n5388 );
  assign n5390 = ( n5339 & ~n5387 ) | ( n5339 & n5389 ) | ( ~n5387 & n5389 );
  assign n5391 = ~n5336 & n5337 ;
  assign n5392 = ( ~n5336 & n5339 ) | ( ~n5336 & n5391 ) | ( n5339 & n5391 );
  assign n5393 = ( n5384 & n5390 ) | ( n5384 & ~n5392 ) | ( n5390 & ~n5392 );
  assign n5394 = ( ~n5380 & n5390 ) | ( ~n5380 & n5393 ) | ( n5390 & n5393 );
  assign n5395 = n5377 & n5394 ;
  assign n5396 = n5377 | n5394 ;
  assign n5397 = n5343 & n5396 ;
  assign n5398 = ~n5395 & n5397 ;
  assign n5399 = ~n5395 & n5396 ;
  assign n5400 = ( n5351 & n5398 ) | ( n5351 & n5399 ) | ( n5398 & n5399 );
  assign n5401 = ( n5346 & n5398 ) | ( n5346 & n5399 ) | ( n5398 & n5399 );
  assign n5402 = ( n5345 & n5398 ) | ( n5345 & n5399 ) | ( n5398 & n5399 );
  assign n5403 = ( n5283 & n5401 ) | ( n5283 & n5402 ) | ( n5401 & n5402 );
  assign n5404 = ( n5055 & n5400 ) | ( n5055 & n5403 ) | ( n5400 & n5403 );
  assign n5405 = n5343 | n5351 ;
  assign n5406 = n5343 | n5346 ;
  assign n5407 = ( n5283 & n5344 ) | ( n5283 & n5406 ) | ( n5344 & n5406 );
  assign n5408 = ( n5055 & n5405 ) | ( n5055 & n5407 ) | ( n5405 & n5407 );
  assign n5409 = ~n5404 & n5408 ;
  assign n5410 = ~n5397 & n5399 ;
  assign n5411 = ~n5351 & n5410 ;
  assign n5412 = ~n5346 & n5410 ;
  assign n5413 = ~n5345 & n5410 ;
  assign n5414 = ( ~n5283 & n5412 ) | ( ~n5283 & n5413 ) | ( n5412 & n5413 );
  assign n5415 = ( ~n5055 & n5411 ) | ( ~n5055 & n5414 ) | ( n5411 & n5414 );
  assign n5416 = n5409 | n5415 ;
  assign n5417 = n5357 & n5416 ;
  assign n5418 = n5295 & n5417 ;
  assign n5419 = n5359 | n5416 ;
  assign n5420 = ~n5418 & n5419 ;
  assign n5421 = ( n3803 & n5362 ) | ( n3803 & n5364 ) | ( n5362 & n5364 );
  assign n5422 = ~n5420 & n5421 ;
  assign n5423 = n5420 & ~n5421 ;
  assign n5424 = n5422 | n5423 ;
  assign n5425 = n5362 | n5420 ;
  assign n5426 = n5363 | n5425 ;
  assign n5427 = n3803 & n5426 ;
  assign n5428 = n133 | n2000 ;
  assign n5429 = n845 | n5428 ;
  assign n5430 = n334 | n2459 ;
  assign n5431 = n207 | n411 ;
  assign n5432 = n5430 | n5431 ;
  assign n5433 = n89 | n338 ;
  assign n5434 = n279 | n370 ;
  assign n5435 = n5433 | n5434 ;
  assign n5436 = n5432 | n5435 ;
  assign n5437 = n5429 | n5436 ;
  assign n5438 = n202 | n504 ;
  assign n5439 = n122 | n910 ;
  assign n5440 = n149 | n5439 ;
  assign n5441 = n5438 | n5440 ;
  assign n5442 = n5437 | n5441 ;
  assign n5443 = n116 | n5442 ;
  assign n5444 = n237 | n5443 ;
  assign n5445 = n5395 & n5444 ;
  assign n5446 = ( n5397 & n5444 ) | ( n5397 & n5445 ) | ( n5444 & n5445 );
  assign n5447 = ( n5399 & n5444 ) | ( n5399 & n5445 ) | ( n5444 & n5445 );
  assign n5448 = ( n5351 & n5446 ) | ( n5351 & n5447 ) | ( n5446 & n5447 );
  assign n5449 = ( n5346 & n5446 ) | ( n5346 & n5447 ) | ( n5446 & n5447 );
  assign n5450 = ( n5345 & n5446 ) | ( n5345 & n5447 ) | ( n5446 & n5447 );
  assign n5451 = ( n5283 & n5449 ) | ( n5283 & n5450 ) | ( n5449 & n5450 );
  assign n5452 = ( n5055 & n5448 ) | ( n5055 & n5451 ) | ( n5448 & n5451 );
  assign n5453 = n5395 | n5444 ;
  assign n5454 = n5397 | n5453 ;
  assign n5455 = n5399 | n5453 ;
  assign n5456 = ( n5351 & n5454 ) | ( n5351 & n5455 ) | ( n5454 & n5455 );
  assign n5457 = ( n5346 & n5454 ) | ( n5346 & n5455 ) | ( n5454 & n5455 );
  assign n5458 = ( n5345 & n5454 ) | ( n5345 & n5455 ) | ( n5454 & n5455 );
  assign n5459 = ( n5283 & n5457 ) | ( n5283 & n5458 ) | ( n5457 & n5458 );
  assign n5460 = ( n5055 & n5456 ) | ( n5055 & n5459 ) | ( n5456 & n5459 );
  assign n5461 = ~n5452 & n5460 ;
  assign n5462 = n5357 & ~n5461 ;
  assign n5463 = n5416 & n5462 ;
  assign n5464 = n5295 & n5463 ;
  assign n5465 = n5461 | n5463 ;
  assign n5466 = ( n5295 & n5461 ) | ( n5295 & n5465 ) | ( n5461 & n5465 );
  assign n5467 = ( ~n5418 & n5464 ) | ( ~n5418 & n5466 ) | ( n5464 & n5466 );
  assign n5468 = n5427 & n5467 ;
  assign n5469 = n5427 | n5467 ;
  assign n5470 = ~n5468 & n5469 ;
  assign n5471 = n5426 | n5467 ;
  assign n5472 = n3803 & n5471 ;
  assign n5473 = n149 | n413 ;
  assign n5474 = n215 | n5473 ;
  assign n5475 = n370 | n474 ;
  assign n5476 = n2053 | n5475 ;
  assign n5477 = n562 | n5476 ;
  assign n5478 = n1065 | n5477 ;
  assign n5479 = n1019 | n5478 ;
  assign n5480 = n908 | n5479 ;
  assign n5481 = n166 | n5480 ;
  assign n5482 = n218 | n5481 ;
  assign n5483 = ( ~n3583 & n3585 ) | ( ~n3583 & n5482 ) | ( n3585 & n5482 );
  assign n5484 = n3583 | n5483 ;
  assign n5485 = n5474 | n5484 ;
  assign n5486 = n5446 | n5485 ;
  assign n5487 = n5447 | n5485 ;
  assign n5488 = ( n5351 & n5486 ) | ( n5351 & n5487 ) | ( n5486 & n5487 );
  assign n5489 = ( n5347 & n5486 ) | ( n5347 & n5487 ) | ( n5486 & n5487 );
  assign n5490 = ( n5055 & n5488 ) | ( n5055 & n5489 ) | ( n5488 & n5489 );
  assign n5491 = n5446 & n5485 ;
  assign n5492 = n5447 & n5485 ;
  assign n5493 = ( n5351 & n5491 ) | ( n5351 & n5492 ) | ( n5491 & n5492 );
  assign n5494 = ( n5347 & n5491 ) | ( n5347 & n5492 ) | ( n5491 & n5492 );
  assign n5495 = ( n5055 & n5493 ) | ( n5055 & n5494 ) | ( n5493 & n5494 );
  assign n5496 = n5490 & ~n5495 ;
  assign n5497 = n5461 | n5496 ;
  assign n5498 = ( n5417 & n5496 ) | ( n5417 & n5497 ) | ( n5496 & n5497 );
  assign n5499 = n5496 & n5497 ;
  assign n5500 = ( n5295 & n5498 ) | ( n5295 & n5499 ) | ( n5498 & n5499 );
  assign n5501 = n5461 & n5490 ;
  assign n5502 = n5500 & ~n5501 ;
  assign n5503 = ( ~n5418 & n5500 ) | ( ~n5418 & n5502 ) | ( n5500 & n5502 );
  assign n5504 = n5472 & ~n5503 ;
  assign n5505 = ~n5472 & n5503 ;
  assign n5506 = n5504 | n5505 ;
  assign n5507 = n5467 | n5503 ;
  assign n5508 = n5426 | n5507 ;
  assign n5509 = n3803 & n5508 ;
  assign n5510 = n5294 & n5501 ;
  assign n5511 = n5136 & n5510 ;
  assign n5512 = n195 | n4400 ;
  assign n5513 = n529 | n5512 ;
  assign n5514 = n5305 | n5513 ;
  assign n5515 = n115 | n870 ;
  assign n5516 = n2431 | n5515 ;
  assign n5517 = n5514 | n5516 ;
  assign n5518 = n128 | n132 ;
  assign n5519 = n153 | n5518 ;
  assign n5520 = n123 | n5519 ;
  assign n5521 = n335 | n5520 ;
  assign n5522 = n410 | n5521 ;
  assign n5523 = n152 | n5522 ;
  assign n5524 = n5517 | n5523 ;
  assign n5525 = n5485 & n5524 ;
  assign n5526 = n5446 & n5525 ;
  assign n5527 = n5447 & n5525 ;
  assign n5528 = ( n5351 & n5526 ) | ( n5351 & n5527 ) | ( n5526 & n5527 );
  assign n5529 = ( n5347 & n5526 ) | ( n5347 & n5527 ) | ( n5526 & n5527 );
  assign n5530 = ( n5055 & n5528 ) | ( n5055 & n5529 ) | ( n5528 & n5529 );
  assign n5531 = n5485 | n5524 ;
  assign n5532 = ( n5446 & n5524 ) | ( n5446 & n5531 ) | ( n5524 & n5531 );
  assign n5533 = ( n5447 & n5524 ) | ( n5447 & n5531 ) | ( n5524 & n5531 );
  assign n5534 = ( n5351 & n5532 ) | ( n5351 & n5533 ) | ( n5532 & n5533 );
  assign n5535 = ( n5347 & n5532 ) | ( n5347 & n5533 ) | ( n5532 & n5533 );
  assign n5536 = ( n5055 & n5534 ) | ( n5055 & n5535 ) | ( n5534 & n5535 );
  assign n5537 = ~n5530 & n5536 ;
  assign n5538 = ~n5417 & n5511 ;
  assign n5539 = ( n5511 & n5537 ) | ( n5511 & n5538 ) | ( n5537 & n5538 );
  assign n5540 = ( n5537 & n5538 ) | ( n5537 & ~n5539 ) | ( n5538 & ~n5539 );
  assign n5541 = ( n5511 & ~n5539 ) | ( n5511 & n5540 ) | ( ~n5539 & n5540 );
  assign n5542 = n5509 & ~n5541 ;
  assign n5543 = ~n5509 & n5541 ;
  assign n5544 = n5542 | n5543 ;
  assign n5545 = n5417 & n5501 ;
  assign n5546 = n179 | n351 ;
  assign n5547 = n408 | n4725 ;
  assign n5548 = n182 | n2002 ;
  assign n5549 = n5547 | n5548 ;
  assign n5550 = n218 | n298 ;
  assign n5551 = n5549 | n5550 ;
  assign n5552 = ( ~n925 & n5546 ) | ( ~n925 & n5551 ) | ( n5546 & n5551 );
  assign n5553 = n206 | n233 ;
  assign n5554 = n205 | n5553 ;
  assign n5555 = n925 | n5554 ;
  assign n5556 = n5552 | n5555 ;
  assign n5557 = n5525 | n5556 ;
  assign n5558 = ( n5446 & n5556 ) | ( n5446 & n5557 ) | ( n5556 & n5557 );
  assign n5559 = n487 | n5558 ;
  assign n5560 = ( n5447 & n5556 ) | ( n5447 & n5557 ) | ( n5556 & n5557 );
  assign n5561 = n487 | n5560 ;
  assign n5562 = ( n5351 & n5559 ) | ( n5351 & n5561 ) | ( n5559 & n5561 );
  assign n5563 = ( n5347 & n5559 ) | ( n5347 & n5561 ) | ( n5559 & n5561 );
  assign n5564 = ( n5055 & n5562 ) | ( n5055 & n5563 ) | ( n5562 & n5563 );
  assign n5565 = ( ~n5501 & n5537 ) | ( ~n5501 & n5564 ) | ( n5537 & n5564 );
  assign n5566 = n5537 | n5564 ;
  assign n5567 = ( ~n5417 & n5565 ) | ( ~n5417 & n5566 ) | ( n5565 & n5566 );
  assign n5568 = n5545 & n5567 ;
  assign n5569 = n5295 & n5568 ;
  assign n5570 = n5525 & n5556 ;
  assign n5571 = n5447 & n5570 ;
  assign n5572 = ( n487 & n5527 ) | ( n487 & n5571 ) | ( n5527 & n5571 );
  assign n5573 = n5446 & n5570 ;
  assign n5574 = ( n487 & n5526 ) | ( n487 & n5573 ) | ( n5526 & n5573 );
  assign n5575 = ( n5351 & n5572 ) | ( n5351 & n5574 ) | ( n5572 & n5574 );
  assign n5576 = ( n5347 & n5572 ) | ( n5347 & n5574 ) | ( n5572 & n5574 );
  assign n5577 = ( n5055 & n5575 ) | ( n5055 & n5576 ) | ( n5575 & n5576 );
  assign n5578 = n5564 & ~n5577 ;
  assign n5579 = n5537 | n5578 ;
  assign n5580 = ( n5501 & n5578 ) | ( n5501 & n5579 ) | ( n5578 & n5579 );
  assign n5581 = ( ~n5295 & n5417 ) | ( ~n5295 & n5580 ) | ( n5417 & n5580 );
  assign n5582 = ( n5295 & n5578 ) | ( n5295 & n5581 ) | ( n5578 & n5581 );
  assign n5583 = ~n5569 & n5582 ;
  assign n5584 = n5508 | n5541 ;
  assign n5585 = n3803 & n5584 ;
  assign n5586 = ~n5583 & n5585 ;
  assign n5587 = n5583 & ~n5585 ;
  assign n5588 = n5586 | n5587 ;
  assign n5589 = ( ~n269 & n391 ) | ( ~n269 & n2516 ) | ( n391 & n2516 );
  assign n5590 = n391 & n2516 ;
  assign n5591 = ( ~n326 & n5589 ) | ( ~n326 & n5590 ) | ( n5589 & n5590 );
  assign n5592 = n327 | n5591 ;
  assign n5593 = n344 | n5592 ;
  assign n5594 = n356 | n5593 ;
  assign n5595 = n5572 & n5594 ;
  assign n5596 = n5574 & n5594 ;
  assign n5597 = ( n5351 & n5595 ) | ( n5351 & n5596 ) | ( n5595 & n5596 );
  assign n5598 = ( n5347 & n5595 ) | ( n5347 & n5596 ) | ( n5595 & n5596 );
  assign n5599 = ( n5055 & n5597 ) | ( n5055 & n5598 ) | ( n5597 & n5598 );
  assign n5600 = n5572 | n5594 ;
  assign n5601 = n5574 | n5594 ;
  assign n5602 = ( n5351 & n5600 ) | ( n5351 & n5601 ) | ( n5600 & n5601 );
  assign n5603 = ( n5347 & n5600 ) | ( n5347 & n5601 ) | ( n5600 & n5601 );
  assign n5604 = ( n5055 & n5602 ) | ( n5055 & n5603 ) | ( n5602 & n5603 );
  assign n5605 = ~n5599 & n5604 ;
  assign n5606 = n5294 & n5605 ;
  assign n5607 = n5136 & n5606 ;
  assign n5608 = n5568 & n5607 ;
  assign n5609 = n5294 | n5605 ;
  assign n5610 = ( n5136 & n5605 ) | ( n5136 & n5609 ) | ( n5605 & n5609 );
  assign n5611 = ( n5568 & n5605 ) | ( n5568 & n5610 ) | ( n5605 & n5610 );
  assign n5612 = ~n5608 & n5611 ;
  assign n5613 = n5541 | n5583 ;
  assign n5614 = ( n3803 & n5509 ) | ( n3803 & n5613 ) | ( n5509 & n5613 );
  assign n5615 = ~n5612 & n5614 ;
  assign n5616 = n5612 & ~n5614 ;
  assign n5617 = n5615 | n5616 ;
  assign n5618 = n5583 | n5612 ;
  assign n5619 = n5541 | n5618 ;
  assign n5620 = ( n3803 & n5509 ) | ( n3803 & n5619 ) | ( n5509 & n5619 );
  assign n5621 = n327 | n427 ;
  assign n5622 = n5573 | n5621 ;
  assign n5623 = n5526 | n5621 ;
  assign n5624 = ( n487 & n5622 ) | ( n487 & n5623 ) | ( n5622 & n5623 );
  assign n5625 = ( n5594 & n5621 ) | ( n5594 & n5624 ) | ( n5621 & n5624 );
  assign n5626 = n5571 | n5621 ;
  assign n5627 = n5527 | n5621 ;
  assign n5628 = ( n487 & n5626 ) | ( n487 & n5627 ) | ( n5626 & n5627 );
  assign n5629 = ( n5594 & n5621 ) | ( n5594 & n5628 ) | ( n5621 & n5628 );
  assign n5630 = ( n5351 & n5625 ) | ( n5351 & n5629 ) | ( n5625 & n5629 );
  assign n5631 = ( n5347 & n5625 ) | ( n5347 & n5629 ) | ( n5625 & n5629 );
  assign n5632 = ( n5055 & n5630 ) | ( n5055 & n5631 ) | ( n5630 & n5631 );
  assign n5633 = n5607 & n5632 ;
  assign n5634 = ( ~n5568 & n5607 ) | ( ~n5568 & n5633 ) | ( n5607 & n5633 );
  assign n5635 = n5573 & n5621 ;
  assign n5636 = n5526 & n5621 ;
  assign n5637 = ( n487 & n5635 ) | ( n487 & n5636 ) | ( n5635 & n5636 );
  assign n5638 = n5594 & n5637 ;
  assign n5639 = n5571 & n5621 ;
  assign n5640 = n5527 & n5621 ;
  assign n5641 = ( n487 & n5639 ) | ( n487 & n5640 ) | ( n5639 & n5640 );
  assign n5642 = n5594 & n5641 ;
  assign n5643 = ( n5351 & n5638 ) | ( n5351 & n5642 ) | ( n5638 & n5642 );
  assign n5644 = ( n5347 & n5638 ) | ( n5347 & n5642 ) | ( n5638 & n5642 );
  assign n5645 = ( n5055 & n5643 ) | ( n5055 & n5644 ) | ( n5643 & n5644 );
  assign n5646 = n5632 & ~n5645 ;
  assign n5647 = ~n5607 & n5646 ;
  assign n5648 = ( ~n5568 & n5646 ) | ( ~n5568 & n5647 ) | ( n5646 & n5647 );
  assign n5649 = ( n5607 & ~n5634 ) | ( n5607 & n5648 ) | ( ~n5634 & n5648 );
  assign n5650 = n5620 & ~n5649 ;
  assign n5651 = ~n5620 & n5649 ;
  assign n5652 = n5650 | n5651 ;
  assign n5653 = n5632 | n5645 ;
  assign n5654 = ( ~n5607 & n5632 ) | ( ~n5607 & n5645 ) | ( n5632 & n5645 );
  assign n5655 = ( ~n5568 & n5653 ) | ( ~n5568 & n5654 ) | ( n5653 & n5654 );
  assign n5656 = n5608 & n5655 ;
  assign n5657 = ( n5607 & n5645 ) | ( n5607 & n5653 ) | ( n5645 & n5653 );
  assign n5658 = n5645 & n5653 ;
  assign n5659 = ( n5568 & n5657 ) | ( n5568 & n5658 ) | ( n5657 & n5658 );
  assign n5660 = ~n5656 & n5659 ;
  assign n5661 = n5619 | n5649 ;
  assign n5662 = ( n3803 & n5509 ) | ( n3803 & n5661 ) | ( n5509 & n5661 );
  assign n5663 = n5660 & n5662 ;
  assign n5664 = n44 | n46 ;
  assign n5665 = ( ~n5662 & n5663 ) | ( ~n5662 & n5664 ) | ( n5663 & n5664 );
  assign n5666 = ( ~n5660 & n5663 ) | ( ~n5660 & n5665 ) | ( n5663 & n5665 );
  assign n5667 = ~n46 & n3803 ;
  assign n5668 = ~n44 & n5667 ;
  assign n5669 = ~n5508 & n5659 ;
  assign n5670 = ( ~n5508 & n5661 ) | ( ~n5508 & n5669 ) | ( n5661 & n5669 );
  assign n5671 = n5508 & n5656 ;
  assign n5672 = ( n5656 & n5661 ) | ( n5656 & n5671 ) | ( n5661 & n5671 );
  assign n5673 = ( n5508 & n5670 ) | ( n5508 & ~n5672 ) | ( n5670 & ~n5672 );
  assign n5674 = ( n3803 & n5668 ) | ( n3803 & n5673 ) | ( n5668 & n5673 );
  assign po0 = n3800 ;
  assign po1 = n3975 ;
  assign po2 = n4116 ;
  assign po3 = n4252 ;
  assign po4 = n4393 ;
  assign po5 = n4499 ;
  assign po6 = n4604 ;
  assign po7 = n4710 ;
  assign po8 = n4805 ;
  assign po9 = n4901 ;
  assign po10 = n4997 ;
  assign po11 = n5066 ;
  assign po12 = n5142 ;
  assign po13 = n5219 ;
  assign po14 = n5302 ;
  assign po15 = n5367 ;
  assign po16 = n5424 ;
  assign po17 = n5470 ;
  assign po18 = n5506 ;
  assign po19 = n5544 ;
  assign po20 = n5588 ;
  assign po21 = n5617 ;
  assign po22 = n5652 ;
  assign po23 = ~n5666 ;
  assign po24 = n5674 ;
endmodule
