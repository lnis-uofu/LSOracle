module top(G1 , G5 , G9 , G13 , G33 , G41 , G17 , G18 , G19 , G20 , G21 , G22 , G23 , G24 , G4 , G8 , G12 , G16 , G36 , G29 , G30 , G31 , G32 , G3 , G7 , G11 , G15 , G35 , G25 , G26 , G27 , G28 , G2 , G6 , G10 , G14 , G34 , G40 , G39 , G38 , G37 , G1324 , G1344 , G1325 , G1326 , G1327 , G1328 , G1329 , G1330 , G1343 , G1331 , G1332 , G1333 , G1334 , G1335 , G1336 , G1337 , G1338 , G1339 , G1340 , G1341 , G1342 , G1345 , G1346 , G1347 , G1348 , G1349 , G1350 , G1351 , G1352 , G1353 , G1354 , G1355 );
  input G1 , G5 , G9 , G13 , G33 , G41 , G17 , G18 , G19 , G20 , G21 , G22 , G23 , G24 , G4 , G8 , G12 , G16 , G36 , G29 , G30 , G31 , G32 , G3 , G7 , G11 , G15 , G35 , G25 , G26 , G27 , G28 , G2 , G6 , G10 , G14 , G34 , G40 , G39 , G38 , G37 ;
  output G1324 , G1344 , G1325 , G1326 , G1327 , G1328 , G1329 , G1330 , G1343 , G1331 , G1332 , G1333 , G1334 , G1335 , G1336 , G1337 , G1338 , G1339 , G1340 , G1341 , G1342 , G1345 , G1346 , G1347 , G1348 , G1349 , G1350 , G1351 , G1352 , G1353 , G1354 , G1355 ;
  wire n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452;
  assign n42 = ~G1 & G9 ;
  assign n43 = G1 & ~G9 ;
  assign n44 = n42 | n43 ;
  assign n45 = G5 | n44 ;
  assign n46 = G5 & n44 ;
  assign n47 = n45 & ~n46 ;
  assign n48 = ~G13 & n47 ;
  assign n49 = G13 & ~n47 ;
  assign n50 = n48 | n49 ;
  assign n51 = G33 & G41 ;
  assign n52 = ~G17 & G19 ;
  assign n53 = G17 & ~G19 ;
  assign n54 = n52 | n53 ;
  assign n55 = G18 | n54 ;
  assign n56 = G18 & n54 ;
  assign n57 = n55 & ~n56 ;
  assign n58 = ~G20 & n57 ;
  assign n59 = G20 & ~n57 ;
  assign n60 = n58 | n59 ;
  assign n61 = n51 & n60 ;
  assign n62 = n51 | n60 ;
  assign n63 = ~n61 & n62 ;
  assign n64 = ~G21 & G23 ;
  assign n65 = G21 & ~G23 ;
  assign n66 = n64 | n65 ;
  assign n67 = G22 | n66 ;
  assign n68 = G22 & n66 ;
  assign n69 = n67 & ~n68 ;
  assign n70 = ~G24 & n69 ;
  assign n71 = G24 & ~n69 ;
  assign n72 = n70 | n71 ;
  assign n73 = n63 & n72 ;
  assign n74 = n63 | n72 ;
  assign n75 = ~n73 & n74 ;
  assign n76 = n50 & n75 ;
  assign n77 = n50 & ~n76 ;
  assign n78 = n75 & ~n76 ;
  assign n79 = n77 | n78 ;
  assign n80 = ~G16 & G15 ;
  assign n81 = G16 & ~G15 ;
  assign n82 = n80 | n81 ;
  assign n83 = ~G13 & G14 ;
  assign n84 = G13 & ~G14 ;
  assign n85 = n83 | n84 ;
  assign n86 = n82 & ~n85 ;
  assign n87 = ~n82 & n85 ;
  assign n88 = n86 | n87 ;
  assign n89 = ~G9 & G11 ;
  assign n90 = G9 & ~G11 ;
  assign n91 = n89 | n90 ;
  assign n92 = G12 | n91 ;
  assign n93 = G12 & n91 ;
  assign n94 = n92 & ~n93 ;
  assign n95 = ~G10 & n94 ;
  assign n96 = G10 & ~n94 ;
  assign n97 = n95 | n96 ;
  assign n98 = G41 & G38 ;
  assign n99 = ~G18 & G30 ;
  assign n100 = G18 & ~G30 ;
  assign n101 = n99 | n100 ;
  assign n102 = G22 | n101 ;
  assign n103 = G22 & n101 ;
  assign n104 = n102 & ~n103 ;
  assign n105 = ~G26 & n104 ;
  assign n106 = G26 & ~n104 ;
  assign n107 = n105 | n106 ;
  assign n108 = n98 & n107 ;
  assign n109 = n98 | n107 ;
  assign n110 = ~n108 & n109 ;
  assign n111 = n97 & n110 ;
  assign n112 = n97 | n110 ;
  assign n113 = ~n111 & n112 ;
  assign n114 = ~n88 & n113 ;
  assign n115 = n88 & ~n113 ;
  assign n116 = n114 | n115 ;
  assign n117 = ~G20 & G24 ;
  assign n118 = G20 & ~G24 ;
  assign n119 = n117 | n118 ;
  assign n120 = ~G5 & G6 ;
  assign n121 = G5 & ~G6 ;
  assign n122 = n120 | n121 ;
  assign n123 = ~G8 & G7 ;
  assign n124 = G8 & ~G7 ;
  assign n125 = n123 | n124 ;
  assign n126 = n122 & ~n125 ;
  assign n127 = ~n122 & n125 ;
  assign n128 = n126 | n127 ;
  assign n129 = G41 & G40 ;
  assign n130 = n88 & n129 ;
  assign n131 = n88 | n129 ;
  assign n132 = ~n130 & n131 ;
  assign n133 = ~n128 & n132 ;
  assign n134 = n128 & ~n132 ;
  assign n135 = n133 | n134 ;
  assign n136 = ~G32 & G28 ;
  assign n137 = G32 & ~G28 ;
  assign n138 = n136 | n137 ;
  assign n139 = n135 & ~n138 ;
  assign n140 = ~n135 & n138 ;
  assign n141 = n139 | n140 ;
  assign n142 = n119 & ~n141 ;
  assign n143 = ~n119 & n141 ;
  assign n144 = n142 | n143 ;
  assign n145 = n116 | n144 ;
  assign n146 = ~G19 & G23 ;
  assign n147 = G19 & ~G23 ;
  assign n148 = n146 | n147 ;
  assign n149 = G41 & G39 ;
  assign n150 = ~G1 & G2 ;
  assign n151 = G1 & ~G2 ;
  assign n152 = n150 | n151 ;
  assign n153 = ~G4 & G3 ;
  assign n154 = G4 & ~G3 ;
  assign n155 = n153 | n154 ;
  assign n156 = n152 & ~n155 ;
  assign n157 = ~n152 & n155 ;
  assign n158 = n156 | n157 ;
  assign n159 = n97 | n158 ;
  assign n160 = n97 & n158 ;
  assign n161 = n159 & ~n160 ;
  assign n162 = n149 | n161 ;
  assign n163 = n149 & n161 ;
  assign n164 = n162 & ~n163 ;
  assign n165 = ~G31 & G27 ;
  assign n166 = G31 & ~G27 ;
  assign n167 = n165 | n166 ;
  assign n168 = n164 & ~n167 ;
  assign n169 = ~n164 & n167 ;
  assign n170 = n168 | n169 ;
  assign n171 = n148 & ~n170 ;
  assign n172 = ~n148 & n170 ;
  assign n173 = n171 | n172 ;
  assign n174 = ~G17 & G21 ;
  assign n175 = G17 & ~G21 ;
  assign n176 = n174 | n175 ;
  assign n177 = G41 & G37 ;
  assign n178 = n128 & ~n158 ;
  assign n179 = ~n128 & n158 ;
  assign n180 = n178 | n179 ;
  assign n181 = n177 | n180 ;
  assign n182 = n177 & n180 ;
  assign n183 = n181 & ~n182 ;
  assign n184 = ~G29 & G25 ;
  assign n185 = G29 & ~G25 ;
  assign n186 = n184 | n185 ;
  assign n187 = n183 & ~n186 ;
  assign n188 = ~n183 & n186 ;
  assign n189 = n187 | n188 ;
  assign n190 = n176 & ~n189 ;
  assign n191 = ~n176 & n189 ;
  assign n192 = n190 | n191 ;
  assign n193 = n173 & n192 ;
  assign n194 = ~G3 & G11 ;
  assign n195 = G3 & ~G11 ;
  assign n196 = n194 | n195 ;
  assign n197 = G7 | n196 ;
  assign n198 = G7 & n196 ;
  assign n199 = n197 & ~n198 ;
  assign n200 = ~G15 & n199 ;
  assign n201 = G15 & ~n199 ;
  assign n202 = n200 | n201 ;
  assign n203 = G41 & G35 ;
  assign n204 = n60 & n203 ;
  assign n205 = n60 | n203 ;
  assign n206 = ~n204 & n205 ;
  assign n207 = ~G25 & G27 ;
  assign n208 = G25 & ~G27 ;
  assign n209 = n207 | n208 ;
  assign n210 = G26 | n209 ;
  assign n211 = G26 & n209 ;
  assign n212 = n210 & ~n211 ;
  assign n213 = ~G28 & n212 ;
  assign n214 = G28 & ~n212 ;
  assign n215 = n213 | n214 ;
  assign n216 = n206 & n215 ;
  assign n217 = n206 | n215 ;
  assign n218 = ~n216 & n217 ;
  assign n219 = n202 & n218 ;
  assign n220 = n202 & ~n219 ;
  assign n221 = n218 & ~n219 ;
  assign n222 = n220 | n221 ;
  assign n223 = G41 & G36 ;
  assign n224 = n72 & n223 ;
  assign n225 = n72 | n223 ;
  assign n226 = ~n224 & n225 ;
  assign n227 = ~G29 & G31 ;
  assign n228 = G29 & ~G31 ;
  assign n229 = n227 | n228 ;
  assign n230 = G30 | n229 ;
  assign n231 = G30 & n229 ;
  assign n232 = n230 & ~n231 ;
  assign n233 = ~G32 & n232 ;
  assign n234 = G32 & ~n232 ;
  assign n235 = n233 | n234 ;
  assign n236 = n226 & n235 ;
  assign n237 = n226 | n235 ;
  assign n238 = ~n236 & n237 ;
  assign n239 = ~G4 & G16 ;
  assign n240 = G4 & ~G16 ;
  assign n241 = n239 | n240 ;
  assign n242 = G8 | n241 ;
  assign n243 = G8 & n241 ;
  assign n244 = n242 & ~n243 ;
  assign n245 = ~G12 & n244 ;
  assign n246 = G12 & ~n244 ;
  assign n247 = n245 | n246 ;
  assign n248 = n238 & n247 ;
  assign n249 = n238 | n247 ;
  assign n250 = ~n248 & n249 ;
  assign n251 = n222 & ~n250 ;
  assign n252 = ~n222 & n250 ;
  assign n253 = n251 | n252 ;
  assign n254 = ~n215 & n235 ;
  assign n255 = n215 & ~n235 ;
  assign n256 = n254 | n255 ;
  assign n257 = G41 & G34 ;
  assign n258 = ~G2 & G14 ;
  assign n259 = G2 & ~G14 ;
  assign n260 = n258 | n259 ;
  assign n261 = ~G6 & G10 ;
  assign n262 = G6 & ~G10 ;
  assign n263 = n261 | n262 ;
  assign n264 = n260 & ~n263 ;
  assign n265 = ~n260 & n263 ;
  assign n266 = n264 | n265 ;
  assign n267 = n257 | n266 ;
  assign n268 = n257 & n266 ;
  assign n269 = n267 & ~n268 ;
  assign n270 = n256 & n269 ;
  assign n271 = n256 | n269 ;
  assign n272 = ~n270 & n271 ;
  assign n273 = n79 | n272 ;
  assign n274 = n253 & ~n273 ;
  assign n275 = n79 & ~n272 ;
  assign n276 = ~n79 & n272 ;
  assign n277 = n275 | n276 ;
  assign n278 = n222 | n250 ;
  assign n279 = n277 & ~n278 ;
  assign n280 = n274 | n279 ;
  assign n281 = n193 & n280 ;
  assign n282 = ~n145 & n281 ;
  assign n283 = n79 & n282 ;
  assign n284 = G1 | n283 ;
  assign n285 = G1 & n283 ;
  assign n286 = n284 & ~n285 ;
  assign n287 = n116 & n144 ;
  assign n288 = n193 | n287 ;
  assign n289 = n173 | n192 ;
  assign n290 = ~n145 & n289 ;
  assign n291 = n145 & ~n289 ;
  assign n292 = n290 | n291 ;
  assign n293 = ~n288 & n292 ;
  assign n294 = n275 & n293 ;
  assign n295 = n252 & n294 ;
  assign n296 = n192 & n295 ;
  assign n297 = G21 | n296 ;
  assign n298 = G21 & n295 ;
  assign n299 = n192 & n298 ;
  assign n300 = n297 & ~n299 ;
  assign n301 = n272 & n282 ;
  assign n302 = ~G2 & n301 ;
  assign n303 = G2 & ~n301 ;
  assign n304 = n302 | n303 ;
  assign n305 = n222 & n282 ;
  assign n306 = G3 | n305 ;
  assign n307 = G3 & n305 ;
  assign n308 = n306 & ~n307 ;
  assign n309 = n250 & n282 ;
  assign n310 = ~G4 & n309 ;
  assign n311 = G4 & ~n309 ;
  assign n312 = n310 | n311 ;
  assign n313 = n144 & ~n173 ;
  assign n314 = n192 & n313 ;
  assign n315 = ~n115 & n314 ;
  assign n316 = ~n114 & n315 ;
  assign n317 = n280 & n316 ;
  assign n318 = n79 & n317 ;
  assign n319 = G5 | n318 ;
  assign n320 = G5 & n318 ;
  assign n321 = n319 & ~n320 ;
  assign n322 = n272 & n317 ;
  assign n323 = ~G6 & n322 ;
  assign n324 = G6 & ~n322 ;
  assign n325 = n323 | n324 ;
  assign n326 = n222 & n317 ;
  assign n327 = G7 | n326 ;
  assign n328 = G7 & n326 ;
  assign n329 = n327 & ~n328 ;
  assign n330 = n251 & n294 ;
  assign n331 = n144 & n330 ;
  assign n332 = G20 | n331 ;
  assign n333 = G20 & n330 ;
  assign n334 = n144 & n333 ;
  assign n335 = n332 & ~n334 ;
  assign n336 = n250 & n317 ;
  assign n337 = ~G8 & n336 ;
  assign n338 = G8 & ~n336 ;
  assign n339 = n337 | n338 ;
  assign n340 = n144 | n192 ;
  assign n341 = n173 & ~n340 ;
  assign n342 = n116 & n341 ;
  assign n343 = n280 & n342 ;
  assign n344 = n79 & n343 ;
  assign n345 = G9 | n344 ;
  assign n346 = G9 & n344 ;
  assign n347 = n345 & ~n346 ;
  assign n348 = n272 & n343 ;
  assign n349 = ~G10 & n348 ;
  assign n350 = G10 & ~n348 ;
  assign n351 = n349 | n350 ;
  assign n352 = n222 & n343 ;
  assign n353 = G11 | n352 ;
  assign n354 = G11 & n352 ;
  assign n355 = n353 & ~n354 ;
  assign n356 = n250 & n343 ;
  assign n357 = ~G12 & n356 ;
  assign n358 = G12 & ~n356 ;
  assign n359 = n357 | n358 ;
  assign n360 = n144 & ~n289 ;
  assign n361 = n116 & n360 ;
  assign n362 = n280 & n361 ;
  assign n363 = n79 & n362 ;
  assign n364 = G13 | n363 ;
  assign n365 = G13 & n363 ;
  assign n366 = n364 & ~n365 ;
  assign n367 = n272 & n362 ;
  assign n368 = ~G14 & n367 ;
  assign n369 = G14 & ~n367 ;
  assign n370 = n368 | n369 ;
  assign n371 = n222 & n362 ;
  assign n372 = G15 | n371 ;
  assign n373 = G15 & n371 ;
  assign n374 = n372 & ~n373 ;
  assign n375 = n250 & n362 ;
  assign n376 = ~G16 & n375 ;
  assign n377 = G16 & ~n375 ;
  assign n378 = n376 | n377 ;
  assign n379 = n192 & n330 ;
  assign n380 = G17 | n379 ;
  assign n381 = G17 & n330 ;
  assign n382 = n192 & n381 ;
  assign n383 = n380 & ~n382 ;
  assign n384 = n116 & n330 ;
  assign n385 = G18 & n384 ;
  assign n386 = G18 | n384 ;
  assign n387 = ~n385 & n386 ;
  assign n388 = n173 & n330 ;
  assign n389 = G19 | n388 ;
  assign n390 = G19 & n330 ;
  assign n391 = n173 & n390 ;
  assign n392 = n389 & ~n391 ;
  assign n393 = n116 & n295 ;
  assign n394 = G22 & n393 ;
  assign n395 = G22 | n393 ;
  assign n396 = ~n394 & n395 ;
  assign n397 = n173 & n295 ;
  assign n398 = G23 | n397 ;
  assign n399 = G23 & n295 ;
  assign n400 = n173 & n399 ;
  assign n401 = n398 & ~n400 ;
  assign n402 = n144 & n295 ;
  assign n403 = G24 | n402 ;
  assign n404 = G24 & n295 ;
  assign n405 = n144 & n404 ;
  assign n406 = n403 & ~n405 ;
  assign n407 = n251 & n293 ;
  assign n408 = n276 & n407 ;
  assign n409 = n192 & n408 ;
  assign n410 = G25 | n409 ;
  assign n411 = G25 & n408 ;
  assign n412 = n192 & n411 ;
  assign n413 = n410 & ~n412 ;
  assign n414 = n116 & n408 ;
  assign n415 = G26 & n414 ;
  assign n416 = G26 | n414 ;
  assign n417 = ~n415 & n416 ;
  assign n418 = n173 & n408 ;
  assign n419 = G27 | n418 ;
  assign n420 = G27 & n408 ;
  assign n421 = n173 & n420 ;
  assign n422 = n419 & ~n421 ;
  assign n423 = n144 & n408 ;
  assign n424 = G28 | n423 ;
  assign n425 = G28 & n408 ;
  assign n426 = n144 & n425 ;
  assign n427 = n424 & ~n426 ;
  assign n428 = n250 & n293 ;
  assign n429 = n78 | n221 ;
  assign n430 = n77 | n220 ;
  assign n431 = n429 | n430 ;
  assign n432 = n272 & ~n431 ;
  assign n433 = n428 & n432 ;
  assign n434 = n192 & n433 ;
  assign n435 = G29 | n434 ;
  assign n436 = G29 & n433 ;
  assign n437 = n192 & n436 ;
  assign n438 = n435 & ~n437 ;
  assign n439 = n116 & n433 ;
  assign n440 = G30 & n439 ;
  assign n441 = G30 | n439 ;
  assign n442 = ~n440 & n441 ;
  assign n443 = n173 & n433 ;
  assign n444 = G31 | n443 ;
  assign n445 = G31 & n433 ;
  assign n446 = n173 & n445 ;
  assign n447 = n444 & ~n446 ;
  assign n448 = n144 & n433 ;
  assign n449 = G32 | n448 ;
  assign n450 = G32 & n433 ;
  assign n451 = n144 & n450 ;
  assign n452 = n449 & ~n451 ;
  assign G1324 = ~n286 ;
  assign G1344 = ~n300 ;
  assign G1325 = ~n304 ;
  assign G1326 = ~n308 ;
  assign G1327 = ~n312 ;
  assign G1328 = ~n321 ;
  assign G1329 = ~n325 ;
  assign G1330 = ~n329 ;
  assign G1343 = ~n335 ;
  assign G1331 = ~n339 ;
  assign G1332 = ~n347 ;
  assign G1333 = ~n351 ;
  assign G1334 = ~n355 ;
  assign G1335 = ~n359 ;
  assign G1336 = ~n366 ;
  assign G1337 = ~n370 ;
  assign G1338 = ~n374 ;
  assign G1339 = ~n378 ;
  assign G1340 = ~n383 ;
  assign G1341 = ~n387 ;
  assign G1342 = ~n392 ;
  assign G1345 = ~n396 ;
  assign G1346 = ~n401 ;
  assign G1347 = ~n406 ;
  assign G1348 = ~n413 ;
  assign G1349 = ~n417 ;
  assign G1350 = ~n422 ;
  assign G1351 = ~n427 ;
  assign G1352 = ~n438 ;
  assign G1353 = ~n442 ;
  assign G1354 = ~n447 ;
  assign G1355 = ~n452 ;
endmodule
