/****************************************************************************
 *                                                                          *
 *  VERILOG VERSION of ORIGINAL NETLIST for c1908                           *
 *                                                                          *  
 *                                                                          *
 *  Generated by: Hakan Yalcin (hyalcin@cadence.com)                        *
 *                                                                          *
 *                Sep 16, 1998                                              *
 *                                                                          *
****************************************************************************/
module c1908g (
        L101, L104, L107, L110, L113, L116, L119,
        L122, L125, L128, L131, L134, L137, L140, L143,
        L146, L210, L214, L217, L221, L224, L227, L234,
        L237, L469, L472, L475, L478, L898, L900, L902,
        L952, L953,
        L3, L6, L9, L12, L30, L45, L48,
        L15, L18, L21, L24, L27, L33, L36, L39,
        L42, L75, L51, L54, L60, L63, L66, L69,
        L72, L57);
 
   input
        L101, L104, L107, L110, L113, L116, L119,
        L122, L125, L128, L131, L134, L137, L140, L143,
        L146, L210, L214, L217, L221, L224, L227, L234,
        L237, L469, L472, L475, L478, L898, L900, L902,
        L952, L953;
 
   output
        L3, L6, L9, L12, L30, L45, L48,
        L15, L18, L21, L24, L27, L33, L36, L39,
        L42, L75, L51, L54, L60, L63, L66, L69,
        L72, L57;


   inv U1 ( L101, L149 ); 
   inv U2 ( L104, L153 ); 
   inv U3 ( L107, L156 ); 
   inv U4 ( L110, L160 ); 
   inv U5 ( L113, L165 ); 
   inv U6 ( L116, L168 ); 
   inv U7 ( L119, L171 ); 
   inv U8 ( L122, L175 ); 
   inv U9 ( L125, L179 ); 
   inv U10 ( L128, L184 ); 
   inv U11 ( L131, L188 ); 
   inv U12 ( L134, L191 ); 
   inv U13 ( L137, L194 ); 
   inv U14 ( L140, L198 ); 
   inv U15 ( L143, L202 ); 
   inv U16 ( L146, L206 ); 
   nand2 U17 ( L224, L898, L231 ); 
   nand2 U18 ( L227, L900, L233 ); 
   inv U19 ( L237, L241 ); 
   inv U20 ( L237, L244 ); 
   buffer U21 ( L234, L245 ); 
   buffer U22 ( L234, L248 ); 
   inv U23 ( L469, L517 ); 
   inv U24 ( L472, L529 ); 
   inv U25 ( L475, L541 ); 
   inv U26 ( L478, L553 ); 
   inv U27 ( L953, L859 ); 
   inv U28 ( L953, L862 ); 
   inv U29 ( L898, L907 ); 
   inv U30 ( L900, L909 ); 
   buffer U31 ( L902, L911 ); 
   inv U32 ( L902, L918 ); 
   buffer U33 ( L902, L919 ); 
   inv U34 ( L902, L922 ); 
   buffer U35 ( L952, L926 ); 
   inv U36 ( L952, L930 ); 
   inv U37 ( L952, L932 ); 
   buffer U38 ( L953, L934 ); 
   inv U39 ( L953, L938 ); 
   buffer U40 ( L953, L943 ); 
   buffer U41 ( L953, L947 ); 
   inv U42 ( L953, L949 ); 
   buffer U43 ( L101, L1506 ); 
   buffer U44 ( L104, L1514 ); 
   buffer U45 ( L107, L1522 ); 
   buffer U46 ( L110, L1530 ); 
   buffer U47 ( L113, L1538 ); 
   buffer U48 ( L116, L1546 ); 
   buffer U49 ( L119, L1554 ); 
   buffer U50 ( L122, L1562 ); 
   buffer U51 ( L125, L1570 ); 
   buffer U52 ( L128, L1578 ); 
   buffer U53 ( L131, L1586 ); 
   buffer U54 ( L134, L1594 ); 
   buffer U55 ( L137, L1602 ); 
   buffer U56 ( L140, L1610 ); 
   buffer U57 ( L143, L1618 ); 
   buffer U58 ( L146, L1626 ); 
   inv U59 ( L1506, L1512 ); 
   inv U60 ( L1514, L1520 ); 
   inv U61 ( L1522, L1528 ); 
   inv U62 ( L1530, L1536 ); 
   inv U63 ( L1538, L1544 ); 
   inv U64 ( L1546, L1552 ); 
   inv U65 ( L1554, L1560 ); 
   inv U66 ( L1562, L1568 ); 
   inv U67 ( L1570, L1576 ); 
   inv U68 ( L1578, L1584 ); 
   inv U69 ( L1586, L1592 ); 
   inv U70 ( L1594, L1600 ); 
   inv U71 ( L1602, L1608 ); 
   inv U72 ( L1610, L1616 ); 
   inv U73 ( L1618, L1624 ); 
   inv U74 ( L1626, L1632 ); 
   nand2 U75 ( L930, L947, L50 ); 
   nand2 U76 ( L930, L947, L52 ); 
   nand2 U77 ( L930, L947, L56 ); 
   nand2 U78 ( L930, L947, L58 ); 
   nand2 U79 ( L930, L947, L62 ); 
   nand2 U80 ( L930, L947, L64 ); 
   buffer U81 ( L149, L251 ); 
   buffer U82 ( L153, L254 ); 
   buffer U83 ( L165, L288 ); 
   buffer U84 ( L168, L291 ); 
   buffer U85 ( L184, L299 ); 
   buffer U86 ( L202, L302 ); 
   and2 U87 ( L224, L938, L318 ); 
   buffer U88 ( L179, L321 ); 
   buffer U89 ( L188, L327 ); 
   buffer U90 ( L191, L330 ); 
   and2 U91 ( L227, L938, L352 ); 
   buffer U92 ( L198, L355 ); 
   and3 U93 ( L210, L241, L938, L369 ); 
   buffer U94 ( L206, L382 ); 
   buffer U95 ( L198, L385 ); 
   nand2 U96 ( L943, L907, L853 ); 
   nand2 U97 ( L943, L909, L856 ); 
   nand2 U98 ( L248, L237, L893 ); 
   nand2 U99 ( L248, L922, L954 ); 
   nand2 U100 ( L244, L922, L955 ); 
   buffer U101 ( L160, L1050 ); 
   buffer U102 ( L175, L1053 ); 
   buffer U103 ( L179, L1176 ); 
   buffer U104 ( L198, L1179 ); 
   buffer U105 ( L149, L1197 ); 
   buffer U106 ( L149, L1207 ); 
   buffer U107 ( L153, L1222 ); 
   buffer U108 ( L188, L1244 ); 
   buffer U109 ( L156, L1278 ); 
   and3 U110 ( L217, L245, L938, L1290 ); 
   buffer U111 ( L191, L1300 ); 
   buffer U112 ( L160, L1312 ); 
   buffer U113 ( L194, L1332 ); 
   and3 U114 ( L221, L245, L938, L1335 ); 
   buffer U115 ( L517, L1442 ); 
   buffer U116 ( L517, L1450 ); 
   buffer U117 ( L529, L1458 ); 
   buffer U118 ( L529, L1466 ); 
   buffer U119 ( L541, L1474 ); 
   buffer U120 ( L541, L1482 ); 
   buffer U121 ( L553, L1490 ); 
   buffer U122 ( L553, L1498 ); 
   and2 U123 ( L231, L934, L1634 ); 
   and2 U124 ( L233, L934, L1644 ); 
   buffer U125 ( L156, L1657 ); 
   buffer U126 ( L156, L1665 ); 
   buffer U127 ( L171, L1697 ); 
   buffer U128 ( L171, L1705 ); 
   buffer U129 ( L206, L1713 ); 
   buffer U130 ( L206, L1721 ); 
   buffer U131 ( L194, L1745 ); 
   buffer U132 ( L194, L1753 ); 
   buffer U133 ( L160, L1785 ); 
   buffer U134 ( L160, L1793 ); 
   buffer U135 ( L165, L1814 ); 
   buffer U136 ( L175, L1817 ); 
   and3 U137 ( L214, L241, L938, L1830 ); 
   buffer U138 ( L202, L1833 ); 
   buffer U139 ( L179, L1841 ); 
   buffer U140 ( L179, L1849 ); 
   buffer U141 ( L168, L1854 ); 
   buffer U142 ( L175, L1857 ); 
   buffer U143 ( L184, L1870 ); 
   buffer U144 ( L202, L1873 ); 
   buffer U145 ( L171, L1878 ); 
   buffer U146 ( L184, L1881 ); 
   inv U147 ( L1634, L1642 ); 
   inv U148 ( L1644, L1652 ); 
   inv U149 ( L1050, L1056 ); 
   inv U150 ( L1053, L1057 ); 
   inv U151 ( L1176, L1182 ); 
   inv U152 ( L1179, L1183 ); 
   inv U153 ( L1207, L1211 ); 
   inv U154 ( L1290, L1298 ); 
   inv U155 ( L1312, L1320 ); 
   inv U156 ( L1332, L1338 ); 
   inv U157 ( L1335, L1339 ); 
   and2 U158 ( L210, L955, L457 ); 
   and2 U159 ( L217, L954, L459 ); 
   nand2 U160 ( L214, L955, L482 ); 
   nand2 U161 ( L221, L954, L487 ); 
   nand2 U162 ( L210, L955, L492 ); 
   nand2 U163 ( L217, L954, L505 ); 
   inv U164 ( L1450, L1456 ); 
   inv U165 ( L1442, L1448 ); 
   inv U166 ( L1466, L1472 ); 
   inv U167 ( L1458, L1464 ); 
   inv U168 ( L1482, L1488 ); 
   inv U169 ( L1474, L1480 ); 
   inv U170 ( L1498, L1504 ); 
   inv U171 ( L1490, L1496 ); 
   nand4 U172 ( L907, L919, L943, L893, L956 ); 
   nand4 U173 ( L909, L919, L943, L893, L967 ); 
   nand3 U174 ( L926, L949, L893, L978 ); 
   and3 U175 ( L926, L949, L893, L979 ); 
   buffer U176 ( L251, L980 ); 
   inv U177 ( L1657, L1661 ); 
   buffer U178 ( L251, L990 ); 
   inv U179 ( L1665, L1669 ); 
   buffer U180 ( L288, L1030 ); 
   inv U181 ( L1697, L1701 ); 
   buffer U182 ( L288, L1040 ); 
   inv U183 ( L1705, L1709 ); 
   buffer U184 ( L299, L1058 ); 
   inv U185 ( L1713, L1717 ); 
   buffer U186 ( L299, L1068 ); 
   inv U187 ( L1721, L1725 ); 
   buffer U188 ( L318, L1078 ); 
   buffer U189 ( L318, L1090 ); 
   buffer U190 ( L327, L1100 ); 
   inv U191 ( L1745, L1749 ); 
   buffer U192 ( L327, L1112 ); 
   inv U193 ( L1753, L1757 ); 
   buffer U194 ( L352, L1154 ); 
   inv U195 ( L1785, L1789 ); 
   buffer U196 ( L352, L1166 ); 
   inv U197 ( L1793, L1797 ); 
   buffer U198 ( L369, L1194 ); 
   inv U199 ( L1197, L1201 ); 
   buffer U200 ( L369, L1204 ); 
   inv U201 ( L1814, L1820 ); 
   inv U202 ( L1817, L1821 ); 
   inv U203 ( L1222, L1230 ); 
   inv U204 ( L1830, L1836 ); 
   inv U205 ( L1833, L1837 ); 
   inv U206 ( L1244, L1252 ); 
   buffer U207 ( L382, L1256 ); 
   inv U208 ( L1841, L1845 ); 
   buffer U209 ( L382, L1268 ); 
   inv U210 ( L1849, L1853 ); 
   inv U211 ( L1854, L1860 ); 
   inv U212 ( L1857, L1861 ); 
   inv U213 ( L1278, L1286 ); 
   inv U214 ( L1870, L1876 ); 
   inv U215 ( L1873, L1877 ); 
   inv U216 ( L1300, L1308 ); 
   inv U217 ( L1878, L1884 ); 
   inv U218 ( L1881, L1885 ); 
   buffer U219 ( L254, L1654 ); 
   buffer U220 ( L254, L1662 ); 
   buffer U221 ( L291, L1694 ); 
   buffer U222 ( L291, L1702 ); 
   buffer U223 ( L302, L1710 ); 
   buffer U224 ( L302, L1718 ); 
   buffer U225 ( L321, L1726 ); 
   buffer U226 ( L321, L1734 ); 
   buffer U227 ( L330, L1742 ); 
   buffer U228 ( L330, L1750 ); 
   buffer U229 ( L355, L1782 ); 
   buffer U230 ( L355, L1790 ); 
   buffer U231 ( L385, L1838 ); 
   buffer U232 ( L385, L1846 ); 
   nand2 U233 ( L1053, L1056, L297 ); 
   nand2 U234 ( L1050, L1057, L298 ); 
   nand2 U235 ( L1179, L1182, L361 ); 
   nand2 U236 ( L1176, L1183, L362 ); 
   nand2 U237 ( L1335, L1338, L404 ); 
   nand2 U238 ( L1332, L1339, L405 ); 
   nand2 U239 ( L1817, L1820, L1225 ); 
   nand2 U240 ( L1814, L1821, L1226 ); 
   nand2 U241 ( L1833, L1836, L1247 ); 
   nand2 U242 ( L1830, L1837, L1248 ); 
   nand2 U243 ( L1857, L1860, L1281 ); 
   nand2 U244 ( L1854, L1861, L1282 ); 
   nand2 U245 ( L1873, L1876, L1303 ); 
   nand2 U246 ( L1870, L1877, L1304 ); 
   nand2 U247 ( L1881, L1884, L1315 ); 
   nand2 U248 ( L1878, L1885, L1316 ); 
   inv U249 ( L990, L998 ); 
   inv U250 ( L980, L988 ); 
   nand2 U251 ( L297, L298, L268 ); 
   inv U252 ( L1030, L1038 ); 
   inv U253 ( L1040, L1048 ); 
   inv U254 ( L1068, L1076 ); 
   inv U255 ( L1058, L1066 ); 
   inv U256 ( L1090, L1098 ); 
   inv U257 ( L1112, L1120 ); 
   inv U258 ( L1166, L1174 ); 
   nand2 U259 ( L361, L362, L363 ); 
   inv U260 ( L1204, L1210 ); 
   nand2 U261 ( L1204, L1211, L373 ); 
   inv U262 ( L1268, L1276 ); 
   nand2 U263 ( L404, L405, L406 ); 
   inv U264 ( L482, L565 ); 
   buffer U265 ( L482, L566 ); 
   inv U266 ( L487, L614 ); 
   buffer U267 ( L487, L615 ); 
   nand2 U268 ( L956, L978, L958 ); 
   nand2 U269 ( L967, L978, L969 ); 
   inv U270 ( L1654, L1660 ); 
   nand2 U271 ( L1654, L1661, L984 ); 
   inv U272 ( L1662, L1668 ); 
   nand2 U273 ( L1662, L1669, L994 ); 
   inv U274 ( L1694, L1700 ); 
   nand2 U275 ( L1694, L1701, L1034 ); 
   inv U276 ( L1702, L1708 ); 
   nand2 U277 ( L1702, L1709, L1044 ); 
   inv U278 ( L1710, L1716 ); 
   nand2 U279 ( L1710, L1717, L1062 ); 
   inv U280 ( L1718, L1724 ); 
   nand2 U281 ( L1718, L1725, L1072 ); 
   inv U282 ( L1726, L1732 ); 
   inv U283 ( L1078, L1086 ); 
   inv U284 ( L1734, L1740 ); 
   inv U285 ( L1742, L1748 ); 
   nand2 U286 ( L1742, L1749, L1104 ); 
   inv U287 ( L1100, L1108 ); 
   inv U288 ( L1750, L1756 ); 
   nand2 U289 ( L1750, L1757, L1116 ); 
   inv U290 ( L1782, L1788 ); 
   nand2 U291 ( L1782, L1789, L1158 ); 
   inv U292 ( L1154, L1162 ); 
   inv U293 ( L1790, L1796 ); 
   nand2 U294 ( L1790, L1797, L1170 ); 
   inv U295 ( L1194, L1200 ); 
   nand2 U296 ( L1194, L1201, L1203 ); 
   nand2 U297 ( L1225, L1226, L1227 ); 
   nand2 U298 ( L1247, L1248, L1249 ); 
   inv U299 ( L1838, L1844 ); 
   nand2 U300 ( L1838, L1845, L1260 ); 
   inv U301 ( L1256, L1264 ); 
   inv U302 ( L1846, L1852 ); 
   nand2 U303 ( L1846, L1853, L1272 ); 
   nand2 U304 ( L1281, L1282, L1283 ); 
   nand2 U305 ( L1303, L1304, L1305 ); 
   nand2 U306 ( L1315, L1316, L1317 ); 
   buffer U307 ( L492, L1410 ); 
   buffer U308 ( L492, L1418 ); 
   buffer U309 ( L505, L1426 ); 
   buffer U310 ( L505, L1434 ); 
   inv U311 ( L268, L269 ); 
   nand2 U312 ( L1207, L1210, L372 ); 
   nand2 U313 ( L1657, L1660, L983 ); 
   nand2 U314 ( L1665, L1668, L993 ); 
   nand2 U315 ( L1697, L1700, L1033 ); 
   nand2 U316 ( L1705, L1708, L1043 ); 
   nand2 U317 ( L1713, L1716, L1061 ); 
   nand2 U318 ( L1721, L1724, L1071 ); 
   nand2 U319 ( L1745, L1748, L1103 ); 
   nand2 U320 ( L1753, L1756, L1115 ); 
   nand2 U321 ( L1785, L1788, L1157 ); 
   nand2 U322 ( L1793, L1796, L1169 ); 
   inv U323 ( L363, L1184 ); 
   nand2 U324 ( L1197, L1200, L1202 ); 
   nand2 U325 ( L1841, L1844, L1259 ); 
   nand2 U326 ( L1849, L1852, L1271 ); 
   inv U327 ( L406, L1322 ); 
   nand2 U328 ( L372, L373, L374 ); 
   nand2 U329 ( L1317, L1320, L396 ); 
   inv U330 ( L1317, L1321 ); 
   inv U331 ( L1418, L1424 ); 
   inv U332 ( L1410, L1416 ); 
   inv U333 ( L1434, L1440 ); 
   inv U334 ( L1426, L1432 ); 
   nand2 U335 ( L983, L984, L985 ); 
   nand2 U336 ( L993, L994, L995 ); 
   nand2 U337 ( L1033, L1034, L1035 ); 
   nand2 U338 ( L1043, L1044, L1045 ); 
   nand2 U339 ( L1061, L1062, L1063 ); 
   nand2 U340 ( L1071, L1072, L1073 ); 
   nand2 U341 ( L1103, L1104, L1105 ); 
   nand2 U342 ( L1115, L1116, L1117 ); 
   nand2 U343 ( L1157, L1158, L1159 ); 
   nand2 U344 ( L1169, L1170, L1171 ); 
   nand2 U345 ( L1202, L1203, L1212 ); 
   inv U346 ( L1227, L1231 ); 
   nand2 U347 ( L1227, L1230, L1232 ); 
   inv U348 ( L1249, L1253 ); 
   nand2 U349 ( L1249, L1252, L1254 ); 
   nand2 U350 ( L1259, L1260, L1261 ); 
   nand2 U351 ( L1271, L1272, L1273 ); 
   inv U352 ( L1283, L1287 ); 
   nand2 U353 ( L1283, L1286, L1288 ); 
   inv U354 ( L1305, L1309 ); 
   nand2 U355 ( L1305, L1308, L1310 ); 
   inv U356 ( L1184, L1192 ); 
   nand2 U357 ( L1312, L1321, L397 ); 
   inv U358 ( L1322, L1330 ); 
   buffer U359 ( L269, L1000 ); 
   buffer U360 ( L269, L1010 ); 
   nand2 U361 ( L1222, L1231, L1233 ); 
   nand2 U362 ( L1244, L1253, L1255 ); 
   nand2 U363 ( L1278, L1287, L1289 ); 
   nand2 U364 ( L1300, L1309, L1311 ); 
   inv U365 ( L374, L1381 ); 
   nand2 U366 ( L995, L998, L257 ); 
   inv U367 ( L995, L999 ); 
   nand2 U368 ( L985, L988, L260 ); 
   inv U369 ( L985, L989 ); 
   nand2 U370 ( L1035, L1038, L272 ); 
   inv U371 ( L1035, L1039 ); 
   nand2 U372 ( L1045, L1048, L294 ); 
   inv U373 ( L1045, L1049 ); 
   nand2 U374 ( L1073, L1076, L305 ); 
   inv U375 ( L1073, L1077 ); 
   nand2 U376 ( L1063, L1066, L308 ); 
   inv U377 ( L1063, L1067 ); 
   nand2 U378 ( L1117, L1120, L333 ); 
   inv U379 ( L1117, L1121 ); 
   nand2 U380 ( L1171, L1174, L358 ); 
   inv U381 ( L1171, L1175 ); 
   inv U382 ( L1212, L1220 ); 
   nand2 U383 ( L1273, L1276, L388 ); 
   inv U384 ( L1273, L1277 ); 
   nand2 U385 ( L396, L397, L398 ); 
   inv U386 ( L1105, L1109 ); 
   nand2 U387 ( L1105, L1108, L1110 ); 
   inv U388 ( L1159, L1163 ); 
   nand2 U389 ( L1159, L1162, L1164 ); 
   nand2 U390 ( L1232, L1233, L1234 ); 
   inv U391 ( L1261, L1265 ); 
   nand2 U392 ( L1261, L1264, L1266 ); 
   nand2 U393 ( L1254, L1255, L1822 ); 
   nand2 U394 ( L1310, L1311, L1862 ); 
   nand2 U395 ( L1288, L1289, L1865 ); 
   nand2 U396 ( L990, L999, L258 ); 
   nand2 U397 ( L980, L989, L261 ); 
   nand2 U398 ( L1030, L1039, L273 ); 
   inv U399 ( L1010, L1018 ); 
   inv U400 ( L1000, L1008 ); 
   nand2 U401 ( L1040, L1049, L295 ); 
   nand2 U402 ( L1068, L1077, L306 ); 
   nand2 U403 ( L1058, L1067, L309 ); 
   nand2 U404 ( L1112, L1121, L334 ); 
   nand2 U405 ( L1166, L1175, L359 ); 
   nand2 U406 ( L1268, L1277, L389 ); 
   inv U407 ( L1381, L1385 ); 
   nand2 U408 ( L1100, L1109, L1111 ); 
   nand2 U409 ( L1154, L1163, L1165 ); 
   nand2 U410 ( L1256, L1265, L1267 ); 
   inv U411 ( L398, L1886 ); 
   nand2 U412 ( L257, L258, L259 ); 
   nand2 U413 ( L260, L261, L262 ); 
   nand2 U414 ( L272, L273, L274 ); 
   nand2 U415 ( L294, L295, L296 ); 
   nand2 U416 ( L305, L306, L307 ); 
   nand2 U417 ( L308, L309, L310 ); 
   nand2 U418 ( L333, L334, L335 ); 
   nand2 U419 ( L358, L359, L360 ); 
   inv U420 ( L1234, L1242 ); 
   nand2 U421 ( L388, L389, L390 ); 
   inv U422 ( L1822, L1828 ); 
   inv U423 ( L1862, L1868 ); 
   inv U424 ( L1865, L1869 ); 
   nand2 U425 ( L1164, L1165, L1373 ); 
   nand2 U426 ( L1110, L1111, L1798 ); 
   nand2 U427 ( L1266, L1267, L1825 ); 
   inv U428 ( L259, L265 ); 
   inv U429 ( L307, L314 ); 
   inv U430 ( L335, L336 ); 
   inv U431 ( L296, L407 ); 
   nand2 U432 ( L1865, L1868, L1293 ); 
   nand2 U433 ( L1862, L1869, L1294 ); 
   inv U434 ( L1886, L1892 ); 
   inv U435 ( L360, L1777 ); 
   inv U436 ( L390, L1889 ); 
   buffer U437 ( L310, L410 ); 
   inv U438 ( L1373, L1377 ); 
   inv U439 ( L1798, L1804 ); 
   nand2 U440 ( L1825, L1828, L1237 ); 
   inv U441 ( L1825, L1829 ); 
   nand2 U442 ( L1293, L1294, L1295 ); 
   buffer U443 ( L274, L1670 ); 
   buffer U444 ( L274, L1678 ); 
   buffer U445 ( L310, L1729 ); 
   buffer U446 ( L310, L1737 ); 
   buffer U447 ( L262, L1761 ); 
   buffer U448 ( L262, L1769 ); 
   buffer U449 ( L336, L340 ); 
   buffer U450 ( L314, L343 ); 
   inv U451 ( L1777, L1781 ); 
   nand2 U452 ( L1822, L1829, L1238 ); 
   nand2 U453 ( L1889, L1892, L1325 ); 
   inv U454 ( L1889, L1893 ); 
   buffer U455 ( L407, L1340 ); 
   buffer U456 ( L407, L1352 ); 
   buffer U457 ( L265, L1673 ); 
   buffer U458 ( L265, L1681 ); 
   buffer U459 ( L314, L1801 ); 
   buffer U460 ( L336, L1897 ); 
   buffer U461 ( L336, L1905 ); 
   nand2 U462 ( L1295, L1298, L391 ); 
   inv U463 ( L1295, L1299 ); 
   inv U464 ( L1670, L1676 ); 
   inv U465 ( L1678, L1684 ); 
   nand2 U466 ( L1729, L1732, L1081 ); 
   inv U467 ( L1729, L1733 ); 
   nand2 U468 ( L1737, L1740, L1093 ); 
   inv U469 ( L1737, L1741 ); 
   inv U470 ( L1761, L1765 ); 
   inv U471 ( L1769, L1773 ); 
   nand2 U472 ( L1237, L1238, L1239 ); 
   nand2 U473 ( L1886, L1893, L1326 ); 
   buffer U474 ( L410, L1894 ); 
   buffer U475 ( L410, L1902 ); 
   nand2 U476 ( L1290, L1299, L392 ); 
   inv U477 ( L1352, L1360 ); 
   nand2 U478 ( L1673, L1676, L1003 ); 
   inv U479 ( L1673, L1677 ); 
   nand2 U480 ( L1681, L1684, L1013 ); 
   inv U481 ( L1681, L1685 ); 
   nand2 U482 ( L1726, L1733, L1082 ); 
   nand2 U483 ( L1734, L1741, L1094 ); 
   buffer U484 ( L340, L1122 ); 
   buffer U485 ( L340, L1134 ); 
   nand2 U486 ( L1801, L1804, L1187 ); 
   inv U487 ( L1801, L1805 ); 
   nand2 U488 ( L1325, L1326, L1327 ); 
   inv U489 ( L1897, L1901 ); 
   inv U490 ( L1340, L1348 ); 
   inv U491 ( L1905, L1909 ); 
   buffer U492 ( L343, L1758 ); 
   buffer U493 ( L343, L1766 ); 
   nand2 U494 ( L1239, L1242, L377 ); 
   inv U495 ( L1239, L1243 ); 
   nand2 U496 ( L391, L392, L393 ); 
   nand2 U497 ( L1670, L1677, L1004 ); 
   nand2 U498 ( L1678, L1685, L1014 ); 
   nand2 U499 ( L1081, L1082, L1083 ); 
   nand2 U500 ( L1093, L1094, L1095 ); 
   nand2 U501 ( L1798, L1805, L1188 ); 
   inv U502 ( L1894, L1900 ); 
   nand2 U503 ( L1894, L1901, L1344 ); 
   inv U504 ( L1902, L1908 ); 
   nand2 U505 ( L1902, L1909, L1356 ); 
   inv U506 ( L1134, L1142 ); 
   nand2 U507 ( L1234, L1243, L378 ); 
   nand2 U508 ( L1327, L1330, L399 ); 
   inv U509 ( L1327, L1331 ); 
   nand2 U510 ( L1003, L1004, L1005 ); 
   nand2 U511 ( L1013, L1014, L1015 ); 
   inv U512 ( L1758, L1764 ); 
   nand2 U513 ( L1758, L1765, L1126 ); 
   inv U514 ( L1122, L1130 ); 
   inv U515 ( L1766, L1772 ); 
   nand2 U516 ( L1766, L1773, L1138 ); 
   nand2 U517 ( L1187, L1188, L1189 ); 
   nand2 U518 ( L1897, L1900, L1343 ); 
   nand2 U519 ( L1905, L1908, L1355 ); 
   nand2 U520 ( L1095, L1098, L324 ); 
   inv U521 ( L1095, L1099 ); 
   nand2 U522 ( L377, L378, L379 ); 
   nand2 U523 ( L1322, L1331, L400 ); 
   nand2 U524 ( L393, L918, L449 ); 
   inv U525 ( L1083, L1087 ); 
   nand2 U526 ( L1083, L1086, L1088 ); 
   nand2 U527 ( L1761, L1764, L1125 ); 
   nand2 U528 ( L1769, L1772, L1137 ); 
   nand2 U529 ( L1343, L1344, L1345 ); 
   nand2 U530 ( L1355, L1356, L1357 ); 
   buffer U531 ( L393, L1397 ); 
   nand2 U532 ( L1015, L1018, L277 ); 
   inv U533 ( L1015, L1019 ); 
   nand2 U534 ( L1005, L1008, L280 ); 
   inv U535 ( L1005, L1009 ); 
   nand2 U536 ( L1090, L1099, L325 ); 
   nand2 U537 ( L1189, L1192, L364 ); 
   inv U538 ( L1189, L1193 ); 
   nand2 U539 ( L399, L400, L401 ); 
   nand2 U540 ( L1078, L1087, L1089 ); 
   nand2 U541 ( L1125, L1126, L1127 ); 
   nand2 U542 ( L1137, L1138, L1139 ); 
   nand2 U543 ( L1010, L1019, L278 ); 
   nand2 U544 ( L1000, L1009, L281 ); 
   nand2 U545 ( L324, L325, L326 ); 
   nand2 U546 ( L1184, L1193, L365 ); 
   nand2 U547 ( L1357, L1360, L413 ); 
   inv U548 ( L1357, L1361 ); 
   inv U549 ( L1397, L1401 ); 
   nand2 U550 ( L379, L918, L445 ); 
   inv U551 ( L1345, L1349 ); 
   nand2 U552 ( L1345, L1348, L1350 ); 
   buffer U553 ( L379, L1389 ); 
   buffer U554 ( L449, L1493 ); 
   buffer U555 ( L449, L1501 ); 
   nand2 U556 ( L1088, L1089, L1689 ); 
   nand2 U557 ( L277, L278, L279 ); 
   nand2 U558 ( L280, L281, L282 ); 
   nand2 U559 ( L1139, L1142, L346 ); 
   inv U560 ( L1139, L1143 ); 
   nand2 U561 ( L364, L365, L366 ); 
   nand2 U562 ( L1352, L1361, L414 ); 
   nand2 U563 ( L401, L918, L453 ); 
   inv U564 ( L1127, L1131 ); 
   nand2 U565 ( L1127, L1130, L1132 ); 
   nand2 U566 ( L1340, L1349, L1351 ); 
   inv U567 ( L326, L1365 ); 
   buffer U568 ( L401, L1405 ); 
   inv U569 ( L279, L285 ); 
   nand2 U570 ( L1134, L1143, L347 ); 
   inv U571 ( L366, L367 ); 
   nand2 U572 ( L413, L414, L415 ); 
   inv U573 ( L1389, L1393 ); 
   nand2 U574 ( L1501, L1504, L556 ); 
   inv U575 ( L1501, L1505 ); 
   nand2 U576 ( L1493, L1496, L559 ); 
   inv U577 ( L1493, L1497 ); 
   inv U578 ( L1689, L1693 ); 
   nand2 U579 ( L1122, L1131, L1133 ); 
   buffer U580 ( L445, L1477 ); 
   buffer U581 ( L445, L1485 ); 
   nand2 U582 ( L1350, L1351, L1809 ); 
   nand2 U583 ( L346, L347, L348 ); 
   inv U584 ( L1365, L1369 ); 
   inv U585 ( L1405, L1409 ); 
   nand2 U586 ( L1498, L1505, L557 ); 
   nand2 U587 ( L1490, L1497, L560 ); 
   buffer U588 ( L282, L1362 ); 
   inv U589 ( L415, L1378 ); 
   buffer U590 ( L453, L1429 ); 
   buffer U591 ( L453, L1437 ); 
   buffer U592 ( L282, L1686 ); 
   nand2 U593 ( L1132, L1133, L1774 ); 
   and2 U594 ( L285, L853, L1910 ); 
   and2 U595 ( L856, L367, L1918 ); 
   nand2 U596 ( L1485, L1488, L544 ); 
   inv U597 ( L1485, L1489 ); 
   nand2 U598 ( L1477, L1480, L547 ); 
   inv U599 ( L1477, L1481 ); 
   nand2 U600 ( L556, L557, L558 ); 
   nand2 U601 ( L559, L560, L561 ); 
   inv U602 ( L1809, L1813 ); 
   inv U603 ( L348, L1370 ); 
   inv U604 ( L1362, L1368 ); 
   nand2 U605 ( L1362, L1369, L417 ); 
   inv U606 ( L1378, L1384 ); 
   nand2 U607 ( L1378, L1385, L424 ); 
   nand2 U608 ( L1437, L1440, L508 ); 
   inv U609 ( L1437, L1441 ); 
   nand2 U610 ( L1429, L1432, L511 ); 
   inv U611 ( L1429, L1433 ); 
   nand2 U612 ( L1482, L1489, L545 ); 
   nand2 U613 ( L1474, L1481, L548 ); 
   inv U614 ( L558, L564 ); 
   inv U615 ( L1686, L1692 ); 
   nand2 U616 ( L1686, L1693, L1024 ); 
   inv U617 ( L1774, L1780 ); 
   nand2 U618 ( L1774, L1781, L1148 ); 
   inv U619 ( L1910, L1916 ); 
   inv U620 ( L1918, L1924 ); 
   nand2 U621 ( L1365, L1368, L416 ); 
   inv U622 ( L1370, L1376 ); 
   nand2 U623 ( L1370, L1377, L421 ); 
   nand2 U624 ( L1381, L1384, L423 ); 
   nand2 U625 ( L1434, L1441, L509 ); 
   nand2 U626 ( L1426, L1433, L512 ); 
   nand2 U627 ( L544, L545, L546 ); 
   nand2 U628 ( L547, L548, L549 ); 
   inv U629 ( L561, L719 ); 
   buffer U630 ( L561, L722 ); 
   nand2 U631 ( L1689, L1692, L1023 ); 
   nand2 U632 ( L1777, L1780, L1147 ); 
   nand2 U633 ( L416, L417, L418 ); 
   nand2 U634 ( L1373, L1376, L420 ); 
   nand2 U635 ( L423, L424, L425 ); 
   nand2 U636 ( L508, L509, L510 ); 
   nand2 U637 ( L511, L512, L513 ); 
   inv U638 ( L546, L552 ); 
   nand2 U639 ( L1023, L1024, L1025 ); 
   nand2 U640 ( L1147, L1148, L1149 ); 
   inv U641 ( L418, L419 ); 
   nand2 U642 ( L420, L421, L422 ); 
   nand2 U643 ( L425, L918, L441 ); 
   inv U644 ( L510, L516 ); 
   inv U645 ( L549, L725 ); 
   buffer U646 ( L549, L728 ); 
   inv U647 ( L1025, L1029 ); 
   inv U648 ( L1149, L1153 ); 
   nand2 U649 ( L419, L918, L433 ); 
   nand2 U650 ( L422, L918, L437 ); 
   inv U651 ( L513, L663 ); 
   buffer U652 ( L513, L666 ); 
   and2 U653 ( L719, L725, L731 ); 
   and2 U654 ( L722, L725, L746 ); 
   and2 U655 ( L719, L728, L756 ); 
   and2 U656 ( L722, L728, L770 ); 
   buffer U657 ( L441, L1461 ); 
   buffer U658 ( L441, L1469 ); 
   buffer U659 ( L433, L1413 ); 
   buffer U660 ( L433, L1421 ); 
   buffer U661 ( L437, L1445 ); 
   buffer U662 ( L437, L1453 ); 
   nand2 U663 ( L1469, L1472, L532 ); 
   inv U664 ( L1469, L1473 ); 
   nand2 U665 ( L1461, L1464, L535 ); 
   inv U666 ( L1461, L1465 ); 
   nand2 U667 ( L1421, L1424, L495 ); 
   inv U668 ( L1421, L1425 ); 
   nand2 U669 ( L1413, L1416, L498 ); 
   inv U670 ( L1413, L1417 ); 
   nand2 U671 ( L1453, L1456, L520 ); 
   inv U672 ( L1453, L1457 ); 
   nand2 U673 ( L1445, L1448, L523 ); 
   inv U674 ( L1445, L1449 ); 
   nand2 U675 ( L1466, L1473, L533 ); 
   nand2 U676 ( L1458, L1465, L536 ); 
   nand2 U677 ( L1418, L1425, L496 ); 
   nand2 U678 ( L1410, L1417, L499 ); 
   nand2 U679 ( L1450, L1457, L521 ); 
   nand2 U680 ( L1442, L1449, L524 ); 
   nand2 U681 ( L532, L533, L534 ); 
   nand2 U682 ( L535, L536, L537 ); 
   nand2 U683 ( L495, L496, L497 ); 
   nand2 U684 ( L498, L499, L500 ); 
   nand2 U685 ( L520, L521, L522 ); 
   nand2 U686 ( L523, L524, L525 ); 
   inv U687 ( L534, L540 ); 
   inv U688 ( L497, L503 ); 
   inv U689 ( L522, L528 ); 
   inv U690 ( L537, L669 ); 
   buffer U691 ( L537, L672 ); 
   inv U692 ( L500, L569 ); 
   and2 U693 ( L566, L500, L588 ); 
   inv U694 ( L525, L618 ); 
   and2 U695 ( L615, L525, L639 ); 
   nand8 U696 ( L516, L564, L552, L540, L482, L528, L503, L487, L867 ); 
   buffer U697 ( L588, L588a ); 
   buffer U698 ( L588, L588b ); 
   buffer U699 ( L639, L639a ); 
   buffer U700 ( L639, L639b ); 
   and2 U701 ( L663, L669, L675 ); 
   and2 U702 ( L666, L669, L688 ); 
   and2 U703 ( L663, L672, L696 ); 
   and2 U704 ( L666, L672, L710 ); 
   and3 U705 ( L949, L867, L932, L73 ); 
   and2 U706 ( L565, L569, L572 ); 
   and2 U707 ( L566, L569, L573 ); 
   and2 U708 ( L614, L618, L621 ); 
   and2 U709 ( L615, L618, L622 ); 
   nand5 U710 ( L588a, L639a, L696, L731, L958, L776 ); 
   nand5 U711 ( L588a, L639a, L675, L756, L958, L780 ); 
   nand5 U712 ( L588a, L639a, L675, L746, L958, L784 ); 
   nand5 U713 ( L588a, L639a, L688, L731, L958, L788 ); 
   nand5 U714 ( L588b, L639a, L710, L746, L969, L812 ); 
   nand5 U715 ( L588b, L639b, L696, L770, L969, L832 ); 
   nand5 U716 ( L588b, L639b, L710, L756, L969, L836 ); 
   and5 U717 ( L588a, L639a, L696, L731, L958, L1509 ); 
   and5 U718 ( L588a, L639a, L675, L756, L958, L1517 ); 
   and5 U719 ( L588a, L639a, L675, L746, L958, L1525 ); 
   and5 U720 ( L588a, L639a, L688, L731, L958, L1533 ); 
   and5 U721 ( L588b, L639a, L710, L746, L969, L1581 ); 
   and5 U722 ( L588b, L639b, L696, L770, L969, L1621 ); 
   and5 U723 ( L588b, L639b, L710, L756, L969, L1629 ); 
   nand5 U724 ( L588a, L622, L696, L756, L958, L792 ); 
   nand5 U725 ( L588b, L622, L696, L746, L958, L796 ); 
   nand5 U726 ( L588b, L622, L710, L731, L958, L800 ); 
   nand5 U727 ( L588b, L622, L675, L770, L958, L804 ); 
   nand5 U728 ( L588b, L622, L688, L756, L969, L808 ); 
   nand5 U729 ( L573, L639b, L696, L756, L969, L816 ); 
   nand5 U730 ( L573, L639b, L696, L746, L969, L820 ); 
   nand5 U731 ( L573, L639b, L710, L731, L969, L824 ); 
   nand5 U732 ( L573, L639b, L688, L756, L969, L828 ); 
   nand5 U733 ( L588b, L622, L675, L731, L979, L871 ); 
   nand5 U734 ( L573, L639b, L675, L731, L979, L873 ); 
   nand5 U735 ( L573, L622, L696, L731, L979, L875 ); 
   nand5 U736 ( L573, L622, L675, L756, L979, L877 ); 
   nand5 U737 ( L573, L622, L675, L746, L979, L879 ); 
   nand5 U738 ( L573, L622, L688, L731, L979, L881 ); 
   nand5 U739 ( L573, L621, L675, L731, L979, L883 ); 
   nand5 U740 ( L572, L622, L675, L731, L979, L885 ); 
   and5 U741 ( L588a, L622, L696, L756, L958, L1541 ); 
   and5 U742 ( L588b, L622, L696, L746, L958, L1549 ); 
   and5 U743 ( L588b, L622, L710, L731, L958, L1557 ); 
   and5 U744 ( L588b, L622, L675, L770, L958, L1565 ); 
   and5 U745 ( L588b, L622, L688, L756, L969, L1573 ); 
   and5 U746 ( L573, L639b, L696, L756, L969, L1589 ); 
   and5 U747 ( L573, L639b, L696, L746, L969, L1597 ); 
   and5 U748 ( L573, L639b, L710, L731, L969, L1605 ); 
   and5 U749 ( L573, L639b, L688, L756, L969, L1613 ); 
   nand2 U750 ( L1509, L1512, L1 ); 
   inv U751 ( L1509, L1513 ); 
   nand2 U752 ( L1517, L1520, L4 ); 
   inv U753 ( L1517, L1521 ); 
   nand2 U754 ( L1525, L1528, L7 ); 
   inv U755 ( L1525, L1529 ); 
   nand2 U756 ( L1533, L1536, L10 ); 
   inv U757 ( L1533, L1537 ); 
   nand2 U758 ( L1581, L1584, L28 ); 
   inv U759 ( L1581, L1585 ); 
   nand2 U760 ( L1621, L1624, L43 ); 
   inv U761 ( L1621, L1625 ); 
   nand2 U762 ( L1629, L1632, L46 ); 
   inv U763 ( L1629, L1633 ); 
   and8 U764 ( L871, L873, L875, L877, L879, L881, L883, L885, L886 ); 
   nand2 U765 ( L1506, L1513, L2 ); 
   nand2 U766 ( L1514, L1521, L5 ); 
   nand2 U767 ( L1522, L1529, L8 ); 
   nand2 U768 ( L1530, L1537, L11 ); 
   nand2 U769 ( L1541, L1544, L13 ); 
   inv U770 ( L1541, L1545 ); 
   nand2 U771 ( L1549, L1552, L16 ); 
   inv U772 ( L1549, L1553 ); 
   nand2 U773 ( L1557, L1560, L19 ); 
   inv U774 ( L1557, L1561 ); 
   nand2 U775 ( L1565, L1568, L22 ); 
   inv U776 ( L1565, L1569 ); 
   nand2 U777 ( L1573, L1576, L25 ); 
   inv U778 ( L1573, L1577 ); 
   nand2 U779 ( L1578, L1585, L29 ); 
   nand2 U780 ( L1589, L1592, L31 ); 
   inv U781 ( L1589, L1593 ); 
   nand2 U782 ( L1597, L1600, L34 ); 
   inv U783 ( L1597, L1601 ); 
   nand2 U784 ( L1605, L1608, L37 ); 
   inv U785 ( L1605, L1609 ); 
   nand2 U786 ( L1613, L1616, L40 ); 
   inv U787 ( L1613, L1617 ); 
   nand2 U788 ( L1618, L1625, L44 ); 
   nand2 U789 ( L1626, L1633, L47 ); 
   nand8 U790 ( L776, L780, L784, L788, L792, L796, L800, L804, L857 ); 
   nand8 U791 ( L808, L812, L816, L820, L824, L828, L832, L836, L860 ); 
   and8 U792 ( L776, L780, L784, L788, L792, L796, L800, L804, L863 ); 
   and8 U793 ( L808, L812, L816, L820, L824, L828, L832, L836, L865 ); 
   nand2 U794 ( L1, L2, L3 ); 
   nand2 U795 ( L4, L5, L6 ); 
   nand2 U796 ( L7, L8, L9 ); 
   nand2 U797 ( L10, L11, L12 ); 
   nand2 U798 ( L1538, L1545, L14 ); 
   nand2 U799 ( L1546, L1553, L17 ); 
   nand2 U800 ( L1554, L1561, L20 ); 
   nand2 U801 ( L1562, L1569, L23 ); 
   nand2 U802 ( L1570, L1577, L26 ); 
   nand2 U803 ( L28, L29, L30 ); 
   nand2 U804 ( L1586, L1593, L32 ); 
   nand2 U805 ( L1594, L1601, L35 ); 
   nand2 U806 ( L1602, L1609, L38 ); 
   nand2 U807 ( L1610, L1617, L41 ); 
   nand2 U808 ( L43, L44, L45 ); 
   nand2 U809 ( L46, L47, L48 ); 
   and2 U810 ( L857, L859, L1913 ); 
   and2 U811 ( L860, L862, L1921 ); 
   nand2 U812 ( L13, L14, L15 ); 
   nand2 U813 ( L16, L17, L18 ); 
   nand2 U814 ( L19, L20, L21 ); 
   nand2 U815 ( L22, L23, L24 ); 
   nand2 U816 ( L25, L26, L27 ); 
   nand2 U817 ( L31, L32, L33 ); 
   nand2 U818 ( L34, L35, L36 ); 
   nand2 U819 ( L37, L38, L39 ); 
   nand2 U820 ( L40, L41, L42 ); 
   and3 U821 ( L863, L865, L886, L887 ); 
   nand2 U822 ( L863, L865, L462 ); 
   and4 U823 ( L949, L867, L952, L887, L74 ); 
   nand2 U824 ( L1913, L1916, L1637 ); 
   inv U825 ( L1913, L1917 ); 
   nand2 U826 ( L1921, L1924, L1647 ); 
   inv U827 ( L1921, L1925 ); 
   nor2 U828 ( L73, L74, L75 ); 
   and3 U829 ( L457, L911, L462, L1020 ); 
   and3 U830 ( L469, L911, L462, L1144 ); 
   and3 U831 ( L475, L911, L462, L1386 ); 
   and3 U832 ( L478, L911, L462, L1394 ); 
   and3 U833 ( L459, L911, L462, L1402 ); 
   nand2 U834 ( L1910, L1917, L1638 ); 
   nand2 U835 ( L1918, L1925, L1648 ); 
   and3 U836 ( L472, L911, L462, L1806 ); 
   nand2 U837 ( L1637, L1638, L1639 ); 
   nand2 U838 ( L1647, L1648, L1649 ); 
   nand2 U839 ( L1020, L1029, L287 ); 
   nand2 U840 ( L1144, L1153, L350 ); 
   nand2 U841 ( L1386, L1393, L427 ); 
   nand2 U842 ( L1394, L1401, L429 ); 
   nand2 U843 ( L1402, L1409, L431 ); 
   inv U844 ( L1020, L1028 ); 
   inv U845 ( L1144, L1152 ); 
   inv U846 ( L1386, L1392 ); 
   inv U847 ( L1394, L1400 ); 
   inv U848 ( L1402, L1408 ); 
   inv U849 ( L1806, L1812 ); 
   nand2 U850 ( L1806, L1813, L1216 ); 
   nand2 U851 ( L1025, L1028, L286 ); 
   nand2 U852 ( L1149, L1152, L349 ); 
   nand2 U853 ( L1389, L1392, L426 ); 
   nand2 U854 ( L1397, L1400, L428 ); 
   nand2 U855 ( L1405, L1408, L430 ); 
   nand2 U856 ( L1639, L1642, L67 ); 
   inv U857 ( L1639, L1643 ); 
   nand2 U858 ( L1649, L1652, L70 ); 
   inv U859 ( L1649, L1653 ); 
   nand2 U860 ( L1809, L1812, L1215 ); 
   nand2 U861 ( L286, L287, L49 ); 
   nand2 U862 ( L349, L350, L53 ); 
   nand2 U863 ( L426, L427, L59 ); 
   nand2 U864 ( L428, L429, L61 ); 
   nand2 U865 ( L430, L431, L65 ); 
   nand2 U866 ( L1634, L1643, L68 ); 
   nand2 U867 ( L1644, L1653, L71 ); 
   nand2 U868 ( L1215, L1216, L1217 ); 
   and2 U869 ( L49, L50, L51 ); 
   and2 U870 ( L52, L53, L54 ); 
   and2 U871 ( L58, L59, L60 ); 
   and2 U872 ( L61, L62, L63 ); 
   and2 U873 ( L64, L65, L66 ); 
   nand2 U874 ( L67, L68, L69 ); 
   nand2 U875 ( L70, L71, L72 ); 
   nand2 U876 ( L1217, L1220, L375 ); 
   inv U877 ( L1217, L1221 ); 
   nand2 U878 ( L1212, L1221, L376 ); 
   nand2 U879 ( L375, L376, L55 ); 
   and2 U880 ( L55, L56, L57 ); 
endmodule

