module top( pi000 , pi001 , pi002 , pi003 , pi004 , pi005 , pi006 , pi007 , pi008 , pi009 , pi010 , pi011 , pi012 , pi013 , pi014 , pi015 , pi016 , pi017 , pi018 , pi019 , pi020 , pi021 , pi022 , pi023 , pi024 , pi025 , pi026 , pi027 , pi028 , pi029 , pi030 , pi031 , pi032 , pi033 , pi034 , pi035 , pi036 , pi037 , pi038 , pi039 , pi040 , pi041 , pi042 , pi043 , pi044 , pi045 , pi046 , pi047 , pi048 , pi049 , pi050 , pi051 , pi052 , pi053 , pi054 , pi055 , pi056 , pi057 , pi058 , pi059 , pi060 , pi061 , pi062 , pi063 , pi064 , pi065 , pi066 , pi067 , pi068 , pi069 , pi070 , pi071 , pi072 , pi073 , pi074 , pi075 , pi076 , pi077 , pi078 , pi079 , pi080 , pi081 , pi082 , pi083 , pi084 , pi085 , pi086 , pi087 , pi088 , pi089 , pi090 , pi091 , pi092 , pi093 , pi094 , pi095 , pi096 , pi097 , pi098 , pi099 , pi100 , pi101 , pi102 , pi103 , pi104 , pi105 , pi106 , pi107 , pi108 , pi109 , pi110 , pi111 , pi112 , pi113 , pi114 , pi115 , pi116 , pi117 , pi118 , pi119 , pi120 , pi121 , pi122 , pi123 , pi124 , pi125 , pi126 , pi127 , pi128 , pi129 , pi130 , pi131 , pi132 , pi133 , pi134 , pi135 , pi136 , pi137 , pi138 , pi139 , pi140 , pi141 , pi142 , pi143 , pi144 , pi145 , pi146 , pi147 , pi148 , pi149 , pi150 , pi151 , pi152 , pi153 , pi154 , pi155 , pi156 , pi157 , pi158 , pi159 , pi160 , pi161 , pi162 , pi163 , pi164 , pi165 , pi166 , pi167 , pi168 , pi169 , pi170 , pi171 , pi172 , pi173 , pi174 , pi175 , pi176 , pi177 , pi178 , pi179 , pi180 , pi181 , pi182 , pi183 , pi184 , pi185 , pi186 , pi187 , pi188 , pi189 , pi190 , pi191 , pi192 , pi193 , pi194 , pi195 , pi196 , pi197 , pi198 , pi199 , pi200 , pi201 , pi202 , pi203 , pi204 , pi205 , pi206 , pi207 , pi208 , pi209 , pi210 , pi211 , pi212 , pi213 , pi214 , pi215 , pi216 , pi217 , pi218 , pi219 , pi220 , pi221 , pi222 , pi223 , pi224 , pi225 , pi226 , pi227 , pi228 , pi229 , pi230 , pi231 , pi232 , pi233 , pi234 , pi235 , pi236 , pi237 , pi238 , pi239 , pi240 , pi241 , pi242 , pi243 , pi244 , pi245 , pi246 , pi247 , pi248 , pi249 , pi250 , pi251 , pi252 , pi253 , pi254 , pi255 , pi256 , pi257 , pi258 , pi259 , pi260 , pi261 , pi262 , pi263 , pi264 , pi265 , pi266 , pi267 , pi268 , pi269 , pi270 , pi271 , pi272 , pi273 , pi274 , pi275 , pi276 , pi277 , pi278 , pi279 , pi280 , pi281 , pi282 , pi283 , pi284 , pi285 , pi286 , pi287 , pi288 , pi289 , pi290 , pi291 , pi292 , pi293 , pi294 , pi295 , pi296 , pi297 , pi298 , pi299 , pi300 , pi301 , pi302 , pi303 , pi304 , pi305 , pi306 , pi307 , pi308 , pi309 , pi310 , pi311 , pi312 , pi313 , pi314 , pi315 , pi316 , pi317 , pi318 , pi319 , pi320 , pi321 , pi322 , pi323 , pi324 , pi325 , pi326 , pi327 , pi328 , pi329 , pi330 , pi331 , pi332 , pi333 , pi334 , pi335 , pi336 , pi337 , pi338 , pi339 , pi340 , pi341 , pi342 , pi343 , pi344 , pi345 , pi346 , pi347 , pi348 , pi349 , pi350 , pi351 , pi352 , pi353 , pi354 , pi355 , pi356 , pi357 , pi358 , pi359 , pi360 , pi361 , pi362 , pi363 , pi364 , pi365 , pi366 , pi367 , pi368 , pi369 , pi370 , pi371 , pi372 , pi373 , pi374 , pi375 , pi376 , pi377 , pi378 , pi379 , pi380 , pi381 , pi382 , pi383 , pi384 , pi385 , pi386 , pi387 , pi388 , pi389 , pi390 , pi391 , pi392 , pi393 , pi394 , pi395 , pi396 , pi397 , pi398 , pi399 , pi400 , pi401 , pi402 , pi403 , pi404 , pi405 , pi406 , pi407 , pi408 , pi409 , pi410 , pi411 , pi412 , pi413 , pi414 , pi415 , pi416 , pi417 , pi418 , pi419 , pi420 , pi421 , pi422 , pi423 , pi424 , pi425 , pi426 , pi427 , pi428 , pi429 , pi430 , pi431 , pi432 , pi433 , pi434 , pi435 , pi436 , pi437 , pi438 , pi439 , pi440 , pi441 , pi442 , pi443 , pi444 , pi445 , pi446 , pi447 , pi448 , pi449 , pi450 , pi451 , pi452 , pi453 , pi454 , pi455 , pi456 , pi457 , pi458 , pi459 , pi460 , pi461 , pi462 , pi463 , po0000 , po0001 , po0002 , po0003 , po0004 , po0005 , po0006 , po0007 , po0008 , po0009 , po0010 , po0011 , po0012 , po0013 , po0014 , po0015 , po0016 , po0017 , po0018 , po0019 , po0020 , po0021 , po0022 , po0023 , po0024 , po0025 , po0026 , po0027 , po0028 , po0029 , po0030 , po0031 , po0032 , po0033 , po0034 , po0035 , po0036 , po0037 , po0038 , po0039 , po0040 , po0041 , po0042 , po0043 , po0044 , po0045 , po0046 , po0047 , po0048 , po0049 , po0050 , po0051 , po0052 , po0053 , po0054 , po0055 , po0056 , po0057 , po0058 , po0059 , po0060 , po0061 , po0062 , po0063 , po0064 , po0065 , po0066 , po0067 , po0068 , po0069 , po0070 , po0071 , po0072 , po0073 , po0074 , po0075 , po0076 , po0077 , po0078 , po0079 , po0080 , po0081 , po0082 , po0083 , po0084 , po0085 , po0086 , po0087 , po0088 , po0089 , po0090 , po0091 , po0092 , po0093 , po0094 , po0095 , po0096 , po0097 , po0098 , po0099 , po0100 , po0101 , po0102 , po0103 , po0104 , po0105 , po0106 , po0107 , po0108 , po0109 , po0110 , po0111 , po0112 , po0113 , po0114 , po0115 , po0116 , po0117 , po0118 , po0119 , po0120 , po0121 , po0122 , po0123 , po0124 , po0125 , po0126 , po0127 , po0128 , po0129 , po0130 , po0131 , po0132 , po0133 , po0134 , po0135 , po0136 , po0137 , po0138 , po0139 , po0140 , po0141 , po0142 , po0143 , po0144 , po0145 , po0146 , po0147 , po0148 , po0149 , po0150 , po0151 , po0152 , po0153 , po0154 , po0155 , po0156 , po0157 , po0158 , po0159 , po0160 , po0161 , po0162 , po0163 , po0164 , po0165 , po0166 , po0167 , po0168 , po0169 , po0170 , po0171 , po0172 , po0173 , po0174 , po0175 , po0176 , po0177 , po0178 , po0179 , po0180 , po0181 , po0182 , po0183 , po0184 , po0185 , po0186 , po0187 , po0188 , po0189 , po0190 , po0191 , po0192 , po0193 , po0194 , po0195 , po0196 , po0197 , po0198 , po0199 , po0200 , po0201 , po0202 , po0203 , po0204 , po0205 , po0206 , po0207 , po0208 , po0209 , po0210 , po0211 , po0212 , po0213 , po0214 , po0215 , po0216 , po0217 , po0218 , po0219 , po0220 , po0221 , po0222 , po0223 , po0224 , po0225 , po0226 , po0227 , po0228 , po0229 , po0230 , po0231 , po0232 , po0233 , po0234 , po0235 , po0236 , po0237 , po0238 , po0239 , po0240 , po0241 , po0242 , po0243 , po0244 , po0245 , po0246 , po0247 , po0248 , po0249 , po0250 , po0251 , po0252 , po0253 , po0254 , po0255 , po0256 , po0257 , po0258 , po0259 , po0260 , po0261 , po0262 , po0263 , po0264 , po0265 , po0266 , po0267 , po0268 , po0269 , po0270 , po0271 , po0272 , po0273 , po0274 , po0275 , po0276 , po0277 , po0278 , po0279 , po0280 , po0281 , po0282 , po0283 , po0284 , po0285 , po0286 , po0287 , po0288 , po0289 , po0290 , po0291 , po0292 , po0293 , po0294 , po0295 , po0296 , po0297 , po0298 , po0299 , po0300 , po0301 , po0302 , po0303 , po0304 , po0305 , po0306 , po0307 , po0308 , po0309 , po0310 , po0311 , po0312 , po0313 , po0314 , po0315 , po0316 , po0317 , po0318 , po0319 , po0320 , po0321 , po0322 , po0323 , po0324 , po0325 , po0326 , po0327 , po0328 , po0329 , po0330 , po0331 , po0332 , po0333 , po0334 , po0335 , po0336 , po0337 , po0338 , po0339 , po0340 , po0341 , po0342 , po0343 , po0344 , po0345 , po0346 , po0347 , po0348 , po0349 , po0350 , po0351 , po0352 , po0353 , po0354 , po0355 , po0356 , po0357 , po0358 , po0359 , po0360 , po0361 , po0362 , po0363 , po0364 , po0365 , po0366 , po0367 , po0368 , po0369 , po0370 , po0371 , po0372 , po0373 , po0374 , po0375 , po0376 , po0377 , po0378 , po0379 , po0380 , po0381 , po0382 , po0383 , po0384 , po0385 , po0386 , po0387 , po0388 , po0389 , po0390 , po0391 , po0392 , po0393 , po0394 , po0395 , po0396 , po0397 , po0398 , po0399 , po0400 , po0401 , po0402 , po0403 , po0404 , po0405 , po0406 , po0407 , po0408 , po0409 , po0410 , po0411 , po0412 , po0413 , po0414 , po0415 , po0416 , po0417 , po0418 , po0419 , po0420 , po0421 , po0422 , po0423 , po0424 , po0425 , po0426 , po0427 , po0428 , po0429 , po0430 , po0431 , po0432 , po0433 , po0434 , po0435 , po0436 , po0437 , po0438 , po0439 , po0440 , po0441 , po0442 , po0443 , po0444 , po0445 , po0446 , po0447 , po0448 , po0449 , po0450 , po0451 , po0452 , po0453 , po0454 , po0455 , po0456 , po0457 , po0458 , po0459 , po0460 , po0461 , po0462 , po0463 , po0464 , po0465 , po0466 , po0467 , po0468 , po0469 , po0470 , po0471 , po0472 , po0473 , po0474 , po0475 , po0476 , po0477 , po0478 , po0479 , po0480 , po0481 , po0482 , po0483 , po0484 , po0485 , po0486 , po0487 , po0488 , po0489 , po0490 , po0491 , po0492 , po0493 , po0494 , po0495 , po0496 , po0497 , po0498 , po0499 , po0500 , po0501 , po0502 , po0503 , po0504 , po0505 , po0506 , po0507 , po0508 , po0509 , po0510 , po0511 , po0512 , po0513 , po0514 , po0515 , po0516 , po0517 , po0518 , po0519 , po0520 , po0521 , po0522 , po0523 , po0524 , po0525 , po0526 , po0527 , po0528 , po0529 , po0530 , po0531 , po0532 , po0533 , po0534 , po0535 , po0536 , po0537 , po0538 , po0539 , po0540 , po0541 , po0542 , po0543 , po0544 , po0545 , po0546 , po0547 , po0548 , po0549 , po0550 , po0551 , po0552 , po0553 , po0554 , po0555 , po0556 , po0557 , po0558 , po0559 , po0560 , po0561 , po0562 , po0563 , po0564 , po0565 , po0566 , po0567 , po0568 , po0569 , po0570 , po0571 , po0572 , po0573 , po0574 , po0575 , po0576 , po0577 , po0578 , po0579 , po0580 , po0581 , po0582 , po0583 , po0584 , po0585 , po0586 , po0587 , po0588 , po0589 , po0590 , po0591 , po0592 , po0593 , po0594 , po0595 , po0596 , po0597 , po0598 , po0599 , po0600 , po0601 , po0602 , po0603 , po0604 , po0605 , po0606 , po0607 , po0608 , po0609 , po0610 , po0611 , po0612 , po0613 , po0614 , po0615 , po0616 , po0617 , po0618 , po0619 , po0620 , po0621 , po0622 , po0623 , po0624 , po0625 , po0626 , po0627 , po0628 , po0629 , po0630 , po0631 , po0632 , po0633 , po0634 , po0635 , po0636 , po0637 , po0638 , po0639 , po0640 , po0641 , po0642 , po0643 , po0644 , po0645 , po0646 , po0647 , po0648 , po0649 , po0650 , po0651 , po0652 , po0653 , po0654 , po0655 , po0656 , po0657 , po0658 , po0659 , po0660 , po0661 , po0662 , po0663 , po0664 , po0665 , po0666 , po0667 , po0668 , po0669 , po0670 , po0671 , po0672 , po0673 , po0674 , po0675 , po0676 , po0677 , po0678 , po0679 , po0680 , po0681 , po0682 , po0683 , po0684 , po0685 , po0686 , po0687 , po0688 , po0689 , po0690 , po0691 , po0692 , po0693 , po0694 , po0695 , po0696 , po0697 , po0698 , po0699 , po0700 , po0701 , po0702 , po0703 , po0704 , po0705 , po0706 , po0707 , po0708 , po0709 , po0710 , po0711 , po0712 , po0713 , po0714 , po0715 , po0716 , po0717 , po0718 , po0719 , po0720 , po0721 , po0722 , po0723 , po0724 , po0725 , po0726 , po0727 , po0728 , po0729 , po0730 , po0731 , po0732 , po0733 , po0734 , po0735 , po0736 , po0737 , po0738 , po0739 , po0740 , po0741 , po0742 , po0743 , po0744 , po0745 , po0746 , po0747 , po0748 , po0749 , po0750 , po0751 , po0752 , po0753 , po0754 , po0755 , po0756 , po0757 , po0758 , po0759 , po0760 , po0761 , po0762 , po0763 , po0764 , po0765 , po0766 , po0767 , po0768 , po0769 , po0770 , po0771 , po0772 , po0773 , po0774 , po0775 , po0776 , po0777 , po0778 , po0779 , po0780 , po0781 , po0782 , po0783 , po0784 , po0785 , po0786 , po0787 , po0788 , po0789 , po0790 , po0791 , po0792 , po0793 , po0794 , po0795 , po0796 , po0797 , po0798 , po0799 , po0800 , po0801 , po0802 , po0803 , po0804 , po0805 , po0806 , po0807 , po0808 , po0809 , po0810 , po0811 , po0812 , po0813 , po0814 , po0815 , po0816 , po0817 , po0818 , po0819 , po0820 , po0821 , po0822 , po0823 , po0824 , po0825 , po0826 , po0827 , po0828 , po0829 , po0830 , po0831 , po0832 , po0833 , po0834 , po0835 , po0836 , po0837 , po0838 , po0839 , po0840 , po0841 , po0842 , po0843 , po0844 , po0845 , po0846 , po0847 , po0848 , po0849 , po0850 , po0851 , po0852 , po0853 , po0854 , po0855 , po0856 , po0857 , po0858 , po0859 , po0860 , po0861 , po0862 , po0863 , po0864 , po0865 , po0866 , po0867 , po0868 , po0869 , po0870 , po0871 , po0872 , po0873 , po0874 , po0875 , po0876 , po0877 , po0878 , po0879 , po0880 , po0881 , po0882 , po0883 , po0884 , po0885 , po0886 , po0887 , po0888 , po0889 , po0890 , po0891 , po0892 , po0893 , po0894 , po0895 , po0896 , po0897 , po0898 , po0899 , po0900 , po0901 , po0902 , po0903 , po0904 , po0905 , po0906 , po0907 , po0908 , po0909 , po0910 , po0911 , po0912 , po0913 , po0914 , po0915 , po0916 , po0917 , po0918 , po0919 , po0920 , po0921 , po0922 , po0923 , po0924 , po0925 , po0926 , po0927 , po0928 , po0929 , po0930 , po0931 , po0932 , po0933 , po0934 , po0935 , po0936 , po0937 , po0938 , po0939 , po0940 , po0941 , po0942 , po0943 , po0944 , po0945 , po0946 , po0947 , po0948 , po0949 , po0950 , po0951 , po0952 , po0953 , po0954 , po0955 , po0956 , po0957 , po0958 , po0959 , po0960 , po0961 , po0962 , po0963 , po0964 , po0965 , po0966 , po0967 , po0968 , po0969 , po0970 , po0971 , po0972 , po0973 , po0974 , po0975 , po0976 , po0977 , po0978 , po0979 , po0980 , po0981 , po0982 , po0983 , po0984 , po0985 , po0986 , po0987 , po0988 , po0989 , po0990 , po0991 , po0992 , po0993 , po0994 , po0995 , po0996 , po0997 , po0998 , po0999 , po1000 , po1001 , po1002 , po1003 , po1004 , po1005 , po1006 , po1007 , po1008 , po1009 , po1010 , po1011 , po1012 , po1013 , po1014 , po1015 , po1016 , po1017 , po1018 , po1019 , po1020 , po1021 , po1022 , po1023 , po1024 , po1025 , po1026 , po1027 , po1028 , po1029 , po1030 , po1031 , po1032 , po1033 , po1034 , po1035 , po1036 , po1037 , po1038 , po1039 , po1040 , po1041 , po1042 , po1043 , po1044 , po1045 , po1046 , po1047 , po1048 , po1049 , po1050 , po1051 , po1052 , po1053 , po1054 , po1055 , po1056 , po1057 , po1058 , po1059 , po1060 , po1061 , po1062 , po1063 , po1064 , po1065 , po1066 , po1067 , po1068 , po1069 , po1070 , po1071 , po1072 , po1073 , po1074 , po1075 , po1076 , po1077 , po1078 , po1079 , po1080 , po1081 , po1082 , po1083 , po1084 , po1085 , po1086 , po1087 , po1088 , po1089 , po1090 , po1091 , po1092 , po1093 , po1094 , po1095 , po1096 , po1097 , po1098 , po1099 , po1100 , po1101 , po1102 , po1103 , po1104 , po1105 , po1106 , po1107 , po1108 , po1109 , po1110 , po1111 , po1112 , po1113 , po1114 , po1115 , po1116 , po1117 , po1118 , po1119 , po1120 , po1121 , po1122 , po1123 , po1124 , po1125 , po1126 , po1127 , po1128 , po1129 , po1130 , po1131 , po1132 , po1133 , po1134 , po1135 , po1136 , po1137 , po1138 , po1139 , po1140 , po1141 , po1142 , po1143 , po1144 , po1145 , po1146 , po1147 , po1148 , po1149 , po1150 , po1151 , po1152 , po1153 , po1154 , po1155 , po1156 , po1157 , po1158 , po1159 , po1160 , po1161 , po1162 , po1163 , po1164 , po1165 , po1166 , po1167 , po1168 , po1169 , po1170 , po1171 , po1172 , po1173 , po1174 , po1175 , po1176 , po1177 , po1178 , po1179 , po1180 , po1181 , po1182 , po1183 , po1184 , po1185 , po1186 , po1187 , po1188 , po1189 , po1190 , po1191 , po1192 , po1193 , po1194 , po1195 , po1196 , po1197 , po1198 , po1199 , po1200 , po1201 , po1202 , po1203 , po1204 , po1205 , po1206 , po1207 , po1208 , po1209 , po1210 , po1211 , po1212 , po1213 , po1214 , po1215 , po1216 , po1217 , po1218 , po1219 , po1220 , po1221 , po1222 , po1223 , po1224 , po1225 , po1226 , po1227 , po1228 , po1229 , po1230 , po1231 , po1232 , po1233 , po1234 , po1235 , po1236 , po1237 , po1238 , po1239 , po1240 , po1241 , po1242 , po1243 , po1244 , po1245 , po1246 , po1247 , po1248 , po1249 , po1250 , po1251 , po1252 , po1253 , po1254 , po1255 , po1256 , po1257 , po1258 , po1259 , po1260 , po1261 , po1262 , po1263 , po1264 , po1265 , po1266 , po1267 , po1268 , po1269 , po1270 , po1271 , po1272 , po1273 , po1274 , po1275 , po1276 , po1277 , po1278 , po1279 , po1280 , po1281 , po1282 , po1283 , po1284 , po1285 , po1286 , po1287 , po1288 , po1289 , po1290 , po1291 , po1292 , po1293 , po1294 , po1295 , po1296 , po1297 , po1298 , po1299 , po1300 , po1301 , po1302 , po1303 , po1304 , po1305 , po1306 , po1307 , po1308 , po1309 , po1310 , po1311 , po1312 , po1313 , po1314 , po1315 , po1316 , po1317 , po1318 , po1319 , po1320 , po1321 , po1322 , po1323 , po1324 , po1325 , po1326 , po1327 , po1328 , po1329 , po1330 , po1331 , po1332 , po1333 , po1334 , po1335 , po1336 , po1337 , po1338 , po1339 , po1340 , po1341 , po1342 , po1343 , po1344 , po1345 , po1346 , po1347 , po1348 , po1349 , po1350 , po1351 , po1352 , po1353 , po1354 , po1355 , po1356 , po1357 , po1358 , po1359 , po1360 , po1361 , po1362 , po1363 , po1364 , po1365 , po1366 , po1367 , po1368 , po1369 , po1370 , po1371 , po1372 , po1373 , po1374 , po1375 , po1376 , po1377 , po1378 , po1379 , po1380 , po1381 , po1382 , po1383 , po1384 , po1385 , po1386 , po1387 , po1388 , po1389 , po1390 , po1391 , po1392 , po1393 , po1394 , po1395 , po1396 , po1397 , po1398 , po1399 , po1400 , po1401 , po1402 , po1403 , po1404 , po1405 , po1406 , po1407 , po1408 , po1409 , po1410 , po1411 , po1412 , po1413 , po1414 , po1415 , po1416 , po1417 , po1418 , po1419 , po1420 , po1421 , po1422 , po1423 , po1424 , po1425 , po1426 , po1427 , po1428 , po1429 , po1430 , po1431 , po1432 , po1433 , po1434 , po1435 , po1436 , po1437 , po1438 , po1439 , po1440 , po1441 , po1442 , po1443 , po1444 , po1445 , po1446 , po1447 , po1448 , po1449 , po1450 , po1451 , po1452 , po1453 , po1454 , po1455 , po1456 , po1457 , po1458 , po1459 , po1460 , po1461 , po1462 , po1463 , po1464 , po1465 , po1466 , po1467 , po1468 , po1469 , po1470 , po1471 , po1472 , po1473 , po1474 , po1475 , po1476 , po1477 , po1478 , po1479 , po1480 , po1481 , po1482 , po1483 , po1484 , po1485 , po1486 , po1487 , po1488 , po1489 , po1490 , po1491 , po1492 , po1493 , po1494 , po1495 , po1496 , po1497 , po1498 , po1499 , po1500 , po1501 , po1502 , po1503 , po1504 , po1505 , po1506 , po1507 , po1508 , po1509 , po1510 , po1511 , po1512 , po1513 , po1514 , po1515 , po1516 , po1517 , po1518 , po1519 , po1520 , po1521 , po1522 , po1523 , po1524 , po1525 , po1526 , po1527 , po1528 , po1529 , po1530 , po1531 , po1532 , po1533 , po1534 , po1535 , po1536 , po1537 , po1538 , po1539 , po1540 , po1541 , po1542 , po1543 , po1544 , po1545 , po1546 , po1547 , po1548 , po1549 , po1550 , po1551 , po1552 , po1553 , po1554 , po1555 , po1556 , po1557 , po1558 , po1559 , po1560 , po1561 , po1562 , po1563 , po1564 , po1565 , po1566 , po1567 , po1568 , po1569 , po1570 , po1571 , po1572 , po1573 , po1574 , po1575 , po1576 , po1577 , po1578 , po1579 , po1580 , po1581 , po1582 , po1583 , po1584 , po1585 , po1586 , po1587 , po1588 , po1589 , po1590 , po1591 , po1592 , po1593 , po1594 , po1595 , po1596 , po1597 , po1598 , po1599 , po1600 , po1601 , po1602 , po1603 , po1604 , po1605 , po1606 , po1607 , po1608 , po1609 , po1610 , po1611 , po1612 , po1613 , po1614 , po1615 , po1616 , po1617 , po1618 , po1619 , po1620 , po1621 , po1622 , po1623 , po1624 , po1625 , po1626 , po1627 , po1628 , po1629 , po1630 , po1631 , po1632 , po1633 , po1634 , po1635 , po1636 , po1637 , po1638 , po1639 , po1640 , po1641 , po1642 , po1643 , po1644 , po1645 , po1646 , po1647 , po1648 , po1649 , po1650 , po1651 , po1652 , po1653 , po1654 , po1655 , po1656 , po1657 , po1658 , po1659 , po1660 , po1661 , po1662 , po1663 , po1664 , po1665 , po1666 , po1667 , po1668 , po1669 , po1670 , po1671 , po1672 , po1673 , po1674 , po1675 , po1676 , po1677 , po1678 , po1679 , po1680 , po1681 , po1682 , po1683 , po1684 , po1685 , po1686 , po1687 , po1688 , po1689 , po1690 , po1691 , po1692 , po1693 , po1694 , po1695 , po1696 , po1697 , po1698 , po1699 , po1700 , po1701 , po1702 , po1703 , po1704 , po1705 , po1706 , po1707 , po1708 , po1709 , po1710 , po1711 , po1712 , po1713 , po1714 , po1715 , po1716 , po1717 , po1718 , po1719 , po1720 , po1721 , po1722 , po1723 , po1724 , po1725 , po1726 , po1727 , po1728 , po1729 , po1730 , po1731 , po1732 , po1733 , po1734 , po1735 , po1736 , po1737 , po1738 , po1739 , po1740 , po1741 , po1742 , po1743 , po1744 , po1745 , po1746 , po1747 , po1748 , po1749 , po1750 , po1751 , po1752 , po1753 , po1754 , po1755 , po1756 , po1757 , po1758 , po1759 , po1760 , po1761 , po1762 , po1763 , po1764 , po1765 , po1766 , po1767 , po1768 , po1769 , po1770 , po1771 , po1772 , po1773 , po1774 , po1775 , po1776 , po1777 , po1778 , po1779 , po1780 , po1781 , po1782 , po1783 , po1784 , po1785 , po1786 , po1787 , po1788 , po1789 , po1790 , po1791 , po1792 , po1793 , po1794 , po1795 , po1796 , po1797 , po1798 , po1799 , po1800 , po1801 , po1802 , po1803 , po1804 , po1805 , po1806 , po1807 , po1808 , po1809 , po1810 , po1811 , po1812 , po1813 , po1814 , po1815 , po1816 , po1817 , po1818 , po1819 , po1820 , po1821 , po1822 , po1823 , po1824 , po1825 , po1826 , po1827 , po1828 , po1829 , po1830 , po1831 , po1832 , po1833 , po1834 , po1835 , po1836 , po1837 , po1838 , po1839 , po1840 , po1841 , po1842 , po1843 , po1844 , po1845 , po1846 , po1847 , po1848 , po1849 , po1850 , po1851 , po1852 , po1853 , po1854 , po1855 , po1856 , po1857 , po1858 , po1859 , po1860 , po1861 , po1862 , po1863 , po1864 , po1865 , po1866 , po1867 , po1868 , po1869 , po1870 , po1871 , po1872 , po1873 , po1874 , po1875 , po1876 , po1877 , po1878 , po1879 , po1880 , po1881 , po1882 , po1883 , po1884 , po1885 , po1886 , po1887 , po1888 , po1889 , po1890 , po1891 , po1892 , po1893 , po1894 , po1895 , po1896 , po1897 , po1898 , po1899 , po1900 , po1901 , po1902 , po1903 , po1904 , po1905 , po1906 , po1907 , po1908 , po1909 , po1910 , po1911 , po1912 , po1913 , po1914 , po1915 , po1916 , po1917 , po1918 , po1919 , po1920 , po1921 , po1922 , po1923 , po1924 , po1925 , po1926 , po1927 , po1928 , po1929 , po1930 , po1931 , po1932 , po1933 , po1934 , po1935 , po1936 , po1937 , po1938 , po1939 , po1940 , po1941 , po1942 , po1943 , po1944 , po1945 , po1946 , po1947 , po1948 , po1949 , po1950 , po1951 , po1952 , po1953 , po1954 , po1955 , po1956 , po1957 , po1958 , po1959 , po1960 , po1961 , po1962 , po1963 , po1964 , po1965 , po1966 , po1967 , po1968 , po1969 , po1970 , po1971 , po1972 , po1973 , po1974 , po1975 , po1976 , po1977 , po1978 , po1979 , po1980 , po1981 , po1982 , po1983 , po1984 , po1985 , po1986 , po1987 , po1988 , po1989 , po1990 , po1991 , po1992 , po1993 , po1994 , po1995 , po1996 , po1997 , po1998 , po1999 , po2000 , po2001 , po2002 , po2003 , po2004 , po2005 , po2006 , po2007 , po2008 , po2009 , po2010 , po2011 , po2012 , po2013 , po2014 , po2015 , po2016 , po2017 , po2018 , po2019 , po2020 , po2021 , po2022 , po2023 , po2024 , po2025 , po2026 , po2027 , po2028 , po2029 , po2030 , po2031 , po2032 , po2033 , po2034 , po2035 , po2036 , po2037 , po2038 , po2039 , po2040 , po2041 , po2042 , po2043 , po2044 , po2045 , po2046 , po2047 , po2048 , po2049 , po2050 , po2051 , po2052 , po2053 , po2054 , po2055 , po2056 , po2057 , po2058 , po2059 , po2060 , po2061 , po2062 , po2063 , po2064 , po2065 , po2066 , po2067 , po2068 , po2069 , po2070 , po2071 , po2072 , po2073 , po2074 , po2075 , po2076 , po2077 , po2078 , po2079 , po2080 , po2081 , po2082 , po2083 , po2084 , po2085 , po2086 , po2087 , po2088 , po2089 , po2090 , po2091 , po2092 , po2093 , po2094 , po2095 , po2096 , po2097 , po2098 , po2099 , po2100 , po2101 , po2102 , po2103 , po2104 , po2105 , po2106 , po2107 , po2108 , po2109 , po2110 , po2111 , po2112 , po2113 , po2114 , po2115 , po2116 , po2117 , po2118 , po2119 , po2120 , po2121 , po2122 , po2123 , po2124 , po2125 , po2126 , po2127 , po2128 , po2129 , po2130 , po2131 , po2132 , po2133 , po2134 , po2135 , po2136 , po2137 , po2138 , po2139 , po2140 , po2141 , po2142 , po2143 , po2144 , po2145 , po2146 , po2147 , po2148 , po2149 , po2150 , po2151 , po2152 , po2153 , po2154 , po2155 , po2156 , po2157 , po2158 , po2159 , po2160 , po2161 , po2162 , po2163 , po2164 , po2165 , po2166 , po2167 , po2168 , po2169 , po2170 , po2171 , po2172 , po2173 , po2174 , po2175 , po2176 , po2177 , po2178 , po2179 , po2180 , po2181 , po2182 , po2183 , po2184 , po2185 , po2186 , po2187 , po2188 , po2189 , po2190 , po2191 , po2192 , po2193 , po2194 , po2195 , po2196 , po2197 , po2198 , po2199 , po2200 , po2201 , po2202 , po2203 , po2204 , po2205 , po2206 , po2207 , po2208 , po2209 , po2210 , po2211 , po2212 , po2213 , po2214 , po2215 , po2216 , po2217 , po2218 , po2219 , po2220 , po2221 , po2222 , po2223 , po2224 , po2225 , po2226 , po2227 , po2228 , po2229 , po2230 , po2231 , po2232 , po2233 , po2234 , po2235 , po2236 , po2237 , po2238 , po2239 , po2240 , po2241 , po2242 , po2243 , po2244 , po2245 , po2246 , po2247 , po2248 , po2249 , po2250 , po2251 , po2252 , po2253 , po2254 , po2255 , po2256 , po2257 , po2258 , po2259 , po2260 , po2261 , po2262 , po2263 , po2264 , po2265 , po2266 , po2267 , po2268 , po2269 , po2270 , po2271 , po2272 , po2273 , po2274 , po2275 , po2276 , po2277 , po2278 , po2279 , po2280 , po2281 , po2282 , po2283 , po2284 , po2285 , po2286 , po2287 , po2288 , po2289 , po2290 , po2291 , po2292 , po2293 , po2294 , po2295 , po2296 , po2297 , po2298 , po2299 , po2300 , po2301 , po2302 , po2303 , po2304 , po2305 , po2306 , po2307 , po2308 , po2309 , po2310 , po2311 , po2312 , po2313 , po2314 , po2315 , po2316 , po2317 , po2318 , po2319 , po2320 , po2321 , po2322 , po2323 , po2324 , po2325 , po2326 , po2327 , po2328 , po2329 , po2330 , po2331 , po2332 , po2333 , po2334 , po2335 , po2336 , po2337 , po2338 , po2339 , po2340 , po2341 , po2342 , po2343 , po2344 , po2345 , po2346 , po2347 , po2348 , po2349 , po2350 , po2351 , po2352 , po2353 , po2354 , po2355 , po2356 , po2357 , po2358 , po2359 , po2360 , po2361 , po2362 , po2363 , po2364 , po2365 , po2366 , po2367 , po2368 , po2369 , po2370 , po2371 , po2372 , po2373 , po2374 , po2375 , po2376 , po2377 , po2378 , po2379 , po2380 , po2381 , po2382 , po2383 , po2384 , po2385 , po2386 , po2387 , po2388 , po2389 , po2390 , po2391 , po2392 , po2393 , po2394 , po2395 , po2396 , po2397 , po2398 , po2399 , po2400 , po2401 , po2402 , po2403 , po2404 , po2405 , po2406 , po2407 , po2408 , po2409 , po2410 , po2411 , po2412 , po2413 , po2414 , po2415 , po2416 , po2417 , po2418 , po2419 , po2420 , po2421 , po2422 , po2423 , po2424 , po2425 , po2426 , po2427 , po2428 , po2429 , po2430 , po2431 , po2432 , po2433 , po2434 , po2435 , po2436 , po2437 , po2438 , po2439 , po2440 , po2441 , po2442 , po2443 , po2444 , po2445 , po2446 , po2447 , po2448 , po2449 , po2450 , po2451 , po2452 , po2453 , po2454 , po2455 , po2456 , po2457 , po2458 , po2459 , po2460 , po2461 , po2462 , po2463 , po2464 , po2465 , po2466 , po2467 , po2468 , po2469 , po2470 , po2471 , po2472 , po2473 , po2474 , po2475 , po2476 , po2477 , po2478 , po2479 , po2480 , po2481 , po2482 , po2483 , po2484 , po2485 , po2486 , po2487 , po2488 , po2489 , po2490 , po2491 , po2492 , po2493 , po2494 , po2495 , po2496 , po2497 , po2498 , po2499 , po2500 , po2501 , po2502 , po2503 , po2504 , po2505 , po2506 , po2507 , po2508 , po2509 , po2510 , po2511 , po2512 , po2513 , po2514 , po2515 , po2516 , po2517 , po2518 , po2519 , po2520 , po2521 , po2522 , po2523 , po2524 , po2525 , po2526 , po2527 , po2528 , po2529 , po2530 , po2531 , po2532 , po2533 , po2534 , po2535 , po2536 , po2537 , po2538 , po2539 , po2540 , po2541 , po2542 , po2543 , po2544 , po2545 , po2546 , po2547 , po2548 , po2549 , po2550 , po2551 , po2552 , po2553 , po2554 , po2555 , po2556 , po2557 , po2558 , po2559 , po2560 , po2561 , po2562 , po2563 , po2564 , po2565 , po2566 , po2567 , po2568 , po2569 , po2570 , po2571 , po2572 , po2573 , po2574 , po2575 , po2576 , po2577 , po2578 , po2579 , po2580 , po2581 , po2582 , po2583 , po2584 , po2585 , po2586 , po2587 , po2588 , po2589 , po2590 , po2591 , po2592 , po2593 , po2594 , po2595 , po2596 , po2597 , po2598 , po2599 , po2600 , po2601 , po2602 , po2603 , po2604 , po2605 , po2606 , po2607 , po2608 , po2609 , po2610 , po2611 , po2612 , po2613 , po2614 , po2615 , po2616 , po2617 , po2618 , po2619 , po2620 , po2621 , po2622 , po2623 , po2624 , po2625 , po2626 , po2627 , po2628 , po2629 , po2630 , po2631 , po2632 , po2633 , po2634 , po2635 , po2636 , po2637 , po2638 , po2639 , po2640 , po2641 , po2642 , po2643 , po2644 , po2645 , po2646 , po2647 , po2648 , po2649 , po2650 , po2651 , po2652 , po2653 , po2654 , po2655 , po2656 , po2657 , po2658 , po2659 , po2660 , po2661 , po2662 , po2663 , po2664 , po2665 , po2666 , po2667 , po2668 , po2669 , po2670 , po2671 , po2672 , po2673 , po2674 , po2675 , po2676 , po2677 , po2678 , po2679 , po2680 , po2681 , po2682 , po2683 , po2684 , po2685 , po2686 , po2687 , po2688 , po2689 , po2690 , po2691 , po2692 , po2693 , po2694 , po2695 , po2696 , po2697 , po2698 , po2699 , po2700 , po2701 , po2702 , po2703 , po2704 , po2705 , po2706 , po2707 , po2708 , po2709 , po2710 , po2711 , po2712 , po2713 , po2714 , po2715 , po2716 , po2717 , po2718 , po2719 , po2720 , po2721 , po2722 , po2723 , po2724 , po2725 , po2726 , po2727 , po2728 , po2729 , po2730 , po2731 , po2732 , po2733 , po2734 , po2735 , po2736 , po2737 , po2738 , po2739 , po2740 , po2741 , po2742 , po2743 , po2744 , po2745 , po2746 , po2747 , po2748 , po2749 , po2750 , po2751 , po2752 , po2753 , po2754 , po2755 , po2756 , po2757 , po2758 , po2759 , po2760 , po2761 , po2762 , po2763 , po2764 , po2765 , po2766 , po2767 , po2768 , po2769 , po2770 , po2771 , po2772 , po2773 , po2774 , po2775 , po2776 , po2777 , po2778 , po2779 , po2780 , po2781 , po2782 , po2783 , po2784 , po2785 , po2786 , po2787 , po2788 , po2789 , po2790 , po2791 , po2792 , po2793 , po2794 , po2795 , po2796 , po2797 , po2798 , po2799 , po2800 , po2801 , po2802 , po2803 , po2804 , po2805 , po2806 , po2807 , po2808 , po2809 , po2810 , po2811 , po2812 , po2813 , po2814 , po2815 , po2816 , po2817 , po2818 , po2819 , po2820 , po2821 , po2822 , po2823 , po2824 , po2825 , po2826 , po2827 , po2828 , po2829 , po2830 , po2831 , po2832 , po2833 , po2834 , po2835 , po2836 , po2837 , po2838 , po2839 , po2840 , po2841 , po2842 , po2843 , po2844 , po2845 , po2846 , po2847 , po2848 , po2849 , po2850 , po2851 , po2852 , po2853 , po2854 , po2855 , po2856 , po2857 , po2858 , po2859 , po2860 , po2861 , po2862 , po2863 , po2864 , po2865 , po2866 , po2867 , po2868 , po2869 , po2870 , po2871 , po2872 , po2873 , po2874 , po2875 , po2876 , po2877 , po2878 , po2879 , po2880 , po2881 , po2882 , po2883 , po2884 , po2885 , po2886 , po2887 , po2888 , po2889 , po2890 , po2891 , po2892 , po2893 , po2894 , po2895 , po2896 , po2897 , po2898 , po2899 , po2900 , po2901 , po2902 , po2903 , po2904 , po2905 , po2906 , po2907 , po2908 , po2909 , po2910 , po2911 , po2912 , po2913 , po2914 , po2915 , po2916 , po2917 , po2918 , po2919 , po2920 , po2921 , po2922 , po2923 , po2924 , po2925 , po2926 , po2927 , po2928 , po2929 , po2930 , po2931 , po2932 , po2933 , po2934 , po2935 , po2936 , po2937 , po2938 , po2939 , po2940 , po2941 , po2942 , po2943 , po2944 , po2945 , po2946 , po2947 , po2948 , po2949 , po2950 , po2951 , po2952 , po2953 , po2954 , po2955 , po2956 , po2957 , po2958 , po2959 , po2960 , po2961 , po2962 , po2963 , po2964 , po2965 , po2966 , po2967 , po2968 , po2969 , po2970 , po2971 , po2972 , po2973 , po2974 , po2975 , po2976 , po2977 , po2978 , po2979 , po2980 , po2981 , po2982 , po2983 , po2984 , po2985 , po2986 , po2987 , po2988 , po2989 , po2990 , po2991 , po2992 , po2993 , po2994 , po2995 , po2996 , po2997 , po2998 , po2999 , po3000 , po3001 , po3002 , po3003 , po3004 , po3005 , po3006 , po3007 , po3008 , po3009 , po3010 , po3011 , po3012 , po3013 , po3014 , po3015 , po3016 , po3017 , po3018 , po3019 , po3020 , po3021 , po3022 , po3023 , po3024 , po3025 , po3026 , po3027 , po3028 , po3029 , po3030 , po3031 , po3032 , po3033 , po3034 , po3035 , po3036 , po3037 , po3038 , po3039 , po3040 , po3041 , po3042 , po3043 , po3044 , po3045 , po3046 , po3047 , po3048 , po3049 , po3050 , po3051 , po3052 , po3053 , po3054 , po3055 , po3056 , po3057 , po3058 , po3059 , po3060 , po3061 , po3062 , po3063 , po3064 , po3065 , po3066 , po3067 , po3068 , po3069 , po3070 , po3071 , po3072 , po3073 , po3074 , po3075 , po3076 , po3077 , po3078 , po3079 , po3080 , po3081 , po3082 , po3083 , po3084 , po3085 , po3086 , po3087 , po3088 , po3089 , po3090 , po3091 , po3092 , po3093 , po3094 , po3095 , po3096 , po3097 , po3098 , po3099 , po3100 , po3101 , po3102 , po3103 , po3104 , po3105 , po3106 , po3107 , po3108 , po3109 , po3110 , po3111 , po3112 , po3113 , po3114 , po3115 , po3116 , po3117 , po3118 , po3119 , po3120 , po3121 , po3122 , po3123 , po3124 , po3125 , po3126 , po3127 , po3128 , po3129 , po3130 , po3131 , po3132 , po3133 , po3134 , po3135 , po3136 , po3137 , po3138 , po3139 , po3140 , po3141 , po3142 , po3143 , po3144 , po3145 , po3146 , po3147 , po3148 , po3149 , po3150 , po3151 , po3152 , po3153 , po3154 , po3155 , po3156 , po3157 , po3158 , po3159 , po3160 , po3161 , po3162 , po3163 , po3164 , po3165 , po3166 , po3167 , po3168 , po3169 , po3170 , po3171 , po3172 , po3173 , po3174 , po3175 , po3176 , po3177 , po3178 , po3179 , po3180 , po3181 , po3182 , po3183 , po3184 , po3185 , po3186 , po3187 , po3188 , po3189 , po3190 , po3191 , po3192 , po3193 , po3194 , po3195 , po3196 , po3197 , po3198 , po3199 , po3200 , po3201 , po3202 , po3203 , po3204 , po3205 , po3206 , po3207 , po3208 , po3209 , po3210 , po3211 , po3212 , po3213 , po3214 , po3215 , po3216 , po3217 , po3218 , po3219 , po3220 , po3221 , po3222 , po3223 , po3224 , po3225 , po3226 , po3227 , po3228 , po3229 , po3230 , po3231 , po3232 , po3233 , po3234 , po3235 , po3236 , po3237 , po3238 , po3239 , po3240 , po3241 , po3242 , po3243 , po3244 , po3245 , po3246 , po3247 , po3248 , po3249 , po3250 , po3251 , po3252 , po3253 , po3254 , po3255 , po3256 , po3257 , po3258 , po3259 , po3260 , po3261 , po3262 , po3263 , po3264 , po3265 , po3266 , po3267 , po3268 , po3269 , po3270 , po3271 , po3272 , po3273 , po3274 , po3275 , po3276 , po3277 , po3278 , po3279 , po3280 , po3281 , po3282 , po3283 , po3284 , po3285 , po3286 , po3287 , po3288 , po3289 , po3290 , po3291 , po3292 , po3293 , po3294 , po3295 , po3296 , po3297 , po3298 , po3299 , po3300 , po3301 , po3302 , po3303 , po3304 , po3305 , po3306 , po3307 , po3308 , po3309 , po3310 , po3311 , po3312 , po3313 , po3314 , po3315 , po3316 , po3317 , po3318 , po3319 , po3320 , po3321 , po3322 , po3323 , po3324 , po3325 , po3326 , po3327 );
  input pi000 , pi001 , pi002 , pi003 , pi004 , pi005 , pi006 , pi007 , pi008 , pi009 , pi010 , pi011 , pi012 , pi013 , pi014 , pi015 , pi016 , pi017 , pi018 , pi019 , pi020 , pi021 , pi022 , pi023 , pi024 , pi025 , pi026 , pi027 , pi028 , pi029 , pi030 , pi031 , pi032 , pi033 , pi034 , pi035 , pi036 , pi037 , pi038 , pi039 , pi040 , pi041 , pi042 , pi043 , pi044 , pi045 , pi046 , pi047 , pi048 , pi049 , pi050 , pi051 , pi052 , pi053 , pi054 , pi055 , pi056 , pi057 , pi058 , pi059 , pi060 , pi061 , pi062 , pi063 , pi064 , pi065 , pi066 , pi067 , pi068 , pi069 , pi070 , pi071 , pi072 , pi073 , pi074 , pi075 , pi076 , pi077 , pi078 , pi079 , pi080 , pi081 , pi082 , pi083 , pi084 , pi085 , pi086 , pi087 , pi088 , pi089 , pi090 , pi091 , pi092 , pi093 , pi094 , pi095 , pi096 , pi097 , pi098 , pi099 , pi100 , pi101 , pi102 , pi103 , pi104 , pi105 , pi106 , pi107 , pi108 , pi109 , pi110 , pi111 , pi112 , pi113 , pi114 , pi115 , pi116 , pi117 , pi118 , pi119 , pi120 , pi121 , pi122 , pi123 , pi124 , pi125 , pi126 , pi127 , pi128 , pi129 , pi130 , pi131 , pi132 , pi133 , pi134 , pi135 , pi136 , pi137 , pi138 , pi139 , pi140 , pi141 , pi142 , pi143 , pi144 , pi145 , pi146 , pi147 , pi148 , pi149 , pi150 , pi151 , pi152 , pi153 , pi154 , pi155 , pi156 , pi157 , pi158 , pi159 , pi160 , pi161 , pi162 , pi163 , pi164 , pi165 , pi166 , pi167 , pi168 , pi169 , pi170 , pi171 , pi172 , pi173 , pi174 , pi175 , pi176 , pi177 , pi178 , pi179 , pi180 , pi181 , pi182 , pi183 , pi184 , pi185 , pi186 , pi187 , pi188 , pi189 , pi190 , pi191 , pi192 , pi193 , pi194 , pi195 , pi196 , pi197 , pi198 , pi199 , pi200 , pi201 , pi202 , pi203 , pi204 , pi205 , pi206 , pi207 , pi208 , pi209 , pi210 , pi211 , pi212 , pi213 , pi214 , pi215 , pi216 , pi217 , pi218 , pi219 , pi220 , pi221 , pi222 , pi223 , pi224 , pi225 , pi226 , pi227 , pi228 , pi229 , pi230 , pi231 , pi232 , pi233 , pi234 , pi235 , pi236 , pi237 , pi238 , pi239 , pi240 , pi241 , pi242 , pi243 , pi244 , pi245 , pi246 , pi247 , pi248 , pi249 , pi250 , pi251 , pi252 , pi253 , pi254 , pi255 , pi256 , pi257 , pi258 , pi259 , pi260 , pi261 , pi262 , pi263 , pi264 , pi265 , pi266 , pi267 , pi268 , pi269 , pi270 , pi271 , pi272 , pi273 , pi274 , pi275 , pi276 , pi277 , pi278 , pi279 , pi280 , pi281 , pi282 , pi283 , pi284 , pi285 , pi286 , pi287 , pi288 , pi289 , pi290 , pi291 , pi292 , pi293 , pi294 , pi295 , pi296 , pi297 , pi298 , pi299 , pi300 , pi301 , pi302 , pi303 , pi304 , pi305 , pi306 , pi307 , pi308 , pi309 , pi310 , pi311 , pi312 , pi313 , pi314 , pi315 , pi316 , pi317 , pi318 , pi319 , pi320 , pi321 , pi322 , pi323 , pi324 , pi325 , pi326 , pi327 , pi328 , pi329 , pi330 , pi331 , pi332 , pi333 , pi334 , pi335 , pi336 , pi337 , pi338 , pi339 , pi340 , pi341 , pi342 , pi343 , pi344 , pi345 , pi346 , pi347 , pi348 , pi349 , pi350 , pi351 , pi352 , pi353 , pi354 , pi355 , pi356 , pi357 , pi358 , pi359 , pi360 , pi361 , pi362 , pi363 , pi364 , pi365 , pi366 , pi367 , pi368 , pi369 , pi370 , pi371 , pi372 , pi373 , pi374 , pi375 , pi376 , pi377 , pi378 , pi379 , pi380 , pi381 , pi382 , pi383 , pi384 , pi385 , pi386 , pi387 , pi388 , pi389 , pi390 , pi391 , pi392 , pi393 , pi394 , pi395 , pi396 , pi397 , pi398 , pi399 , pi400 , pi401 , pi402 , pi403 , pi404 , pi405 , pi406 , pi407 , pi408 , pi409 , pi410 , pi411 , pi412 , pi413 , pi414 , pi415 , pi416 , pi417 , pi418 , pi419 , pi420 , pi421 , pi422 , pi423 , pi424 , pi425 , pi426 , pi427 , pi428 , pi429 , pi430 , pi431 , pi432 , pi433 , pi434 , pi435 , pi436 , pi437 , pi438 , pi439 , pi440 , pi441 , pi442 , pi443 , pi444 , pi445 , pi446 , pi447 , pi448 , pi449 , pi450 , pi451 , pi452 , pi453 , pi454 , pi455 , pi456 , pi457 , pi458 , pi459 , pi460 , pi461 , pi462 , pi463 ;
  output po0000 , po0001 , po0002 , po0003 , po0004 , po0005 , po0006 , po0007 , po0008 , po0009 , po0010 , po0011 , po0012 , po0013 , po0014 , po0015 , po0016 , po0017 , po0018 , po0019 , po0020 , po0021 , po0022 , po0023 , po0024 , po0025 , po0026 , po0027 , po0028 , po0029 , po0030 , po0031 , po0032 , po0033 , po0034 , po0035 , po0036 , po0037 , po0038 , po0039 , po0040 , po0041 , po0042 , po0043 , po0044 , po0045 , po0046 , po0047 , po0048 , po0049 , po0050 , po0051 , po0052 , po0053 , po0054 , po0055 , po0056 , po0057 , po0058 , po0059 , po0060 , po0061 , po0062 , po0063 , po0064 , po0065 , po0066 , po0067 , po0068 , po0069 , po0070 , po0071 , po0072 , po0073 , po0074 , po0075 , po0076 , po0077 , po0078 , po0079 , po0080 , po0081 , po0082 , po0083 , po0084 , po0085 , po0086 , po0087 , po0088 , po0089 , po0090 , po0091 , po0092 , po0093 , po0094 , po0095 , po0096 , po0097 , po0098 , po0099 , po0100 , po0101 , po0102 , po0103 , po0104 , po0105 , po0106 , po0107 , po0108 , po0109 , po0110 , po0111 , po0112 , po0113 , po0114 , po0115 , po0116 , po0117 , po0118 , po0119 , po0120 , po0121 , po0122 , po0123 , po0124 , po0125 , po0126 , po0127 , po0128 , po0129 , po0130 , po0131 , po0132 , po0133 , po0134 , po0135 , po0136 , po0137 , po0138 , po0139 , po0140 , po0141 , po0142 , po0143 , po0144 , po0145 , po0146 , po0147 , po0148 , po0149 , po0150 , po0151 , po0152 , po0153 , po0154 , po0155 , po0156 , po0157 , po0158 , po0159 , po0160 , po0161 , po0162 , po0163 , po0164 , po0165 , po0166 , po0167 , po0168 , po0169 , po0170 , po0171 , po0172 , po0173 , po0174 , po0175 , po0176 , po0177 , po0178 , po0179 , po0180 , po0181 , po0182 , po0183 , po0184 , po0185 , po0186 , po0187 , po0188 , po0189 , po0190 , po0191 , po0192 , po0193 , po0194 , po0195 , po0196 , po0197 , po0198 , po0199 , po0200 , po0201 , po0202 , po0203 , po0204 , po0205 , po0206 , po0207 , po0208 , po0209 , po0210 , po0211 , po0212 , po0213 , po0214 , po0215 , po0216 , po0217 , po0218 , po0219 , po0220 , po0221 , po0222 , po0223 , po0224 , po0225 , po0226 , po0227 , po0228 , po0229 , po0230 , po0231 , po0232 , po0233 , po0234 , po0235 , po0236 , po0237 , po0238 , po0239 , po0240 , po0241 , po0242 , po0243 , po0244 , po0245 , po0246 , po0247 , po0248 , po0249 , po0250 , po0251 , po0252 , po0253 , po0254 , po0255 , po0256 , po0257 , po0258 , po0259 , po0260 , po0261 , po0262 , po0263 , po0264 , po0265 , po0266 , po0267 , po0268 , po0269 , po0270 , po0271 , po0272 , po0273 , po0274 , po0275 , po0276 , po0277 , po0278 , po0279 , po0280 , po0281 , po0282 , po0283 , po0284 , po0285 , po0286 , po0287 , po0288 , po0289 , po0290 , po0291 , po0292 , po0293 , po0294 , po0295 , po0296 , po0297 , po0298 , po0299 , po0300 , po0301 , po0302 , po0303 , po0304 , po0305 , po0306 , po0307 , po0308 , po0309 , po0310 , po0311 , po0312 , po0313 , po0314 , po0315 , po0316 , po0317 , po0318 , po0319 , po0320 , po0321 , po0322 , po0323 , po0324 , po0325 , po0326 , po0327 , po0328 , po0329 , po0330 , po0331 , po0332 , po0333 , po0334 , po0335 , po0336 , po0337 , po0338 , po0339 , po0340 , po0341 , po0342 , po0343 , po0344 , po0345 , po0346 , po0347 , po0348 , po0349 , po0350 , po0351 , po0352 , po0353 , po0354 , po0355 , po0356 , po0357 , po0358 , po0359 , po0360 , po0361 , po0362 , po0363 , po0364 , po0365 , po0366 , po0367 , po0368 , po0369 , po0370 , po0371 , po0372 , po0373 , po0374 , po0375 , po0376 , po0377 , po0378 , po0379 , po0380 , po0381 , po0382 , po0383 , po0384 , po0385 , po0386 , po0387 , po0388 , po0389 , po0390 , po0391 , po0392 , po0393 , po0394 , po0395 , po0396 , po0397 , po0398 , po0399 , po0400 , po0401 , po0402 , po0403 , po0404 , po0405 , po0406 , po0407 , po0408 , po0409 , po0410 , po0411 , po0412 , po0413 , po0414 , po0415 , po0416 , po0417 , po0418 , po0419 , po0420 , po0421 , po0422 , po0423 , po0424 , po0425 , po0426 , po0427 , po0428 , po0429 , po0430 , po0431 , po0432 , po0433 , po0434 , po0435 , po0436 , po0437 , po0438 , po0439 , po0440 , po0441 , po0442 , po0443 , po0444 , po0445 , po0446 , po0447 , po0448 , po0449 , po0450 , po0451 , po0452 , po0453 , po0454 , po0455 , po0456 , po0457 , po0458 , po0459 , po0460 , po0461 , po0462 , po0463 , po0464 , po0465 , po0466 , po0467 , po0468 , po0469 , po0470 , po0471 , po0472 , po0473 , po0474 , po0475 , po0476 , po0477 , po0478 , po0479 , po0480 , po0481 , po0482 , po0483 , po0484 , po0485 , po0486 , po0487 , po0488 , po0489 , po0490 , po0491 , po0492 , po0493 , po0494 , po0495 , po0496 , po0497 , po0498 , po0499 , po0500 , po0501 , po0502 , po0503 , po0504 , po0505 , po0506 , po0507 , po0508 , po0509 , po0510 , po0511 , po0512 , po0513 , po0514 , po0515 , po0516 , po0517 , po0518 , po0519 , po0520 , po0521 , po0522 , po0523 , po0524 , po0525 , po0526 , po0527 , po0528 , po0529 , po0530 , po0531 , po0532 , po0533 , po0534 , po0535 , po0536 , po0537 , po0538 , po0539 , po0540 , po0541 , po0542 , po0543 , po0544 , po0545 , po0546 , po0547 , po0548 , po0549 , po0550 , po0551 , po0552 , po0553 , po0554 , po0555 , po0556 , po0557 , po0558 , po0559 , po0560 , po0561 , po0562 , po0563 , po0564 , po0565 , po0566 , po0567 , po0568 , po0569 , po0570 , po0571 , po0572 , po0573 , po0574 , po0575 , po0576 , po0577 , po0578 , po0579 , po0580 , po0581 , po0582 , po0583 , po0584 , po0585 , po0586 , po0587 , po0588 , po0589 , po0590 , po0591 , po0592 , po0593 , po0594 , po0595 , po0596 , po0597 , po0598 , po0599 , po0600 , po0601 , po0602 , po0603 , po0604 , po0605 , po0606 , po0607 , po0608 , po0609 , po0610 , po0611 , po0612 , po0613 , po0614 , po0615 , po0616 , po0617 , po0618 , po0619 , po0620 , po0621 , po0622 , po0623 , po0624 , po0625 , po0626 , po0627 , po0628 , po0629 , po0630 , po0631 , po0632 , po0633 , po0634 , po0635 , po0636 , po0637 , po0638 , po0639 , po0640 , po0641 , po0642 , po0643 , po0644 , po0645 , po0646 , po0647 , po0648 , po0649 , po0650 , po0651 , po0652 , po0653 , po0654 , po0655 , po0656 , po0657 , po0658 , po0659 , po0660 , po0661 , po0662 , po0663 , po0664 , po0665 , po0666 , po0667 , po0668 , po0669 , po0670 , po0671 , po0672 , po0673 , po0674 , po0675 , po0676 , po0677 , po0678 , po0679 , po0680 , po0681 , po0682 , po0683 , po0684 , po0685 , po0686 , po0687 , po0688 , po0689 , po0690 , po0691 , po0692 , po0693 , po0694 , po0695 , po0696 , po0697 , po0698 , po0699 , po0700 , po0701 , po0702 , po0703 , po0704 , po0705 , po0706 , po0707 , po0708 , po0709 , po0710 , po0711 , po0712 , po0713 , po0714 , po0715 , po0716 , po0717 , po0718 , po0719 , po0720 , po0721 , po0722 , po0723 , po0724 , po0725 , po0726 , po0727 , po0728 , po0729 , po0730 , po0731 , po0732 , po0733 , po0734 , po0735 , po0736 , po0737 , po0738 , po0739 , po0740 , po0741 , po0742 , po0743 , po0744 , po0745 , po0746 , po0747 , po0748 , po0749 , po0750 , po0751 , po0752 , po0753 , po0754 , po0755 , po0756 , po0757 , po0758 , po0759 , po0760 , po0761 , po0762 , po0763 , po0764 , po0765 , po0766 , po0767 , po0768 , po0769 , po0770 , po0771 , po0772 , po0773 , po0774 , po0775 , po0776 , po0777 , po0778 , po0779 , po0780 , po0781 , po0782 , po0783 , po0784 , po0785 , po0786 , po0787 , po0788 , po0789 , po0790 , po0791 , po0792 , po0793 , po0794 , po0795 , po0796 , po0797 , po0798 , po0799 , po0800 , po0801 , po0802 , po0803 , po0804 , po0805 , po0806 , po0807 , po0808 , po0809 , po0810 , po0811 , po0812 , po0813 , po0814 , po0815 , po0816 , po0817 , po0818 , po0819 , po0820 , po0821 , po0822 , po0823 , po0824 , po0825 , po0826 , po0827 , po0828 , po0829 , po0830 , po0831 , po0832 , po0833 , po0834 , po0835 , po0836 , po0837 , po0838 , po0839 , po0840 , po0841 , po0842 , po0843 , po0844 , po0845 , po0846 , po0847 , po0848 , po0849 , po0850 , po0851 , po0852 , po0853 , po0854 , po0855 , po0856 , po0857 , po0858 , po0859 , po0860 , po0861 , po0862 , po0863 , po0864 , po0865 , po0866 , po0867 , po0868 , po0869 , po0870 , po0871 , po0872 , po0873 , po0874 , po0875 , po0876 , po0877 , po0878 , po0879 , po0880 , po0881 , po0882 , po0883 , po0884 , po0885 , po0886 , po0887 , po0888 , po0889 , po0890 , po0891 , po0892 , po0893 , po0894 , po0895 , po0896 , po0897 , po0898 , po0899 , po0900 , po0901 , po0902 , po0903 , po0904 , po0905 , po0906 , po0907 , po0908 , po0909 , po0910 , po0911 , po0912 , po0913 , po0914 , po0915 , po0916 , po0917 , po0918 , po0919 , po0920 , po0921 , po0922 , po0923 , po0924 , po0925 , po0926 , po0927 , po0928 , po0929 , po0930 , po0931 , po0932 , po0933 , po0934 , po0935 , po0936 , po0937 , po0938 , po0939 , po0940 , po0941 , po0942 , po0943 , po0944 , po0945 , po0946 , po0947 , po0948 , po0949 , po0950 , po0951 , po0952 , po0953 , po0954 , po0955 , po0956 , po0957 , po0958 , po0959 , po0960 , po0961 , po0962 , po0963 , po0964 , po0965 , po0966 , po0967 , po0968 , po0969 , po0970 , po0971 , po0972 , po0973 , po0974 , po0975 , po0976 , po0977 , po0978 , po0979 , po0980 , po0981 , po0982 , po0983 , po0984 , po0985 , po0986 , po0987 , po0988 , po0989 , po0990 , po0991 , po0992 , po0993 , po0994 , po0995 , po0996 , po0997 , po0998 , po0999 , po1000 , po1001 , po1002 , po1003 , po1004 , po1005 , po1006 , po1007 , po1008 , po1009 , po1010 , po1011 , po1012 , po1013 , po1014 , po1015 , po1016 , po1017 , po1018 , po1019 , po1020 , po1021 , po1022 , po1023 , po1024 , po1025 , po1026 , po1027 , po1028 , po1029 , po1030 , po1031 , po1032 , po1033 , po1034 , po1035 , po1036 , po1037 , po1038 , po1039 , po1040 , po1041 , po1042 , po1043 , po1044 , po1045 , po1046 , po1047 , po1048 , po1049 , po1050 , po1051 , po1052 , po1053 , po1054 , po1055 , po1056 , po1057 , po1058 , po1059 , po1060 , po1061 , po1062 , po1063 , po1064 , po1065 , po1066 , po1067 , po1068 , po1069 , po1070 , po1071 , po1072 , po1073 , po1074 , po1075 , po1076 , po1077 , po1078 , po1079 , po1080 , po1081 , po1082 , po1083 , po1084 , po1085 , po1086 , po1087 , po1088 , po1089 , po1090 , po1091 , po1092 , po1093 , po1094 , po1095 , po1096 , po1097 , po1098 , po1099 , po1100 , po1101 , po1102 , po1103 , po1104 , po1105 , po1106 , po1107 , po1108 , po1109 , po1110 , po1111 , po1112 , po1113 , po1114 , po1115 , po1116 , po1117 , po1118 , po1119 , po1120 , po1121 , po1122 , po1123 , po1124 , po1125 , po1126 , po1127 , po1128 , po1129 , po1130 , po1131 , po1132 , po1133 , po1134 , po1135 , po1136 , po1137 , po1138 , po1139 , po1140 , po1141 , po1142 , po1143 , po1144 , po1145 , po1146 , po1147 , po1148 , po1149 , po1150 , po1151 , po1152 , po1153 , po1154 , po1155 , po1156 , po1157 , po1158 , po1159 , po1160 , po1161 , po1162 , po1163 , po1164 , po1165 , po1166 , po1167 , po1168 , po1169 , po1170 , po1171 , po1172 , po1173 , po1174 , po1175 , po1176 , po1177 , po1178 , po1179 , po1180 , po1181 , po1182 , po1183 , po1184 , po1185 , po1186 , po1187 , po1188 , po1189 , po1190 , po1191 , po1192 , po1193 , po1194 , po1195 , po1196 , po1197 , po1198 , po1199 , po1200 , po1201 , po1202 , po1203 , po1204 , po1205 , po1206 , po1207 , po1208 , po1209 , po1210 , po1211 , po1212 , po1213 , po1214 , po1215 , po1216 , po1217 , po1218 , po1219 , po1220 , po1221 , po1222 , po1223 , po1224 , po1225 , po1226 , po1227 , po1228 , po1229 , po1230 , po1231 , po1232 , po1233 , po1234 , po1235 , po1236 , po1237 , po1238 , po1239 , po1240 , po1241 , po1242 , po1243 , po1244 , po1245 , po1246 , po1247 , po1248 , po1249 , po1250 , po1251 , po1252 , po1253 , po1254 , po1255 , po1256 , po1257 , po1258 , po1259 , po1260 , po1261 , po1262 , po1263 , po1264 , po1265 , po1266 , po1267 , po1268 , po1269 , po1270 , po1271 , po1272 , po1273 , po1274 , po1275 , po1276 , po1277 , po1278 , po1279 , po1280 , po1281 , po1282 , po1283 , po1284 , po1285 , po1286 , po1287 , po1288 , po1289 , po1290 , po1291 , po1292 , po1293 , po1294 , po1295 , po1296 , po1297 , po1298 , po1299 , po1300 , po1301 , po1302 , po1303 , po1304 , po1305 , po1306 , po1307 , po1308 , po1309 , po1310 , po1311 , po1312 , po1313 , po1314 , po1315 , po1316 , po1317 , po1318 , po1319 , po1320 , po1321 , po1322 , po1323 , po1324 , po1325 , po1326 , po1327 , po1328 , po1329 , po1330 , po1331 , po1332 , po1333 , po1334 , po1335 , po1336 , po1337 , po1338 , po1339 , po1340 , po1341 , po1342 , po1343 , po1344 , po1345 , po1346 , po1347 , po1348 , po1349 , po1350 , po1351 , po1352 , po1353 , po1354 , po1355 , po1356 , po1357 , po1358 , po1359 , po1360 , po1361 , po1362 , po1363 , po1364 , po1365 , po1366 , po1367 , po1368 , po1369 , po1370 , po1371 , po1372 , po1373 , po1374 , po1375 , po1376 , po1377 , po1378 , po1379 , po1380 , po1381 , po1382 , po1383 , po1384 , po1385 , po1386 , po1387 , po1388 , po1389 , po1390 , po1391 , po1392 , po1393 , po1394 , po1395 , po1396 , po1397 , po1398 , po1399 , po1400 , po1401 , po1402 , po1403 , po1404 , po1405 , po1406 , po1407 , po1408 , po1409 , po1410 , po1411 , po1412 , po1413 , po1414 , po1415 , po1416 , po1417 , po1418 , po1419 , po1420 , po1421 , po1422 , po1423 , po1424 , po1425 , po1426 , po1427 , po1428 , po1429 , po1430 , po1431 , po1432 , po1433 , po1434 , po1435 , po1436 , po1437 , po1438 , po1439 , po1440 , po1441 , po1442 , po1443 , po1444 , po1445 , po1446 , po1447 , po1448 , po1449 , po1450 , po1451 , po1452 , po1453 , po1454 , po1455 , po1456 , po1457 , po1458 , po1459 , po1460 , po1461 , po1462 , po1463 , po1464 , po1465 , po1466 , po1467 , po1468 , po1469 , po1470 , po1471 , po1472 , po1473 , po1474 , po1475 , po1476 , po1477 , po1478 , po1479 , po1480 , po1481 , po1482 , po1483 , po1484 , po1485 , po1486 , po1487 , po1488 , po1489 , po1490 , po1491 , po1492 , po1493 , po1494 , po1495 , po1496 , po1497 , po1498 , po1499 , po1500 , po1501 , po1502 , po1503 , po1504 , po1505 , po1506 , po1507 , po1508 , po1509 , po1510 , po1511 , po1512 , po1513 , po1514 , po1515 , po1516 , po1517 , po1518 , po1519 , po1520 , po1521 , po1522 , po1523 , po1524 , po1525 , po1526 , po1527 , po1528 , po1529 , po1530 , po1531 , po1532 , po1533 , po1534 , po1535 , po1536 , po1537 , po1538 , po1539 , po1540 , po1541 , po1542 , po1543 , po1544 , po1545 , po1546 , po1547 , po1548 , po1549 , po1550 , po1551 , po1552 , po1553 , po1554 , po1555 , po1556 , po1557 , po1558 , po1559 , po1560 , po1561 , po1562 , po1563 , po1564 , po1565 , po1566 , po1567 , po1568 , po1569 , po1570 , po1571 , po1572 , po1573 , po1574 , po1575 , po1576 , po1577 , po1578 , po1579 , po1580 , po1581 , po1582 , po1583 , po1584 , po1585 , po1586 , po1587 , po1588 , po1589 , po1590 , po1591 , po1592 , po1593 , po1594 , po1595 , po1596 , po1597 , po1598 , po1599 , po1600 , po1601 , po1602 , po1603 , po1604 , po1605 , po1606 , po1607 , po1608 , po1609 , po1610 , po1611 , po1612 , po1613 , po1614 , po1615 , po1616 , po1617 , po1618 , po1619 , po1620 , po1621 , po1622 , po1623 , po1624 , po1625 , po1626 , po1627 , po1628 , po1629 , po1630 , po1631 , po1632 , po1633 , po1634 , po1635 , po1636 , po1637 , po1638 , po1639 , po1640 , po1641 , po1642 , po1643 , po1644 , po1645 , po1646 , po1647 , po1648 , po1649 , po1650 , po1651 , po1652 , po1653 , po1654 , po1655 , po1656 , po1657 , po1658 , po1659 , po1660 , po1661 , po1662 , po1663 , po1664 , po1665 , po1666 , po1667 , po1668 , po1669 , po1670 , po1671 , po1672 , po1673 , po1674 , po1675 , po1676 , po1677 , po1678 , po1679 , po1680 , po1681 , po1682 , po1683 , po1684 , po1685 , po1686 , po1687 , po1688 , po1689 , po1690 , po1691 , po1692 , po1693 , po1694 , po1695 , po1696 , po1697 , po1698 , po1699 , po1700 , po1701 , po1702 , po1703 , po1704 , po1705 , po1706 , po1707 , po1708 , po1709 , po1710 , po1711 , po1712 , po1713 , po1714 , po1715 , po1716 , po1717 , po1718 , po1719 , po1720 , po1721 , po1722 , po1723 , po1724 , po1725 , po1726 , po1727 , po1728 , po1729 , po1730 , po1731 , po1732 , po1733 , po1734 , po1735 , po1736 , po1737 , po1738 , po1739 , po1740 , po1741 , po1742 , po1743 , po1744 , po1745 , po1746 , po1747 , po1748 , po1749 , po1750 , po1751 , po1752 , po1753 , po1754 , po1755 , po1756 , po1757 , po1758 , po1759 , po1760 , po1761 , po1762 , po1763 , po1764 , po1765 , po1766 , po1767 , po1768 , po1769 , po1770 , po1771 , po1772 , po1773 , po1774 , po1775 , po1776 , po1777 , po1778 , po1779 , po1780 , po1781 , po1782 , po1783 , po1784 , po1785 , po1786 , po1787 , po1788 , po1789 , po1790 , po1791 , po1792 , po1793 , po1794 , po1795 , po1796 , po1797 , po1798 , po1799 , po1800 , po1801 , po1802 , po1803 , po1804 , po1805 , po1806 , po1807 , po1808 , po1809 , po1810 , po1811 , po1812 , po1813 , po1814 , po1815 , po1816 , po1817 , po1818 , po1819 , po1820 , po1821 , po1822 , po1823 , po1824 , po1825 , po1826 , po1827 , po1828 , po1829 , po1830 , po1831 , po1832 , po1833 , po1834 , po1835 , po1836 , po1837 , po1838 , po1839 , po1840 , po1841 , po1842 , po1843 , po1844 , po1845 , po1846 , po1847 , po1848 , po1849 , po1850 , po1851 , po1852 , po1853 , po1854 , po1855 , po1856 , po1857 , po1858 , po1859 , po1860 , po1861 , po1862 , po1863 , po1864 , po1865 , po1866 , po1867 , po1868 , po1869 , po1870 , po1871 , po1872 , po1873 , po1874 , po1875 , po1876 , po1877 , po1878 , po1879 , po1880 , po1881 , po1882 , po1883 , po1884 , po1885 , po1886 , po1887 , po1888 , po1889 , po1890 , po1891 , po1892 , po1893 , po1894 , po1895 , po1896 , po1897 , po1898 , po1899 , po1900 , po1901 , po1902 , po1903 , po1904 , po1905 , po1906 , po1907 , po1908 , po1909 , po1910 , po1911 , po1912 , po1913 , po1914 , po1915 , po1916 , po1917 , po1918 , po1919 , po1920 , po1921 , po1922 , po1923 , po1924 , po1925 , po1926 , po1927 , po1928 , po1929 , po1930 , po1931 , po1932 , po1933 , po1934 , po1935 , po1936 , po1937 , po1938 , po1939 , po1940 , po1941 , po1942 , po1943 , po1944 , po1945 , po1946 , po1947 , po1948 , po1949 , po1950 , po1951 , po1952 , po1953 , po1954 , po1955 , po1956 , po1957 , po1958 , po1959 , po1960 , po1961 , po1962 , po1963 , po1964 , po1965 , po1966 , po1967 , po1968 , po1969 , po1970 , po1971 , po1972 , po1973 , po1974 , po1975 , po1976 , po1977 , po1978 , po1979 , po1980 , po1981 , po1982 , po1983 , po1984 , po1985 , po1986 , po1987 , po1988 , po1989 , po1990 , po1991 , po1992 , po1993 , po1994 , po1995 , po1996 , po1997 , po1998 , po1999 , po2000 , po2001 , po2002 , po2003 , po2004 , po2005 , po2006 , po2007 , po2008 , po2009 , po2010 , po2011 , po2012 , po2013 , po2014 , po2015 , po2016 , po2017 , po2018 , po2019 , po2020 , po2021 , po2022 , po2023 , po2024 , po2025 , po2026 , po2027 , po2028 , po2029 , po2030 , po2031 , po2032 , po2033 , po2034 , po2035 , po2036 , po2037 , po2038 , po2039 , po2040 , po2041 , po2042 , po2043 , po2044 , po2045 , po2046 , po2047 , po2048 , po2049 , po2050 , po2051 , po2052 , po2053 , po2054 , po2055 , po2056 , po2057 , po2058 , po2059 , po2060 , po2061 , po2062 , po2063 , po2064 , po2065 , po2066 , po2067 , po2068 , po2069 , po2070 , po2071 , po2072 , po2073 , po2074 , po2075 , po2076 , po2077 , po2078 , po2079 , po2080 , po2081 , po2082 , po2083 , po2084 , po2085 , po2086 , po2087 , po2088 , po2089 , po2090 , po2091 , po2092 , po2093 , po2094 , po2095 , po2096 , po2097 , po2098 , po2099 , po2100 , po2101 , po2102 , po2103 , po2104 , po2105 , po2106 , po2107 , po2108 , po2109 , po2110 , po2111 , po2112 , po2113 , po2114 , po2115 , po2116 , po2117 , po2118 , po2119 , po2120 , po2121 , po2122 , po2123 , po2124 , po2125 , po2126 , po2127 , po2128 , po2129 , po2130 , po2131 , po2132 , po2133 , po2134 , po2135 , po2136 , po2137 , po2138 , po2139 , po2140 , po2141 , po2142 , po2143 , po2144 , po2145 , po2146 , po2147 , po2148 , po2149 , po2150 , po2151 , po2152 , po2153 , po2154 , po2155 , po2156 , po2157 , po2158 , po2159 , po2160 , po2161 , po2162 , po2163 , po2164 , po2165 , po2166 , po2167 , po2168 , po2169 , po2170 , po2171 , po2172 , po2173 , po2174 , po2175 , po2176 , po2177 , po2178 , po2179 , po2180 , po2181 , po2182 , po2183 , po2184 , po2185 , po2186 , po2187 , po2188 , po2189 , po2190 , po2191 , po2192 , po2193 , po2194 , po2195 , po2196 , po2197 , po2198 , po2199 , po2200 , po2201 , po2202 , po2203 , po2204 , po2205 , po2206 , po2207 , po2208 , po2209 , po2210 , po2211 , po2212 , po2213 , po2214 , po2215 , po2216 , po2217 , po2218 , po2219 , po2220 , po2221 , po2222 , po2223 , po2224 , po2225 , po2226 , po2227 , po2228 , po2229 , po2230 , po2231 , po2232 , po2233 , po2234 , po2235 , po2236 , po2237 , po2238 , po2239 , po2240 , po2241 , po2242 , po2243 , po2244 , po2245 , po2246 , po2247 , po2248 , po2249 , po2250 , po2251 , po2252 , po2253 , po2254 , po2255 , po2256 , po2257 , po2258 , po2259 , po2260 , po2261 , po2262 , po2263 , po2264 , po2265 , po2266 , po2267 , po2268 , po2269 , po2270 , po2271 , po2272 , po2273 , po2274 , po2275 , po2276 , po2277 , po2278 , po2279 , po2280 , po2281 , po2282 , po2283 , po2284 , po2285 , po2286 , po2287 , po2288 , po2289 , po2290 , po2291 , po2292 , po2293 , po2294 , po2295 , po2296 , po2297 , po2298 , po2299 , po2300 , po2301 , po2302 , po2303 , po2304 , po2305 , po2306 , po2307 , po2308 , po2309 , po2310 , po2311 , po2312 , po2313 , po2314 , po2315 , po2316 , po2317 , po2318 , po2319 , po2320 , po2321 , po2322 , po2323 , po2324 , po2325 , po2326 , po2327 , po2328 , po2329 , po2330 , po2331 , po2332 , po2333 , po2334 , po2335 , po2336 , po2337 , po2338 , po2339 , po2340 , po2341 , po2342 , po2343 , po2344 , po2345 , po2346 , po2347 , po2348 , po2349 , po2350 , po2351 , po2352 , po2353 , po2354 , po2355 , po2356 , po2357 , po2358 , po2359 , po2360 , po2361 , po2362 , po2363 , po2364 , po2365 , po2366 , po2367 , po2368 , po2369 , po2370 , po2371 , po2372 , po2373 , po2374 , po2375 , po2376 , po2377 , po2378 , po2379 , po2380 , po2381 , po2382 , po2383 , po2384 , po2385 , po2386 , po2387 , po2388 , po2389 , po2390 , po2391 , po2392 , po2393 , po2394 , po2395 , po2396 , po2397 , po2398 , po2399 , po2400 , po2401 , po2402 , po2403 , po2404 , po2405 , po2406 , po2407 , po2408 , po2409 , po2410 , po2411 , po2412 , po2413 , po2414 , po2415 , po2416 , po2417 , po2418 , po2419 , po2420 , po2421 , po2422 , po2423 , po2424 , po2425 , po2426 , po2427 , po2428 , po2429 , po2430 , po2431 , po2432 , po2433 , po2434 , po2435 , po2436 , po2437 , po2438 , po2439 , po2440 , po2441 , po2442 , po2443 , po2444 , po2445 , po2446 , po2447 , po2448 , po2449 , po2450 , po2451 , po2452 , po2453 , po2454 , po2455 , po2456 , po2457 , po2458 , po2459 , po2460 , po2461 , po2462 , po2463 , po2464 , po2465 , po2466 , po2467 , po2468 , po2469 , po2470 , po2471 , po2472 , po2473 , po2474 , po2475 , po2476 , po2477 , po2478 , po2479 , po2480 , po2481 , po2482 , po2483 , po2484 , po2485 , po2486 , po2487 , po2488 , po2489 , po2490 , po2491 , po2492 , po2493 , po2494 , po2495 , po2496 , po2497 , po2498 , po2499 , po2500 , po2501 , po2502 , po2503 , po2504 , po2505 , po2506 , po2507 , po2508 , po2509 , po2510 , po2511 , po2512 , po2513 , po2514 , po2515 , po2516 , po2517 , po2518 , po2519 , po2520 , po2521 , po2522 , po2523 , po2524 , po2525 , po2526 , po2527 , po2528 , po2529 , po2530 , po2531 , po2532 , po2533 , po2534 , po2535 , po2536 , po2537 , po2538 , po2539 , po2540 , po2541 , po2542 , po2543 , po2544 , po2545 , po2546 , po2547 , po2548 , po2549 , po2550 , po2551 , po2552 , po2553 , po2554 , po2555 , po2556 , po2557 , po2558 , po2559 , po2560 , po2561 , po2562 , po2563 , po2564 , po2565 , po2566 , po2567 , po2568 , po2569 , po2570 , po2571 , po2572 , po2573 , po2574 , po2575 , po2576 , po2577 , po2578 , po2579 , po2580 , po2581 , po2582 , po2583 , po2584 , po2585 , po2586 , po2587 , po2588 , po2589 , po2590 , po2591 , po2592 , po2593 , po2594 , po2595 , po2596 , po2597 , po2598 , po2599 , po2600 , po2601 , po2602 , po2603 , po2604 , po2605 , po2606 , po2607 , po2608 , po2609 , po2610 , po2611 , po2612 , po2613 , po2614 , po2615 , po2616 , po2617 , po2618 , po2619 , po2620 , po2621 , po2622 , po2623 , po2624 , po2625 , po2626 , po2627 , po2628 , po2629 , po2630 , po2631 , po2632 , po2633 , po2634 , po2635 , po2636 , po2637 , po2638 , po2639 , po2640 , po2641 , po2642 , po2643 , po2644 , po2645 , po2646 , po2647 , po2648 , po2649 , po2650 , po2651 , po2652 , po2653 , po2654 , po2655 , po2656 , po2657 , po2658 , po2659 , po2660 , po2661 , po2662 , po2663 , po2664 , po2665 , po2666 , po2667 , po2668 , po2669 , po2670 , po2671 , po2672 , po2673 , po2674 , po2675 , po2676 , po2677 , po2678 , po2679 , po2680 , po2681 , po2682 , po2683 , po2684 , po2685 , po2686 , po2687 , po2688 , po2689 , po2690 , po2691 , po2692 , po2693 , po2694 , po2695 , po2696 , po2697 , po2698 , po2699 , po2700 , po2701 , po2702 , po2703 , po2704 , po2705 , po2706 , po2707 , po2708 , po2709 , po2710 , po2711 , po2712 , po2713 , po2714 , po2715 , po2716 , po2717 , po2718 , po2719 , po2720 , po2721 , po2722 , po2723 , po2724 , po2725 , po2726 , po2727 , po2728 , po2729 , po2730 , po2731 , po2732 , po2733 , po2734 , po2735 , po2736 , po2737 , po2738 , po2739 , po2740 , po2741 , po2742 , po2743 , po2744 , po2745 , po2746 , po2747 , po2748 , po2749 , po2750 , po2751 , po2752 , po2753 , po2754 , po2755 , po2756 , po2757 , po2758 , po2759 , po2760 , po2761 , po2762 , po2763 , po2764 , po2765 , po2766 , po2767 , po2768 , po2769 , po2770 , po2771 , po2772 , po2773 , po2774 , po2775 , po2776 , po2777 , po2778 , po2779 , po2780 , po2781 , po2782 , po2783 , po2784 , po2785 , po2786 , po2787 , po2788 , po2789 , po2790 , po2791 , po2792 , po2793 , po2794 , po2795 , po2796 , po2797 , po2798 , po2799 , po2800 , po2801 , po2802 , po2803 , po2804 , po2805 , po2806 , po2807 , po2808 , po2809 , po2810 , po2811 , po2812 , po2813 , po2814 , po2815 , po2816 , po2817 , po2818 , po2819 , po2820 , po2821 , po2822 , po2823 , po2824 , po2825 , po2826 , po2827 , po2828 , po2829 , po2830 , po2831 , po2832 , po2833 , po2834 , po2835 , po2836 , po2837 , po2838 , po2839 , po2840 , po2841 , po2842 , po2843 , po2844 , po2845 , po2846 , po2847 , po2848 , po2849 , po2850 , po2851 , po2852 , po2853 , po2854 , po2855 , po2856 , po2857 , po2858 , po2859 , po2860 , po2861 , po2862 , po2863 , po2864 , po2865 , po2866 , po2867 , po2868 , po2869 , po2870 , po2871 , po2872 , po2873 , po2874 , po2875 , po2876 , po2877 , po2878 , po2879 , po2880 , po2881 , po2882 , po2883 , po2884 , po2885 , po2886 , po2887 , po2888 , po2889 , po2890 , po2891 , po2892 , po2893 , po2894 , po2895 , po2896 , po2897 , po2898 , po2899 , po2900 , po2901 , po2902 , po2903 , po2904 , po2905 , po2906 , po2907 , po2908 , po2909 , po2910 , po2911 , po2912 , po2913 , po2914 , po2915 , po2916 , po2917 , po2918 , po2919 , po2920 , po2921 , po2922 , po2923 , po2924 , po2925 , po2926 , po2927 , po2928 , po2929 , po2930 , po2931 , po2932 , po2933 , po2934 , po2935 , po2936 , po2937 , po2938 , po2939 , po2940 , po2941 , po2942 , po2943 , po2944 , po2945 , po2946 , po2947 , po2948 , po2949 , po2950 , po2951 , po2952 , po2953 , po2954 , po2955 , po2956 , po2957 , po2958 , po2959 , po2960 , po2961 , po2962 , po2963 , po2964 , po2965 , po2966 , po2967 , po2968 , po2969 , po2970 , po2971 , po2972 , po2973 , po2974 , po2975 , po2976 , po2977 , po2978 , po2979 , po2980 , po2981 , po2982 , po2983 , po2984 , po2985 , po2986 , po2987 , po2988 , po2989 , po2990 , po2991 , po2992 , po2993 , po2994 , po2995 , po2996 , po2997 , po2998 , po2999 , po3000 , po3001 , po3002 , po3003 , po3004 , po3005 , po3006 , po3007 , po3008 , po3009 , po3010 , po3011 , po3012 , po3013 , po3014 , po3015 , po3016 , po3017 , po3018 , po3019 , po3020 , po3021 , po3022 , po3023 , po3024 , po3025 , po3026 , po3027 , po3028 , po3029 , po3030 , po3031 , po3032 , po3033 , po3034 , po3035 , po3036 , po3037 , po3038 , po3039 , po3040 , po3041 , po3042 , po3043 , po3044 , po3045 , po3046 , po3047 , po3048 , po3049 , po3050 , po3051 , po3052 , po3053 , po3054 , po3055 , po3056 , po3057 , po3058 , po3059 , po3060 , po3061 , po3062 , po3063 , po3064 , po3065 , po3066 , po3067 , po3068 , po3069 , po3070 , po3071 , po3072 , po3073 , po3074 , po3075 , po3076 , po3077 , po3078 , po3079 , po3080 , po3081 , po3082 , po3083 , po3084 , po3085 , po3086 , po3087 , po3088 , po3089 , po3090 , po3091 , po3092 , po3093 , po3094 , po3095 , po3096 , po3097 , po3098 , po3099 , po3100 , po3101 , po3102 , po3103 , po3104 , po3105 , po3106 , po3107 , po3108 , po3109 , po3110 , po3111 , po3112 , po3113 , po3114 , po3115 , po3116 , po3117 , po3118 , po3119 , po3120 , po3121 , po3122 , po3123 , po3124 , po3125 , po3126 , po3127 , po3128 , po3129 , po3130 , po3131 , po3132 , po3133 , po3134 , po3135 , po3136 , po3137 , po3138 , po3139 , po3140 , po3141 , po3142 , po3143 , po3144 , po3145 , po3146 , po3147 , po3148 , po3149 , po3150 , po3151 , po3152 , po3153 , po3154 , po3155 , po3156 , po3157 , po3158 , po3159 , po3160 , po3161 , po3162 , po3163 , po3164 , po3165 , po3166 , po3167 , po3168 , po3169 , po3170 , po3171 , po3172 , po3173 , po3174 , po3175 , po3176 , po3177 , po3178 , po3179 , po3180 , po3181 , po3182 , po3183 , po3184 , po3185 , po3186 , po3187 , po3188 , po3189 , po3190 , po3191 , po3192 , po3193 , po3194 , po3195 , po3196 , po3197 , po3198 , po3199 , po3200 , po3201 , po3202 , po3203 , po3204 , po3205 , po3206 , po3207 , po3208 , po3209 , po3210 , po3211 , po3212 , po3213 , po3214 , po3215 , po3216 , po3217 , po3218 , po3219 , po3220 , po3221 , po3222 , po3223 , po3224 , po3225 , po3226 , po3227 , po3228 , po3229 , po3230 , po3231 , po3232 , po3233 , po3234 , po3235 , po3236 , po3237 , po3238 , po3239 , po3240 , po3241 , po3242 , po3243 , po3244 , po3245 , po3246 , po3247 , po3248 , po3249 , po3250 , po3251 , po3252 , po3253 , po3254 , po3255 , po3256 , po3257 , po3258 , po3259 , po3260 , po3261 , po3262 , po3263 , po3264 , po3265 , po3266 , po3267 , po3268 , po3269 , po3270 , po3271 , po3272 , po3273 , po3274 , po3275 , po3276 , po3277 , po3278 , po3279 , po3280 , po3281 , po3282 , po3283 , po3284 , po3285 , po3286 , po3287 , po3288 , po3289 , po3290 , po3291 , po3292 , po3293 , po3294 , po3295 , po3296 , po3297 , po3298 , po3299 , po3300 , po3301 , po3302 , po3303 , po3304 , po3305 , po3306 , po3307 , po3308 , po3309 , po3310 , po3311 , po3312 , po3313 , po3314 , po3315 , po3316 , po3317 , po3318 , po3319 , po3320 , po3321 , po3322 , po3323 , po3324 , po3325 , po3326 , po3327 ;
  reg lo0000 , lo0001 , lo0002 , lo0003 , lo0004 , lo0005 , lo0006 , lo0007 , lo0008 , lo0009 , lo0010 , lo0011 , lo0012 , lo0013 , lo0014 , lo0015 , lo0016 , lo0017 , lo0018 , lo0019 , lo0020 , lo0021 , lo0022 , lo0023 , lo0024 , lo0025 , lo0026 , lo0027 , lo0028 , lo0029 , lo0030 , lo0031 , lo0032 , lo0033 , lo0034 , lo0035 , lo0036 , lo0037 , lo0038 , lo0039 , lo0040 , lo0041 , lo0042 , lo0043 , lo0044 , lo0045 , lo0046 , lo0047 , lo0048 , lo0049 , lo0050 , lo0051 , lo0052 , lo0053 , lo0054 , lo0055 , lo0056 , lo0057 , lo0058 , lo0059 , lo0060 , lo0061 , lo0062 , lo0063 , lo0064 , lo0065 , lo0066 , lo0067 , lo0068 , lo0069 , lo0070 , lo0071 , lo0072 , lo0073 , lo0074 , lo0075 , lo0076 , lo0077 , lo0078 , lo0079 , lo0080 , lo0081 , lo0082 , lo0083 , lo0084 , lo0085 , lo0086 , lo0087 , lo0088 , lo0089 , lo0090 , lo0091 , lo0092 , lo0093 , lo0094 , lo0095 , lo0096 , lo0097 , lo0098 , lo0099 , lo0100 , lo0101 , lo0102 , lo0103 , lo0104 , lo0105 , lo0106 , lo0107 , lo0108 , lo0109 , lo0110 , lo0111 , lo0112 , lo0113 , lo0114 , lo0115 , lo0116 , lo0117 , lo0118 , lo0119 , lo0120 , lo0121 , lo0122 , lo0123 , lo0124 , lo0125 , lo0126 , lo0127 , lo0128 , lo0129 , lo0130 , lo0131 , lo0132 , lo0133 , lo0134 , lo0135 , lo0136 , lo0137 , lo0138 , lo0139 , lo0140 , lo0141 , lo0142 , lo0143 , lo0144 , lo0145 , lo0146 , lo0147 , lo0148 , lo0149 , lo0150 , lo0151 , lo0152 , lo0153 , lo0154 , lo0155 , lo0156 , lo0157 , lo0158 , lo0159 , lo0160 , lo0161 , lo0162 , lo0163 , lo0164 , lo0165 , lo0166 , lo0167 , lo0168 , lo0169 , lo0170 , lo0171 , lo0172 , lo0173 , lo0174 , lo0175 , lo0176 , lo0177 , lo0178 , lo0179 , lo0180 , lo0181 , lo0182 , lo0183 , lo0184 , lo0185 , lo0186 , lo0187 , lo0188 , lo0189 , lo0190 , lo0191 , lo0192 , lo0193 , lo0194 , lo0195 , lo0196 , lo0197 , lo0198 , lo0199 , lo0200 , lo0201 , lo0202 , lo0203 , lo0204 , lo0205 , lo0206 , lo0207 , lo0208 , lo0209 , lo0210 , lo0211 , lo0212 , lo0213 , lo0214 , lo0215 , lo0216 , lo0217 , lo0218 , lo0219 , lo0220 , lo0221 , lo0222 , lo0223 , lo0224 , lo0225 , lo0226 , lo0227 , lo0228 , lo0229 , lo0230 , lo0231 , lo0232 , lo0233 , lo0234 , lo0235 , lo0236 , lo0237 , lo0238 , lo0239 , lo0240 , lo0241 , lo0242 , lo0243 , lo0244 , lo0245 , lo0246 , lo0247 , lo0248 , lo0249 , lo0250 , lo0251 , lo0252 , lo0253 , lo0254 , lo0255 , lo0256 , lo0257 , lo0258 , lo0259 , lo0260 , lo0261 , lo0262 , lo0263 , lo0264 , lo0265 , lo0266 , lo0267 , lo0268 , lo0269 , lo0270 , lo0271 , lo0272 , lo0273 , lo0274 , lo0275 , lo0276 , lo0277 , lo0278 , lo0279 , lo0280 , lo0281 , lo0282 , lo0283 , lo0284 , lo0285 , lo0286 , lo0287 , lo0288 , lo0289 , lo0290 , lo0291 , lo0292 , lo0293 , lo0294 , lo0295 , lo0296 , lo0297 , lo0298 , lo0299 , lo0300 , lo0301 , lo0302 , lo0303 , lo0304 , lo0305 , lo0306 , lo0307 , lo0308 , lo0309 , lo0310 , lo0311 , lo0312 , lo0313 , lo0314 , lo0315 , lo0316 , lo0317 , lo0318 , lo0319 , lo0320 , lo0321 , lo0322 , lo0323 , lo0324 , lo0325 , lo0326 , lo0327 , lo0328 , lo0329 , lo0330 , lo0331 , lo0332 , lo0333 , lo0334 , lo0335 , lo0336 , lo0337 , lo0338 , lo0339 , lo0340 , lo0341 , lo0342 , lo0343 , lo0344 , lo0345 , lo0346 , lo0347 , lo0348 , lo0349 , lo0350 , lo0351 , lo0352 , lo0353 , lo0354 , lo0355 , lo0356 , lo0357 , lo0358 , lo0359 , lo0360 , lo0361 , lo0362 , lo0363 , lo0364 , lo0365 , lo0366 , lo0367 , lo0368 , lo0369 , lo0370 , lo0371 , lo0372 , lo0373 , lo0374 , lo0375 , lo0376 , lo0377 , lo0378 , lo0379 , lo0380 , lo0381 , lo0382 , lo0383 , lo0384 , lo0385 , lo0386 , lo0387 , lo0388 , lo0389 , lo0390 , lo0391 , lo0392 , lo0393 , lo0394 , lo0395 , lo0396 , lo0397 , lo0398 , lo0399 , lo0400 , lo0401 , lo0402 , lo0403 , lo0404 , lo0405 , lo0406 , lo0407 , lo0408 , lo0409 , lo0410 , lo0411 , lo0412 , lo0413 , lo0414 , lo0415 , lo0416 , lo0417 , lo0418 , lo0419 , lo0420 , lo0421 , lo0422 , lo0423 , lo0424 , lo0425 , lo0426 , lo0427 , lo0428 , lo0429 , lo0430 , lo0431 , lo0432 , lo0433 , lo0434 , lo0435 , lo0436 , lo0437 , lo0438 , lo0439 , lo0440 , lo0441 , lo0442 , lo0443 , lo0444 , lo0445 , lo0446 , lo0447 , lo0448 , lo0449 , lo0450 , lo0451 , lo0452 , lo0453 , lo0454 , lo0455 , lo0456 , lo0457 , lo0458 , lo0459 , lo0460 , lo0461 , lo0462 , lo0463 , lo0464 , lo0465 , lo0466 , lo0467 , lo0468 , lo0469 , lo0470 , lo0471 , lo0472 , lo0473 , lo0474 , lo0475 , lo0476 , lo0477 , lo0478 , lo0479 , lo0480 , lo0481 , lo0482 , lo0483 , lo0484 , lo0485 , lo0486 , lo0487 , lo0488 , lo0489 , lo0490 , lo0491 , lo0492 , lo0493 , lo0494 , lo0495 , lo0496 , lo0497 , lo0498 , lo0499 , lo0500 , lo0501 , lo0502 , lo0503 , lo0504 , lo0505 , lo0506 , lo0507 , lo0508 , lo0509 , lo0510 , lo0511 , lo0512 , lo0513 , lo0514 , lo0515 , lo0516 , lo0517 , lo0518 , lo0519 , lo0520 , lo0521 , lo0522 , lo0523 , lo0524 , lo0525 , lo0526 , lo0527 , lo0528 , lo0529 , lo0530 , lo0531 , lo0532 , lo0533 , lo0534 , lo0535 , lo0536 , lo0537 , lo0538 , lo0539 , lo0540 , lo0541 , lo0542 , lo0543 , lo0544 , lo0545 , lo0546 , lo0547 , lo0548 , lo0549 , lo0550 , lo0551 , lo0552 , lo0553 , lo0554 , lo0555 , lo0556 , lo0557 , lo0558 , lo0559 , lo0560 , lo0561 , lo0562 , lo0563 , lo0564 , lo0565 , lo0566 , lo0567 , lo0568 , lo0569 , lo0570 , lo0571 , lo0572 , lo0573 , lo0574 , lo0575 , lo0576 , lo0577 , lo0578 , lo0579 , lo0580 , lo0581 , lo0582 , lo0583 , lo0584 , lo0585 , lo0586 , lo0587 , lo0588 , lo0589 , lo0590 , lo0591 , lo0592 , lo0593 , lo0594 , lo0595 , lo0596 , lo0597 , lo0598 , lo0599 , lo0600 , lo0601 , lo0602 , lo0603 , lo0604 , lo0605 , lo0606 , lo0607 , lo0608 , lo0609 , lo0610 , lo0611 , lo0612 , lo0613 , lo0614 , lo0615 , lo0616 , lo0617 , lo0618 , lo0619 , lo0620 , lo0621 , lo0622 , lo0623 , lo0624 , lo0625 , lo0626 , lo0627 , lo0628 , lo0629 , lo0630 , lo0631 , lo0632 , lo0633 , lo0634 , lo0635 , lo0636 , lo0637 , lo0638 , lo0639 , lo0640 , lo0641 , lo0642 , lo0643 , lo0644 , lo0645 , lo0646 , lo0647 , lo0648 , lo0649 , lo0650 , lo0651 , lo0652 , lo0653 , lo0654 , lo0655 , lo0656 , lo0657 , lo0658 , lo0659 , lo0660 , lo0661 , lo0662 , lo0663 , lo0664 , lo0665 , lo0666 , lo0667 , lo0668 , lo0669 , lo0670 , lo0671 , lo0672 , lo0673 , lo0674 , lo0675 , lo0676 , lo0677 , lo0678 , lo0679 , lo0680 , lo0681 , lo0682 , lo0683 , lo0684 , lo0685 , lo0686 , lo0687 , lo0688 , lo0689 , lo0690 , lo0691 , lo0692 , lo0693 , lo0694 , lo0695 , lo0696 , lo0697 , lo0698 , lo0699 , lo0700 , lo0701 , lo0702 , lo0703 , lo0704 , lo0705 , lo0706 , lo0707 , lo0708 , lo0709 , lo0710 , lo0711 , lo0712 , lo0713 , lo0714 , lo0715 , lo0716 , lo0717 , lo0718 , lo0719 , lo0720 , lo0721 , lo0722 , lo0723 , lo0724 , lo0725 , lo0726 , lo0727 , lo0728 , lo0729 , lo0730 , lo0731 , lo0732 , lo0733 , lo0734 , lo0735 , lo0736 , lo0737 , lo0738 , lo0739 , lo0740 , lo0741 , lo0742 , lo0743 , lo0744 , lo0745 , lo0746 , lo0747 , lo0748 , lo0749 , lo0750 , lo0751 , lo0752 , lo0753 , lo0754 , lo0755 , lo0756 , lo0757 , lo0758 , lo0759 , lo0760 , lo0761 , lo0762 , lo0763 , lo0764 , lo0765 , lo0766 , lo0767 , lo0768 , lo0769 , lo0770 , lo0771 , lo0772 , lo0773 , lo0774 , lo0775 , lo0776 , lo0777 , lo0778 , lo0779 , lo0780 , lo0781 , lo0782 , lo0783 , lo0784 , lo0785 , lo0786 , lo0787 , lo0788 , lo0789 , lo0790 , lo0791 , lo0792 , lo0793 , lo0794 , lo0795 , lo0796 , lo0797 , lo0798 , lo0799 , lo0800 , lo0801 , lo0802 , lo0803 , lo0804 , lo0805 , lo0806 , lo0807 , lo0808 , lo0809 , lo0810 , lo0811 , lo0812 , lo0813 , lo0814 , lo0815 , lo0816 , lo0817 , lo0818 , lo0819 , lo0820 , lo0821 , lo0822 , lo0823 , lo0824 , lo0825 , lo0826 , lo0827 , lo0828 , lo0829 , lo0830 , lo0831 , lo0832 , lo0833 , lo0834 , lo0835 , lo0836 , lo0837 , lo0838 , lo0839 , lo0840 , lo0841 , lo0842 , lo0843 , lo0844 , lo0845 , lo0846 , lo0847 , lo0848 , lo0849 , lo0850 , lo0851 , lo0852 , lo0853 , lo0854 , lo0855 , lo0856 , lo0857 , lo0858 , lo0859 , lo0860 , lo0861 , lo0862 , lo0863 , lo0864 , lo0865 , lo0866 , lo0867 , lo0868 , lo0869 , lo0870 , lo0871 , lo0872 , lo0873 , lo0874 , lo0875 , lo0876 , lo0877 , lo0878 , lo0879 , lo0880 , lo0881 , lo0882 , lo0883 , lo0884 , lo0885 , lo0886 , lo0887 , lo0888 , lo0889 , lo0890 , lo0891 , lo0892 , lo0893 , lo0894 , lo0895 , lo0896 , lo0897 , lo0898 , lo0899 , lo0900 , lo0901 , lo0902 , lo0903 , lo0904 , lo0905 , lo0906 , lo0907 , lo0908 , lo0909 , lo0910 , lo0911 , lo0912 , lo0913 , lo0914 , lo0915 , lo0916 , lo0917 , lo0918 , lo0919 , lo0920 , lo0921 , lo0922 , lo0923 , lo0924 , lo0925 , lo0926 , lo0927 , lo0928 , lo0929 , lo0930 , lo0931 , lo0932 , lo0933 , lo0934 , lo0935 , lo0936 , lo0937 , lo0938 , lo0939 , lo0940 , lo0941 , lo0942 , lo0943 , lo0944 , lo0945 , lo0946 , lo0947 , lo0948 , lo0949 , lo0950 , lo0951 , lo0952 , lo0953 , lo0954 , lo0955 , lo0956 , lo0957 , lo0958 , lo0959 , lo0960 , lo0961 , lo0962 , lo0963 , lo0964 , lo0965 , lo0966 , lo0967 , lo0968 , lo0969 , lo0970 , lo0971 , lo0972 , lo0973 , lo0974 , lo0975 , lo0976 , lo0977 , lo0978 , lo0979 , lo0980 , lo0981 , lo0982 , lo0983 , lo0984 , lo0985 , lo0986 , lo0987 , lo0988 , lo0989 , lo0990 , lo0991 , lo0992 , lo0993 , lo0994 , lo0995 , lo0996 , lo0997 , lo0998 , lo0999 , lo1000 , lo1001 , lo1002 , lo1003 , lo1004 , lo1005 , lo1006 , lo1007 , lo1008 , lo1009 , lo1010 , lo1011 , lo1012 , lo1013 , lo1014 , lo1015 , lo1016 , lo1017 , lo1018 , lo1019 , lo1020 , lo1021 , lo1022 , lo1023 , lo1024 , lo1025 , lo1026 , lo1027 , lo1028 , lo1029 , lo1030 , lo1031 , lo1032 , lo1033 , lo1034 , lo1035 , lo1036 , lo1037 , lo1038 , lo1039 , lo1040 , lo1041 , lo1042 , lo1043 , lo1044 , lo1045 , lo1046 , lo1047 , lo1048 , lo1049 , lo1050 , lo1051 , lo1052 , lo1053 , lo1054 , lo1055 , lo1056 , lo1057 , lo1058 , lo1059 , lo1060 , lo1061 , lo1062 , lo1063 , lo1064 , lo1065 , lo1066 , lo1067 , lo1068 , lo1069 , lo1070 , lo1071 , lo1072 , lo1073 , lo1074 , lo1075 , lo1076 , lo1077 , lo1078 , lo1079 , lo1080 , lo1081 , lo1082 , lo1083 , lo1084 , lo1085 , lo1086 , lo1087 , lo1088 , lo1089 , lo1090 , lo1091 , lo1092 , lo1093 , lo1094 , lo1095 , lo1096 , lo1097 , lo1098 , lo1099 , lo1100 , lo1101 , lo1102 , lo1103 , lo1104 , lo1105 , lo1106 , lo1107 , lo1108 , lo1109 , lo1110 , lo1111 , lo1112 , lo1113 , lo1114 , lo1115 , lo1116 , lo1117 , lo1118 , lo1119 , lo1120 , lo1121 , lo1122 , lo1123 , lo1124 , lo1125 , lo1126 , lo1127 , lo1128 , lo1129 , lo1130 , lo1131 , lo1132 , lo1133 , lo1134 , lo1135 , lo1136 , lo1137 , lo1138 , lo1139 , lo1140 , lo1141 , lo1142 , lo1143 , lo1144 , lo1145 , lo1146 , lo1147 , lo1148 , lo1149 , lo1150 , lo1151 , lo1152 , lo1153 , lo1154 , lo1155 , lo1156 , lo1157 , lo1158 , lo1159 , lo1160 , lo1161 , lo1162 , lo1163 , lo1164 , lo1165 , lo1166 , lo1167 , lo1168 , lo1169 , lo1170 , lo1171 , lo1172 , lo1173 , lo1174 , lo1175 , lo1176 , lo1177 , lo1178 , lo1179 , lo1180 , lo1181 , lo1182 , lo1183 , lo1184 , lo1185 , lo1186 , lo1187 , lo1188 , lo1189 , lo1190 , lo1191 , lo1192 , lo1193 , lo1194 , lo1195 , lo1196 , lo1197 , lo1198 , lo1199 , lo1200 , lo1201 , lo1202 , lo1203 , lo1204 , lo1205 , lo1206 , lo1207 , lo1208 , lo1209 , lo1210 , lo1211 , lo1212 , lo1213 , lo1214 , lo1215 , lo1216 , lo1217 , lo1218 , lo1219 , lo1220 , lo1221 , lo1222 , lo1223 , lo1224 , lo1225 , lo1226 , lo1227 , lo1228 , lo1229 , lo1230 , lo1231 , lo1232 , lo1233 , lo1234 , lo1235 , lo1236 , lo1237 , lo1238 , lo1239 , lo1240 , lo1241 , lo1242 , lo1243 , lo1244 , lo1245 , lo1246 , lo1247 , lo1248 , lo1249 , lo1250 , lo1251 , lo1252 , lo1253 , lo1254 , lo1255 , lo1256 , lo1257 , lo1258 , lo1259 , lo1260 , lo1261 , lo1262 , lo1263 , lo1264 , lo1265 , lo1266 , lo1267 , lo1268 , lo1269 , lo1270 , lo1271 , lo1272 , lo1273 , lo1274 , lo1275 , lo1276 , lo1277 , lo1278 , lo1279 , lo1280 , lo1281 , lo1282 , lo1283 , lo1284 , lo1285 , lo1286 , lo1287 , lo1288 , lo1289 , lo1290 , lo1291 , lo1292 , lo1293 , lo1294 , lo1295 , lo1296 , lo1297 , lo1298 , lo1299 , lo1300 , lo1301 , lo1302 , lo1303 , lo1304 , lo1305 , lo1306 , lo1307 , lo1308 , lo1309 , lo1310 , lo1311 , lo1312 , lo1313 , lo1314 , lo1315 , lo1316 , lo1317 , lo1318 , lo1319 , lo1320 , lo1321 , lo1322 , lo1323 , lo1324 , lo1325 , lo1326 , lo1327 , lo1328 , lo1329 , lo1330 , lo1331 , lo1332 , lo1333 , lo1334 , lo1335 , lo1336 , lo1337 , lo1338 , lo1339 , lo1340 , lo1341 , lo1342 , lo1343 , lo1344 , lo1345 , lo1346 , lo1347 , lo1348 , lo1349 , lo1350 , lo1351 , lo1352 , lo1353 , lo1354 , lo1355 , lo1356 , lo1357 , lo1358 , lo1359 , lo1360 , lo1361 , lo1362 , lo1363 , lo1364 , lo1365 , lo1366 , lo1367 , lo1368 , lo1369 , lo1370 , lo1371 , lo1372 , lo1373 , lo1374 , lo1375 , lo1376 , lo1377 , lo1378 , lo1379 , lo1380 , lo1381 , lo1382 , lo1383 , lo1384 , lo1385 , lo1386 , lo1387 , lo1388 , lo1389 , lo1390 , lo1391 , lo1392 , lo1393 , lo1394 , lo1395 , lo1396 , lo1397 , lo1398 , lo1399 , lo1400 , lo1401 , lo1402 , lo1403 , lo1404 , lo1405 , lo1406 , lo1407 , lo1408 , lo1409 , lo1410 , lo1411 , lo1412 , lo1413 , lo1414 , lo1415 , lo1416 , lo1417 , lo1418 , lo1419 , lo1420 , lo1421 , lo1422 , lo1423 , lo1424 , lo1425 , lo1426 , lo1427 , lo1428 , lo1429 , lo1430 , lo1431 , lo1432 , lo1433 , lo1434 , lo1435 , lo1436 , lo1437 , lo1438 , lo1439 , lo1440 , lo1441 , lo1442 , lo1443 , lo1444 , lo1445 , lo1446 , lo1447 , lo1448 , lo1449 , lo1450 , lo1451 , lo1452 , lo1453 , lo1454 , lo1455 , lo1456 , lo1457 , lo1458 , lo1459 , lo1460 , lo1461 , lo1462 , lo1463 , lo1464 , lo1465 , lo1466 , lo1467 , lo1468 , lo1469 , lo1470 , lo1471 , lo1472 , lo1473 , lo1474 , lo1475 , lo1476 ;
  wire new_n1942, new_n1943, new_n1944, new_n1945, new_n1946, new_n1947, new_n1948, new_n1949, new_n1950, new_n1951, new_n1952, new_n1953, new_n1954, new_n1955, new_n1956, new_n1957, new_n1958, new_n1959, new_n1960, new_n1961, new_n1962, new_n1963, new_n1964, new_n1965, new_n1966, new_n1967, new_n1968, new_n1969, new_n1970, new_n1971, new_n1972, new_n1973, new_n1974, new_n1975, new_n1976, new_n1977, new_n1978, new_n1979, new_n1980, new_n1981, new_n1982, new_n1983, new_n1984, new_n1985, new_n1986, new_n1987, new_n1988, new_n1989, new_n1990, new_n1991, new_n1992, new_n1993, new_n1994, new_n1995, new_n1996, new_n1997, new_n1998, new_n1999, new_n2000, new_n2001, new_n2002, new_n2003, new_n2004, new_n2005, new_n2006, new_n2007, new_n2008, new_n2009, new_n2010, new_n2011, new_n2012, new_n2013, new_n2014, new_n2015, new_n2016, new_n2017, new_n2018, new_n2019, new_n2020, new_n2021, new_n2022, new_n2023, new_n2024, new_n2025, new_n2026, new_n2027, new_n2028, new_n2029, new_n2030, new_n2031, new_n2032, new_n2033, new_n2034, new_n2035, new_n2036, new_n2037, new_n2038, new_n2039, new_n2040, new_n2041, new_n2042, new_n2043, new_n2044, new_n2045, new_n2046, new_n2047, new_n2048, new_n2049, new_n2050, new_n2051, new_n2052, new_n2053, new_n2054, new_n2055, new_n2056, new_n2057, new_n2058, new_n2059, new_n2060, new_n2061, new_n2062, new_n2063, new_n2064, new_n2065, new_n2066, new_n2067, new_n2068, new_n2069, new_n2070, new_n2071, new_n2072, new_n2073, new_n2074, new_n2075, new_n2076, new_n2077, new_n2078, new_n2079, new_n2080, new_n2081, new_n2082, new_n2083, new_n2084, new_n2085, new_n2086, new_n2087, new_n2088, new_n2089, new_n2090, new_n2091, new_n2092, new_n2093, new_n2094, new_n2095, new_n2096, new_n2097, new_n2098, new_n2099, new_n2100, new_n2101, new_n2102, new_n2103, new_n2104, new_n2105, new_n2106, new_n2107, new_n2108, new_n2109, new_n2110, new_n2111, new_n2112, new_n2113, new_n2114, new_n2115, new_n2116, new_n2117, new_n2118, new_n2119, new_n2120, new_n2121, new_n2122, new_n2123, new_n2124, new_n2125, new_n2126, new_n2127, new_n2128, new_n2129, new_n2130, new_n2131, new_n2132, new_n2133, new_n2134, new_n2135, new_n2136, new_n2137, new_n2138, new_n2139, new_n2140, new_n2141, new_n2142, new_n2143, new_n2144, new_n2145, new_n2146, new_n2147, new_n2148, new_n2149, new_n2150, new_n2151, new_n2152, new_n2153, new_n2154, new_n2155, new_n2156, new_n2157, new_n2158, new_n2159, new_n2160, new_n2161, new_n2162, new_n2163, new_n2164, new_n2165, new_n2166, new_n2167, new_n2168, new_n2169, new_n2170, new_n2171, new_n2172, new_n2173, new_n2174, new_n2175, new_n2176, new_n2177, new_n2178, new_n2179, new_n2180, new_n2181, new_n2182, new_n2183, new_n2184, new_n2185, new_n2186, new_n2187, new_n2188, new_n2189, new_n2190, new_n2191, new_n2192, new_n2193, new_n2194, new_n2195, new_n2196, new_n2197, new_n2198, new_n2199, new_n2200, new_n2201, new_n2202, new_n2203, new_n2204, new_n2205, new_n2206, new_n2207, new_n2208, new_n2209, new_n2210, new_n2211, new_n2212, new_n2213, new_n2214, new_n2215, new_n2216, new_n2217, new_n2218, new_n2219, new_n2220, new_n2221, new_n2222, new_n2223, new_n2224, new_n2225, new_n2226, new_n2227, new_n2228, new_n2229, new_n2230, new_n2231, new_n2232, new_n2233, new_n2234, new_n2235, new_n2236, new_n2237, new_n2238, new_n2239, new_n2240, new_n2241, new_n2242, new_n2243, new_n2244, new_n2245, new_n2246, new_n2247, new_n2248, new_n2249, new_n2250, new_n2251, new_n2252, new_n2253, new_n2254, new_n2255, new_n2256, new_n2257, new_n2258, new_n2259, new_n2260, new_n2261, new_n2262, new_n2263, new_n2264, new_n2265, new_n2266, new_n2267, new_n2268, new_n2269, new_n2270, new_n2271, new_n2272, new_n2273, new_n2274, new_n2275, new_n2276, new_n2277, new_n2278, new_n2279, new_n2280, new_n2281, new_n2282, new_n2283, new_n2284, new_n2285, new_n2286, new_n2287, new_n2288, new_n2289, new_n2290, new_n2291, new_n2292, new_n2293, new_n2294, new_n2295, new_n2296, new_n2297, new_n2298, new_n2299, new_n2300, new_n2301, new_n2302, new_n2303, new_n2304, new_n2305, new_n2306, new_n2307, new_n2308, new_n2309, new_n2310, new_n2311, new_n2312, new_n2313, new_n2314, new_n2315, new_n2316, new_n2317, new_n2318, new_n2319, new_n2320, new_n2321, new_n2322, new_n2323, new_n2324, new_n2325, new_n2326, new_n2327, new_n2328, new_n2329, new_n2330, new_n2331, new_n2332, new_n2333, new_n2334, new_n2335, new_n2336, new_n2337, new_n2338, new_n2339, new_n2340, new_n2341, new_n2342, new_n2343, new_n2344, new_n2345, new_n2346, new_n2347, new_n2348, new_n2349, new_n2350, new_n2351, new_n2352, new_n2353, new_n2354, new_n2355, new_n2356, new_n2357, new_n2358, new_n2359, new_n2360, new_n2361, new_n2362, new_n2363, new_n2364, new_n2365, new_n2366, new_n2367, new_n2368, new_n2369, new_n2370, new_n2371, new_n2372, new_n2373, new_n2374, new_n2375, new_n2376, new_n2377, new_n2378, new_n2379, new_n2380, new_n2381, new_n2382, new_n2383, new_n2384, new_n2385, new_n2386, new_n2387, new_n2388, new_n2389, new_n2390, new_n2391, new_n2392, new_n2393, new_n2394, new_n2395, new_n2396, new_n2397, new_n2398, new_n2399, new_n2400, new_n2401, new_n2402, new_n2403, new_n2404, new_n2405, new_n2406, new_n2407, new_n2408, new_n2409, new_n2410, new_n2411, new_n2412, new_n2413, new_n2414, new_n2415, new_n2416, new_n2417, new_n2418, new_n2419, new_n2420, new_n2421, new_n2422, new_n2423, new_n2424, new_n2425, new_n2426, new_n2427, new_n2428, new_n2429, new_n2430, new_n2431, new_n2432, new_n2433, new_n2434, new_n2435, new_n2436, new_n2437, new_n2438, new_n2439, new_n2440, new_n2441, new_n2442, new_n2443, new_n2444, new_n2445, new_n2446, new_n2447, new_n2448, new_n2449, new_n2450, new_n2451, new_n2452, new_n2453, new_n2454, new_n2455, new_n2456, new_n2457, new_n2458, new_n2459, new_n2460, new_n2461, new_n2462, new_n2463, new_n2464, new_n2465, new_n2466, new_n2467, new_n2468, new_n2469, new_n2470, new_n2471, new_n2472, new_n2473, new_n2474, new_n2475, new_n2476, new_n2477, new_n2478, new_n2479, new_n2480, new_n2481, new_n2482, new_n2483, new_n2484, new_n2485, new_n2486, new_n2487, new_n2488, new_n2489, new_n2490, new_n2491, new_n2492, new_n2493, new_n2494, new_n2495, new_n2496, new_n2497, new_n2498, new_n2499, new_n2500, new_n2501, new_n2502, new_n2503, new_n2504, new_n2505, new_n2506, new_n2507, new_n2508, new_n2509, new_n2510, new_n2511, new_n2512, new_n2513, new_n2514, new_n2515, new_n2516, new_n2517, new_n2518, new_n2519, new_n2520, new_n2521, new_n2522, new_n2523, new_n2524, new_n2525, new_n2526, new_n2527, new_n2528, new_n2529, new_n2530, new_n2531, new_n2532, new_n2533, new_n2534, new_n2535, new_n2536, new_n2537, new_n2538, new_n2539, new_n2540, new_n2541, new_n2542, new_n2543, new_n2544, new_n2545, new_n2546, new_n2547, new_n2548, new_n2549, new_n2550, new_n2551, new_n2552, new_n2553, new_n2554, new_n2555, new_n2556, new_n2557, new_n2558, new_n2559, new_n2560, new_n2561, new_n2562, new_n2563, new_n2564, new_n2565, new_n2566, new_n2567, new_n2568, new_n2569, new_n2570, new_n2571, new_n2572, new_n2573, new_n2574, new_n2575, new_n2576, new_n2577, new_n2578, new_n2579, new_n2580, new_n2581, new_n2582, new_n2583, new_n2584, new_n2585, new_n2586, new_n2587, new_n2588, new_n2589, new_n2590, new_n2591, new_n2592, new_n2593, new_n2594, new_n2595, new_n2596, new_n2597, new_n2598, new_n2599, new_n2600, new_n2601, new_n2602, new_n2603, new_n2604, new_n2605, new_n2606, new_n2607, new_n2608, new_n2609, new_n2610, new_n2611, new_n2612, new_n2613, new_n2614, new_n2615, new_n2616, new_n2617, new_n2618, new_n2619, new_n2620, new_n2621, new_n2622, new_n2623, new_n2624, new_n2625, new_n2626, new_n2627, new_n2628, new_n2629, new_n2630, new_n2631, new_n2632, new_n2633, new_n2634, new_n2635, new_n2636, new_n2637, new_n2638, new_n2639, new_n2640, new_n2641, new_n2642, new_n2643, new_n2644, new_n2645, new_n2646, new_n2647, new_n2648, new_n2649, new_n2650, new_n2651, new_n2652, new_n2653, new_n2654, new_n2655, new_n2656, new_n2657, new_n2658, new_n2659, new_n2660, new_n2661, new_n2662, new_n2663, new_n2664, new_n2665, new_n2666, new_n2667, new_n2668, new_n2669, new_n2670, new_n2671, new_n2672, new_n2673, new_n2674, new_n2675, new_n2676, new_n2677, new_n2678, new_n2679, new_n2680, new_n2681, new_n2682, new_n2683, new_n2684, new_n2685, new_n2686, new_n2687, new_n2688, new_n2689, new_n2690, new_n2691, new_n2692, new_n2693, new_n2694, new_n2695, new_n2696, new_n2697, new_n2698, new_n2699, new_n2700, new_n2701, new_n2702, new_n2703, new_n2704, new_n2705, new_n2706, new_n2707, new_n2708, new_n2709, new_n2710, new_n2711, new_n2712, new_n2713, new_n2714, new_n2715, new_n2716, new_n2717, new_n2718, new_n2719, new_n2720, new_n2721, new_n2722, new_n2723, new_n2724, new_n2725, new_n2726, new_n2727, new_n2728, new_n2729, new_n2730, new_n2731, new_n2732, new_n2733, new_n2734, new_n2735, new_n2736, new_n2737, new_n2738, new_n2739, new_n2740, new_n2741, new_n2742, new_n2743, new_n2744, new_n2745, new_n2746, new_n2747, new_n2748, new_n2749, new_n2750, new_n2751, new_n2752, new_n2753, new_n2754, new_n2755, new_n2756, new_n2757, new_n2758, new_n2759, new_n2760, new_n2761, new_n2762, new_n2763, new_n2764, new_n2765, new_n2766, new_n2767, new_n2768, new_n2769, new_n2770, new_n2771, new_n2772, new_n2773, new_n2774, new_n2775, new_n2776, new_n2777, new_n2778, new_n2779, new_n2780, new_n2781, new_n2782, new_n2783, new_n2784, new_n2785, new_n2786, new_n2787, new_n2788, new_n2789, new_n2790, new_n2791, new_n2792, new_n2793, new_n2794, new_n2795, new_n2796, new_n2797, new_n2798, new_n2799, new_n2800, new_n2801, new_n2802, new_n2803, new_n2804, new_n2805, new_n2806, new_n2807, new_n2808, new_n2809, new_n2810, new_n2811, new_n2812, new_n2813, new_n2814, new_n2815, new_n2816, new_n2817, new_n2818, new_n2819, new_n2820, new_n2821, new_n2822, new_n2823, new_n2824, new_n2825, new_n2826, new_n2827, new_n2828, new_n2829, new_n2830, new_n2831, new_n2832, new_n2833, new_n2834, new_n2835, new_n2836, new_n2837, new_n2838, new_n2839, new_n2840, new_n2841, new_n2842, new_n2843, new_n2844, new_n2845, new_n2846, new_n2847, new_n2848, new_n2849, new_n2850, new_n2851, new_n2852, new_n2853, new_n2854, new_n2855, new_n2856, new_n2857, new_n2858, new_n2859, new_n2860, new_n2861, new_n2862, new_n2863, new_n2864, new_n2865, new_n2866, new_n2867, new_n2868, new_n2869, new_n2870, new_n2871, new_n2872, new_n2873, new_n2874, new_n2875, new_n2876, new_n2877, new_n2878, new_n2879, new_n2880, new_n2881, new_n2882, new_n2883, new_n2884, new_n2885, new_n2886, new_n2887, new_n2888, new_n2889, new_n2890, new_n2891, new_n2892, new_n2893, new_n2894, new_n2895, new_n2896, new_n2897, new_n2898, new_n2899, new_n2900, new_n2901, new_n2902, new_n2903, new_n2904, new_n2905, new_n2906, new_n2907, new_n2908, new_n2909, new_n2910, new_n2911, new_n2912, new_n2913, new_n2914, new_n2915, new_n2916, new_n2917, new_n2918, new_n2919, new_n2920, new_n2921, new_n2922, new_n2923, new_n2924, new_n2925, new_n2926, new_n2927, new_n2928, new_n2929, new_n2930, new_n2931, new_n2932, new_n2933, new_n2934, new_n2935, new_n2936, new_n2937, new_n2938, new_n2939, new_n2940, new_n2941, new_n2942, new_n2943, new_n2944, new_n2945, new_n2946, new_n2947, new_n2948, new_n2949, new_n2950, new_n2951, new_n2952, new_n2953, new_n2954, new_n2955, new_n2956, new_n2957, new_n2958, new_n2959, new_n2960, new_n2961, new_n2962, new_n2963, new_n2964, new_n2965, new_n2966, new_n2967, new_n2968, new_n2969, new_n2970, new_n2971, new_n2972, new_n2973, new_n2974, new_n2975, new_n2976, new_n2977, new_n2978, new_n2979, new_n2980, new_n2981, new_n2982, new_n2983, new_n2984, new_n2985, new_n2986, new_n2987, new_n2988, new_n2989, new_n2990, new_n2991, new_n2992, new_n2993, new_n2994, new_n2995, new_n2996, new_n2997, new_n2998, new_n2999, new_n3000, new_n3001, new_n3002, new_n3003, new_n3004, new_n3005, new_n3006, new_n3007, new_n3008, new_n3009, new_n3010, new_n3011, new_n3012, new_n3013, new_n3014, new_n3015, new_n3016, new_n3017, new_n3018, new_n3019, new_n3020, new_n3021, new_n3022, new_n3023, new_n3024, new_n3025, new_n3026, new_n3027, new_n3028, new_n3029, new_n3030, new_n3031, new_n3032, new_n3033, new_n3034, new_n3035, new_n3036, new_n3037, new_n3038, new_n3039, new_n3040, new_n3041, new_n3042, new_n3043, new_n3044, new_n3045, new_n3046, new_n3047, new_n3048, new_n3049, new_n3050, new_n3051, new_n3052, new_n3053, new_n3054, new_n3055, new_n3056, new_n3057, new_n3058, new_n3059, new_n3060, new_n3061, new_n3062, new_n3063, new_n3064, new_n3065, new_n3066, new_n3067, new_n3068, new_n3069, new_n3070, new_n3071, new_n3072, new_n3073, new_n3074, new_n3075, new_n3076, new_n3077, new_n3078, new_n3079, new_n3080, new_n3081, new_n3082, new_n3083, new_n3084, new_n3085, new_n3086, new_n3087, new_n3088, new_n3089, new_n3090, new_n3091, new_n3092, new_n3093, new_n3094, new_n3095, new_n3096, new_n3097, new_n3098, new_n3099, new_n3100, new_n3101, new_n3102, new_n3103, new_n3104, new_n3105, new_n3106, new_n3107, new_n3108, new_n3109, new_n3110, new_n3111, new_n3112, new_n3113, new_n3114, new_n3115, new_n3116, new_n3117, new_n3118, new_n3119, new_n3120, new_n3121, new_n3122, new_n3123, new_n3124, new_n3125, new_n3126, new_n3127, new_n3128, new_n3129, new_n3130, new_n3131, new_n3132, new_n3133, new_n3134, new_n3135, new_n3136, new_n3137, new_n3138, new_n3139, new_n3140, new_n3141, new_n3142, new_n3143, new_n3144, new_n3145, new_n3146, new_n3147, new_n3148, new_n3149, new_n3150, new_n3151, new_n3152, new_n3153, new_n3154, new_n3155, new_n3156, new_n3157, new_n3158, new_n3159, new_n3160, new_n3161, new_n3162, new_n3163, new_n3164, new_n3165, new_n3166, new_n3167, new_n3168, new_n3169, new_n3170, new_n3171, new_n3172, new_n3173, new_n3174, new_n3175, new_n3176, new_n3177, new_n3178, new_n3179, new_n3180, new_n3181, new_n3182, new_n3183, new_n3184, new_n3185, new_n3186, new_n3187, new_n3188, new_n3189, new_n3190, new_n3191, new_n3192, new_n3193, new_n3194, new_n3195, new_n3196, new_n3197, new_n3198, new_n3199, new_n3200, new_n3201, new_n3202, new_n3203, new_n3204, new_n3205, new_n3206, new_n3207, new_n3208, new_n3209, new_n3210, new_n3211, new_n3212, new_n3213, new_n3214, new_n3215, new_n3216, new_n3217, new_n3218, new_n3219, new_n3220, new_n3221, new_n3222, new_n3223, new_n3224, new_n3225, new_n3226, new_n3227, new_n3228, new_n3229, new_n3230, new_n3231, new_n3232, new_n3233, new_n3234, new_n3235, new_n3236, new_n3237, new_n3238, new_n3239, new_n3240, new_n3241, new_n3242, new_n3243, new_n3244, new_n3245, new_n3246, new_n3247, new_n3248, new_n3249, new_n3250, new_n3251, new_n3252, new_n3253, new_n3254, new_n3255, new_n3256, new_n3257, new_n3258, new_n3259, new_n3260, new_n3261, new_n3262, new_n3263, new_n3264, new_n3265, new_n3266, new_n3267, new_n3268, new_n3269, new_n3270, new_n3271, new_n3272, new_n3273, new_n3274, new_n3275, new_n3276, new_n3277, new_n3278, new_n3279, new_n3280, new_n3281, new_n3282, new_n3283, new_n3284, new_n3285, new_n3286, new_n3287, new_n3288, new_n3289, new_n3290, new_n3291, new_n3292, new_n3293, new_n3294, new_n3295, new_n3296, new_n3297, new_n3298, new_n3299, new_n3300, new_n3301, new_n3302, new_n3303, new_n3304, new_n3305, new_n3306, new_n3307, new_n3308, new_n3309, new_n3310, new_n3311, new_n3312, new_n3313, new_n3314, new_n3315, new_n3316, new_n3317, new_n3318, new_n3319, new_n3320, new_n3321, new_n3322, new_n3323, new_n3324, new_n3325, new_n3326, new_n3327, new_n3328, new_n3329, new_n3330, new_n3331, new_n3332, new_n3333, new_n3334, new_n3335, new_n3336, new_n3337, new_n3338, new_n3339, new_n3340, new_n3341, new_n3342, new_n3343, new_n3344, new_n3345, new_n3346, new_n3347, new_n3348, new_n3349, new_n3350, new_n3351, new_n3352, new_n3353, new_n3354, new_n3355, new_n3356, new_n3357, new_n3358, new_n3359, new_n3360, new_n3361, new_n3362, new_n3363, new_n3364, new_n3365, new_n3366, new_n3367, new_n3368, new_n3369, new_n3370, new_n3371, new_n3372, new_n3373, new_n3374, new_n3375, new_n3376, new_n3377, new_n3378, new_n3379, new_n3380, new_n3381, new_n3382, new_n3383, new_n3384, new_n3385, new_n3386, new_n3387, new_n3388, new_n3389, new_n3390, new_n3391, new_n3392, new_n3393, new_n3394, new_n3395, new_n3396, new_n3397, new_n3398, new_n3399, new_n3400, new_n3401, new_n3402, new_n3403, new_n3404, new_n3405, new_n3406, new_n3407, new_n3408, new_n3409, new_n3410, new_n3411, new_n3412, new_n3413, new_n3414, new_n3415, new_n3416, new_n3417, new_n3418, new_n3419, new_n3420, new_n3421, new_n3422, new_n3423, new_n3424, new_n3425, new_n3426, new_n3427, new_n3428, new_n3429, new_n3430, new_n3431, new_n3432, new_n3433, new_n3434, new_n3435, new_n3436, new_n3437, new_n3438, new_n3439, new_n3440, new_n3441, new_n3442, new_n3443, new_n3444, new_n3445, new_n3446, new_n3447, new_n3448, new_n3449, new_n3450, new_n3451, new_n3452, new_n3453, new_n3454, new_n3455, new_n3456, new_n3457, new_n3458, new_n3459, new_n3460, new_n3461, new_n3462, new_n3463, new_n3464, new_n3465, new_n3466, new_n3467, new_n3468, new_n3469, new_n3470, new_n3471, new_n3472, new_n3473, new_n3474, new_n3475, new_n3476, new_n3477, new_n3478, new_n3479, new_n3480, new_n3481, new_n3482, new_n3483, new_n3484, new_n3485, new_n3486, new_n3487, new_n3488, new_n3489, new_n3490, new_n3491, new_n3492, new_n3493, new_n3494, new_n3495, new_n3496, new_n3497, new_n3498, new_n3499, new_n3500, new_n3501, new_n3502, new_n3503, new_n3504, new_n3505, new_n3506, new_n3507, new_n3508, new_n3509, new_n3510, new_n3511, new_n3512, new_n3513, new_n3514, new_n3515, new_n3516, new_n3517, new_n3518, new_n3519, new_n3520, new_n3521, new_n3522, new_n3523, new_n3524, new_n3525, new_n3526, new_n3527, new_n3528, new_n3529, new_n3530, new_n3531, new_n3532, new_n3533, new_n3534, new_n3535, new_n3536, new_n3537, new_n3538, new_n3539, new_n3540, new_n3541, new_n3542, new_n3543, new_n3544, new_n3545, new_n3546, new_n3547, new_n3548, new_n3549, new_n3550, new_n3551, new_n3552, new_n3553, new_n3554, new_n3555, new_n3556, new_n3557, new_n3558, new_n3559, new_n3560, new_n3561, new_n3562, new_n3563, new_n3564, new_n3565, new_n3566, new_n3567, new_n3568, new_n3569, new_n3570, new_n3571, new_n3572, new_n3573, new_n3574, new_n3575, new_n3576, new_n3577, new_n3578, new_n3579, new_n3580, new_n3581, new_n3582, new_n3583, new_n3584, new_n3585, new_n3586, new_n3587, new_n3588, new_n3589, new_n3590, new_n3591, new_n3592, new_n3593, new_n3594, new_n3595, new_n3596, new_n3597, new_n3598, new_n3599, new_n3600, new_n3601, new_n3602, new_n3603, new_n3604, new_n3605, new_n3606, new_n3607, new_n3608, new_n3609, new_n3610, new_n3611, new_n3612, new_n3613, new_n3614, new_n3615, new_n3616, new_n3617, new_n3618, new_n3619, new_n3620, new_n3621, new_n3622, new_n3623, new_n3624, new_n3625, new_n3626, new_n3627, new_n3628, new_n3629, new_n3630, new_n3631, new_n3632, new_n3633, new_n3634, new_n3635, new_n3636, new_n3637, new_n3638, new_n3639, new_n3640, new_n3641, new_n3642, new_n3643, new_n3644, new_n3645, new_n3646, new_n3647, new_n3648, new_n3649, new_n3650, new_n3651, new_n3652, new_n3653, new_n3654, new_n3655, new_n3656, new_n3657, new_n3658, new_n3659, new_n3660, new_n3661, new_n3662, new_n3663, new_n3664, new_n3665, new_n3666, new_n3667, new_n3668, new_n3669, new_n3670, new_n3671, new_n3672, new_n3673, new_n3674, new_n3675, new_n3676, new_n3677, new_n3678, new_n3679, new_n3680, new_n3681, new_n3682, new_n3683, new_n3684, new_n3685, new_n3686, new_n3687, new_n3688, new_n3689, new_n3690, new_n3691, new_n3692, new_n3693, new_n3694, new_n3695, new_n3696, new_n3697, new_n3698, new_n3699, new_n3700, new_n3701, new_n3702, new_n3703, new_n3704, new_n3705, new_n3706, new_n3707, new_n3708, new_n3709, new_n3710, new_n3711, new_n3712, new_n3713, new_n3714, new_n3715, new_n3716, new_n3717, new_n3718, new_n3719, new_n3720, new_n3721, new_n3722, new_n3723, new_n3724, new_n3725, new_n3726, new_n3727, new_n3728, new_n3729, new_n3730, new_n3731, new_n3732, new_n3733, new_n3734, new_n3735, new_n3736, new_n3737, new_n3738, new_n3739, new_n3740, new_n3741, new_n3742, new_n3743, new_n3744, new_n3745, new_n3746, new_n3747, new_n3748, new_n3749, new_n3750, new_n3751, new_n3752, new_n3753, new_n3754, new_n3755, new_n3756, new_n3757, new_n3758, new_n3759, new_n3760, new_n3761, new_n3762, new_n3763, new_n3764, new_n3765, new_n3766, new_n3767, new_n3768, new_n3769, new_n3770, new_n3771, new_n3772, new_n3773, new_n3774, new_n3775, new_n3776, new_n3777, new_n3778, new_n3779, new_n3780, new_n3781, new_n3782, new_n3783, new_n3784, new_n3785, new_n3786, new_n3787, new_n3788, new_n3789, new_n3790, new_n3791, new_n3792, new_n3793, new_n3794, new_n3795, new_n3796, new_n3797, new_n3798, new_n3799, new_n3800, new_n3801, new_n3802, new_n3803, new_n3804, new_n3805, new_n3806, new_n3807, new_n3808, new_n3809, new_n3810, new_n3811, new_n3812, new_n3813, new_n3814, new_n3815, new_n3816, new_n3817, new_n3818, new_n3819, new_n3820, new_n3821, new_n3822, new_n3823, new_n3824, new_n3825, new_n3826, new_n3827, new_n3828, new_n3829, new_n3830, new_n3831, new_n3832, new_n3833, new_n3834, new_n3835, new_n3836, new_n3837, new_n3838, new_n3839, new_n3840, new_n3841, new_n3842, new_n3843, new_n3844, new_n3845, new_n3846, new_n3847, new_n3848, new_n3849, new_n3850, new_n3851, new_n3852, new_n3853, new_n3854, new_n3855, new_n3856, new_n3857, new_n3858, new_n3859, new_n3860, new_n3861, new_n3862, new_n3863, new_n3864, new_n3865, new_n3866, new_n3867, new_n3868, new_n3869, new_n3870, new_n3871, new_n3872, new_n3873, new_n3874, new_n3875, new_n3876, new_n3877, new_n3878, new_n3879, new_n3880, new_n3881, new_n3882, new_n3883, new_n3884, new_n3885, new_n3886, new_n3887, new_n3888, new_n3889, new_n3890, new_n3891, new_n3892, new_n3893, new_n3894, new_n3895, new_n3896, new_n3897, new_n3898, new_n3899, new_n3900, new_n3901, new_n3902, new_n3903, new_n3904, new_n3905, new_n3906, new_n3907, new_n3908, new_n3909, new_n3910, new_n3911, new_n3912, new_n3913, new_n3914, new_n3915, new_n3916, new_n3917, new_n3918, new_n3919, new_n3920, new_n3921, new_n3922, new_n3923, new_n3924, new_n3925, new_n3926, new_n3927, new_n3928, new_n3929, new_n3930, new_n3931, new_n3932, new_n3933, new_n3934, new_n3935, new_n3936, new_n3937, new_n3938, new_n3939, new_n3940, new_n3941, new_n3942, new_n3943, new_n3944, new_n3945, new_n3946, new_n3947, new_n3948, new_n3949, new_n3950, new_n3951, new_n3952, new_n3953, new_n3954, new_n3955, new_n3956, new_n3957, new_n3958, new_n3959, new_n3960, new_n3961, new_n3962, new_n3963, new_n3964, new_n3965, new_n3966, new_n3967, new_n3968, new_n3969, new_n3970, new_n3971, new_n3972, new_n3973, new_n3974, new_n3975, new_n3976, new_n3977, new_n3978, new_n3979, new_n3980, new_n3981, new_n3982, new_n3983, new_n3984, new_n3985, new_n3986, new_n3987, new_n3988, new_n3989, new_n3990, new_n3991, new_n3992, new_n3993, new_n3994, new_n3995, new_n3996, new_n3997, new_n3998, new_n3999, new_n4000, new_n4001, new_n4002, new_n4003, new_n4004, new_n4005, new_n4006, new_n4007, new_n4008, new_n4009, new_n4010, new_n4011, new_n4012, new_n4013, new_n4014, new_n4015, new_n4016, new_n4017, new_n4018, new_n4019, new_n4020, new_n4021, new_n4022, new_n4023, new_n4024, new_n4025, new_n4026, new_n4027, new_n4028, new_n4029, new_n4030, new_n4031, new_n4032, new_n4033, new_n4034, new_n4035, new_n4036, new_n4037, new_n4038, new_n4039, new_n4040, new_n4041, new_n4042, new_n4043, new_n4044, new_n4045, new_n4046, new_n4047, new_n4048, new_n4049, new_n4050, new_n4051, new_n4052, new_n4053, new_n4054, new_n4055, new_n4056, new_n4057, new_n4058, new_n4059, new_n4060, new_n4061, new_n4062, new_n4063, new_n4064, new_n4065, new_n4066, new_n4067, new_n4068, new_n4069, new_n4070, new_n4071, new_n4072, new_n4073, new_n4074, new_n4075, new_n4076, new_n4077, new_n4078, new_n4079, new_n4080, new_n4081, new_n4082, new_n4083, new_n4084, new_n4085, new_n4086, new_n4087, new_n4088, new_n4089, new_n4090, new_n4091, new_n4092, new_n4093, new_n4094, new_n4095, new_n4096, new_n4097, new_n4098, new_n4099, new_n4100, new_n4101, new_n4102, new_n4103, new_n4104, new_n4105, new_n4106, new_n4107, new_n4108, new_n4109, new_n4110, new_n4111, new_n4112, new_n4113, new_n4114, new_n4115, new_n4116, new_n4117, new_n4118, new_n4119, new_n4120, new_n4121, new_n4122, new_n4123, new_n4124, new_n4125, new_n4126, new_n4127, new_n4128, new_n4129, new_n4130, new_n4131, new_n4132, new_n4133, new_n4134, new_n4135, new_n4136, new_n4137, new_n4138, new_n4139, new_n4140, new_n4141, new_n4142, new_n4143, new_n4144, new_n4145, new_n4146, new_n4147, new_n4148, new_n4149, new_n4150, new_n4151, new_n4152, new_n4153, new_n4154, new_n4155, new_n4156, new_n4157, new_n4158, new_n4159, new_n4160, new_n4161, new_n4162, new_n4163, new_n4164, new_n4165, new_n4166, new_n4167, new_n4168, new_n4169, new_n4170, new_n4171, new_n4172, new_n4173, new_n4174, new_n4175, new_n4176, new_n4177, new_n4178, new_n4179, new_n4180, new_n4181, new_n4182, new_n4183, new_n4184, new_n4185, new_n4186, new_n4187, new_n4188, new_n4189, new_n4190, new_n4191, new_n4192, new_n4193, new_n4194, new_n4195, new_n4196, new_n4197, new_n4198, new_n4199, new_n4200, new_n4201, new_n4202, new_n4203, new_n4204, new_n4205, new_n4206, new_n4207, new_n4208, new_n4209, new_n4210, new_n4211, new_n4212, new_n4213, new_n4214, new_n4215, new_n4216, new_n4217, new_n4218, new_n4219, new_n4220, new_n4221, new_n4222, new_n4223, new_n4224, new_n4225, new_n4226, new_n4227, new_n4228, new_n4229, new_n4230, new_n4231, new_n4232, new_n4233, new_n4234, new_n4235, new_n4236, new_n4237, new_n4238, new_n4239, new_n4240, new_n4241, new_n4242, new_n4243, new_n4244, new_n4245, new_n4246, new_n4247, new_n4248, new_n4249, new_n4250, new_n4251, new_n4252, new_n4253, new_n4254, new_n4255, new_n4256, new_n4257, new_n4258, new_n4259, new_n4260, new_n4261, new_n4262, new_n4263, new_n4264, new_n4265, new_n4266, new_n4267, new_n4268, new_n4269, new_n4270, new_n4271, new_n4272, new_n4273, new_n4274, new_n4275, new_n4276, new_n4277, new_n4278, new_n4279, new_n4280, new_n4281, new_n4282, new_n4283, new_n4284, new_n4285, new_n4286, new_n4287, new_n4288, new_n4289, new_n4290, new_n4291, new_n4292, new_n4293, new_n4294, new_n4295, new_n4296, new_n4297, new_n4298, new_n4299, new_n4300, new_n4301, new_n4302, new_n4303, new_n4304, new_n4305, new_n4306, new_n4307, new_n4308, new_n4309, new_n4310, new_n4311, new_n4312, new_n4313, new_n4314, new_n4315, new_n4316, new_n4317, new_n4318, new_n4319, new_n4320, new_n4321, new_n4322, new_n4323, new_n4324, new_n4325, new_n4326, new_n4327, new_n4328, new_n4329, new_n4330, new_n4331, new_n4332, new_n4333, new_n4334, new_n4335, new_n4336, new_n4337, new_n4338, new_n4339, new_n4340, new_n4341, new_n4342, new_n4343, new_n4344, new_n4345, new_n4346, new_n4347, new_n4348, new_n4349, new_n4350, new_n4351, new_n4352, new_n4353, new_n4354, new_n4355, new_n4356, new_n4357, new_n4358, new_n4359, new_n4360, new_n4361, new_n4362, new_n4363, new_n4364, new_n4365, new_n4366, new_n4367, new_n4368, new_n4369, new_n4370, new_n4371, new_n4372, new_n4373, new_n4374, new_n4375, new_n4376, new_n4377, new_n4378, new_n4379, new_n4380, new_n4381, new_n4382, new_n4383, new_n4384, new_n4385, new_n4386, new_n4387, new_n4388, new_n4389, new_n4390, new_n4391, new_n4392, new_n4393, new_n4394, new_n4395, new_n4396, new_n4397, new_n4398, new_n4399, new_n4400, new_n4401, new_n4402, new_n4403, new_n4404, new_n4405, new_n4406, new_n4407, new_n4408, new_n4409, new_n4410, new_n4411, new_n4412, new_n4413, new_n4414, new_n4415, new_n4416, new_n4417, new_n4418, new_n4419, new_n4420, new_n4421, new_n4422, new_n4423, new_n4424, new_n4425, new_n4426, new_n4427, new_n4428, new_n4429, new_n4430, new_n4431, new_n4432, new_n4433, new_n4434, new_n4435, new_n4436, new_n4437, new_n4438, new_n4439, new_n4440, new_n4441, new_n4442, new_n4443, new_n4444, new_n4445, new_n4446, new_n4447, new_n4448, new_n4449, new_n4450, new_n4451, new_n4452, new_n4453, new_n4454, new_n4455, new_n4456, new_n4457, new_n4458, new_n4459, new_n4460, new_n4461, new_n4462, new_n4463, new_n4464, new_n4465, new_n4466, new_n4467, new_n4468, new_n4469, new_n4470, new_n4471, new_n4472, new_n4473, new_n4474, new_n4475, new_n4476, new_n4477, new_n4478, new_n4479, new_n4480, new_n4481, new_n4482, new_n4483, new_n4484, new_n4485, new_n4486, new_n4487, new_n4488, new_n4489, new_n4490, new_n4491, new_n4492, new_n4493, new_n4494, new_n4495, new_n4496, new_n4497, new_n4498, new_n4499, new_n4500, new_n4501, new_n4502, new_n4503, new_n4504, new_n4505, new_n4506, new_n4507, new_n4508, new_n4509, new_n4510, new_n4511, new_n4512, new_n4513, new_n4514, new_n4515, new_n4516, new_n4517, new_n4518, new_n4519, new_n4520, new_n4521, new_n4522, new_n4523, new_n4524, new_n4525, new_n4526, new_n4527, new_n4528, new_n4529, new_n4530, new_n4531, new_n4532, new_n4533, new_n4534, new_n4535, new_n4536, new_n4537, new_n4538, new_n4539, new_n4540, new_n4541, new_n4542, new_n4543, new_n4544, new_n4545, new_n4546, new_n4547, new_n4548, new_n4549, new_n4550, new_n4551, new_n4552, new_n4553, new_n4554, new_n4555, new_n4556, new_n4557, new_n4558, new_n4559, new_n4560, new_n4561, new_n4562, new_n4563, new_n4564, new_n4565, new_n4566, new_n4567, new_n4568, new_n4569, new_n4570, new_n4571, new_n4572, new_n4573, new_n4574, new_n4575, new_n4576, new_n4577, new_n4578, new_n4579, new_n4580, new_n4581, new_n4582, new_n4583, new_n4584, new_n4585, new_n4586, new_n4587, new_n4588, new_n4589, new_n4590, new_n4591, new_n4592, new_n4593, new_n4594, new_n4595, new_n4596, new_n4597, new_n4598, new_n4599, new_n4600, new_n4601, new_n4602, new_n4603, new_n4604, new_n4605, new_n4606, new_n4607, new_n4608, new_n4609, new_n4610, new_n4611, new_n4612, new_n4613, new_n4614, new_n4615, new_n4616, new_n4617, new_n4618, new_n4619, new_n4620, new_n4621, new_n4622, new_n4623, new_n4624, new_n4625, new_n4626, new_n4627, new_n4628, new_n4629, new_n4630, new_n4631, new_n4632, new_n4633, new_n4634, new_n4635, new_n4636, new_n4637, new_n4638, new_n4639, new_n4640, new_n4641, new_n4642, new_n4643, new_n4644, new_n4645, new_n4646, new_n4647, new_n4648, new_n4649, new_n4650, new_n4651, new_n4652, new_n4653, new_n4654, new_n4655, new_n4656, new_n4657, new_n4658, new_n4659, new_n4660, new_n4661, new_n4662, new_n4663, new_n4664, new_n4665, new_n4666, new_n4667, new_n4668, new_n4669, new_n4670, new_n4671, new_n4672, new_n4673, new_n4674, new_n4675, new_n4676, new_n4677, new_n4678, new_n4679, new_n4680, new_n4681, new_n4682, new_n4683, new_n4684, new_n4685, new_n4686, new_n4687, new_n4688, new_n4689, new_n4690, new_n4691, new_n4692, new_n4693, new_n4694, new_n4695, new_n4696, new_n4697, new_n4698, new_n4699, new_n4700, new_n4701, new_n4702, new_n4703, new_n4704, new_n4705, new_n4706, new_n4707, new_n4708, new_n4709, new_n4710, new_n4711, new_n4712, new_n4713, new_n4714, new_n4715, new_n4716, new_n4717, new_n4718, new_n4719, new_n4720, new_n4721, new_n4722, new_n4723, new_n4724, new_n4725, new_n4726, new_n4727, new_n4728, new_n4729, new_n4730, new_n4731, new_n4732, new_n4733, new_n4734, new_n4735, new_n4736, new_n4737, new_n4738, new_n4739, new_n4740, new_n4741, new_n4742, new_n4743, new_n4744, new_n4745, new_n4746, new_n4747, new_n4748, new_n4749, new_n4750, new_n4751, new_n4752, new_n4753, new_n4754, new_n4755, new_n4756, new_n4757, new_n4758, new_n4759, new_n4760, new_n4761, new_n4762, new_n4763, new_n4764, new_n4765, new_n4766, new_n4767, new_n4768, new_n4769, new_n4770, new_n4771, new_n4772, new_n4773, new_n4774, new_n4775, new_n4776, new_n4777, new_n4778, new_n4779, new_n4780, new_n4781, new_n4782, new_n4783, new_n4784, new_n4785, new_n4786, new_n4787, new_n4788, new_n4789, new_n4790, new_n4791, new_n4792, new_n4793, new_n4794, new_n4795, new_n4796, new_n4797, new_n4798, new_n4799, new_n4800, new_n4801, new_n4802, new_n4803, new_n4804, new_n4805, new_n4806, new_n4807, new_n4808, new_n4809, new_n4810, new_n4811, new_n4812, new_n4813, new_n4814, new_n4815, new_n4816, new_n4817, new_n4818, new_n4819, new_n4820, new_n4821, new_n4822, new_n4823, new_n4824, new_n4825, new_n4826, new_n4827, new_n4828, new_n4829, new_n4830, new_n4831, new_n4832, new_n4833, new_n4834, new_n4835, new_n4836, new_n4837, new_n4838, new_n4839, new_n4840, new_n4841, new_n4842, new_n4843, new_n4844, new_n4845, new_n4846, new_n4847, new_n4848, new_n4849, new_n4850, new_n4851, new_n4852, new_n4853, new_n4854, new_n4855, new_n4856, new_n4857, new_n4858, new_n4859, new_n4860, new_n4861, new_n4862, new_n4863, new_n4864, new_n4865, new_n4866, new_n4867, new_n4868, new_n4869, new_n4870, new_n4871, new_n4872, new_n4873, new_n4874, new_n4875, new_n4876, new_n4877, new_n4878, new_n4879, new_n4880, new_n4881, new_n4882, new_n4883, new_n4884, new_n4885, new_n4886, new_n4887, new_n4888, new_n4889, new_n4890, new_n4891, new_n4892, new_n4893, new_n4894, new_n4895, new_n4896, new_n4897, new_n4898, new_n4899, new_n4900, new_n4901, new_n4902, new_n4903, new_n4904, new_n4905, new_n4906, new_n4907, new_n4908, new_n4909, new_n4910, new_n4911, new_n4912, new_n4913, new_n4914, new_n4915, new_n4916, new_n4917, new_n4918, new_n4919, new_n4920, new_n4921, new_n4922, new_n4923, new_n4924, new_n4925, new_n4926, new_n4927, new_n4928, new_n4929, new_n4930, new_n4931, new_n4932, new_n4933, new_n4934, new_n4935, new_n4936, new_n4937, new_n4938, new_n4939, new_n4940, new_n4941, new_n4942, new_n4943, new_n4944, new_n4945, new_n4946, new_n4947, new_n4948, new_n4949, new_n4950, new_n4951, new_n4952, new_n4953, new_n4954, new_n4955, new_n4956, new_n4957, new_n4958, new_n4959, new_n4960, new_n4961, new_n4962, new_n4963, new_n4964, new_n4965, new_n4966, new_n4967, new_n4968, new_n4969, new_n4970, new_n4971, new_n4972, new_n4973, new_n4974, new_n4975, new_n4976, new_n4977, new_n4978, new_n4979, new_n4980, new_n4981, new_n4982, new_n4983, new_n4984, new_n4985, new_n4986, new_n4987, new_n4988, new_n4989, new_n4990, new_n4991, new_n4992, new_n4993, new_n4994, new_n4995, new_n4996, new_n4997, new_n4998, new_n4999, new_n5000, new_n5001, new_n5002, new_n5003, new_n5004, new_n5005, new_n5006, new_n5007, new_n5008, new_n5009, new_n5010, new_n5011, new_n5012, new_n5013, new_n5014, new_n5015, new_n5016, new_n5017, new_n5018, new_n5019, new_n5020, new_n5021, new_n5022, new_n5023, new_n5024, new_n5025, new_n5026, new_n5027, new_n5028, new_n5029, new_n5030, new_n5031, new_n5032, new_n5033, new_n5034, new_n5035, new_n5036, new_n5037, new_n5038, new_n5039, new_n5040, new_n5041, new_n5042, new_n5043, new_n5044, new_n5045, new_n5046, new_n5047, new_n5048, new_n5049, new_n5050, new_n5051, new_n5052, new_n5053, new_n5054, new_n5055, new_n5056, new_n5057, new_n5058, new_n5059, new_n5060, new_n5061, new_n5062, new_n5063, new_n5064, new_n5065, new_n5066, new_n5067, new_n5068, new_n5069, new_n5070, new_n5071, new_n5072, new_n5073, new_n5074, new_n5075, new_n5076, new_n5077, new_n5078, new_n5079, new_n5080, new_n5081, new_n5082, new_n5083, new_n5084, new_n5085, new_n5086, new_n5087, new_n5088, new_n5089, new_n5090, new_n5091, new_n5092, new_n5093, new_n5094, new_n5095, new_n5096, new_n5097, new_n5098, new_n5099, new_n5100, new_n5101, new_n5102, new_n5103, new_n5104, new_n5105, new_n5106, new_n5107, new_n5108, new_n5109, new_n5110, new_n5111, new_n5112, new_n5113, new_n5114, new_n5115, new_n5116, new_n5117, new_n5118, new_n5119, new_n5120, new_n5121, new_n5122, new_n5123, new_n5124, new_n5125, new_n5126, new_n5127, new_n5128, new_n5129, new_n5130, new_n5131, new_n5132, new_n5133, new_n5134, new_n5135, new_n5136, new_n5137, new_n5138, new_n5139, new_n5140, new_n5141, new_n5142, new_n5143, new_n5144, new_n5145, new_n5146, new_n5147, new_n5148, new_n5149, new_n5150, new_n5151, new_n5152, new_n5153, new_n5154, new_n5155, new_n5156, new_n5157, new_n5158, new_n5159, new_n5160, new_n5161, new_n5162, new_n5163, new_n5164, new_n5165, new_n5166, new_n5167, new_n5168, new_n5169, new_n5170, new_n5171, new_n5172, new_n5173, new_n5174, new_n5175, new_n5176, new_n5177, new_n5178, new_n5179, new_n5180, new_n5181, new_n5182, new_n5183, new_n5184, new_n5185, new_n5186, new_n5187, new_n5188, new_n5189, new_n5190, new_n5191, new_n5192, new_n5193, new_n5194, new_n5195, new_n5196, new_n5197, new_n5198, new_n5199, new_n5200, new_n5201, new_n5202, new_n5203, new_n5204, new_n5205, new_n5206, new_n5207, new_n5208, new_n5209, new_n5210, new_n5211, new_n5212, new_n5213, new_n5214, new_n5215, new_n5216, new_n5217, new_n5218, new_n5219, new_n5220, new_n5221, new_n5222, new_n5223, new_n5224, new_n5225, new_n5226, new_n5227, new_n5228, new_n5229, new_n5230, new_n5231, new_n5232, new_n5233, new_n5234, new_n5235, new_n5236, new_n5237, new_n5238, new_n5239, new_n5240, new_n5241, new_n5242, new_n5243, new_n5244, new_n5245, new_n5246, new_n5247, new_n5248, new_n5249, new_n5250, new_n5251, new_n5252, new_n5253, new_n5254, new_n5255, new_n5256, new_n5257, new_n5258, new_n5259, new_n5260, new_n5261, new_n5262, new_n5263, new_n5264, new_n5265, new_n5266, new_n5267, new_n5268, new_n5269, new_n5270, new_n5271, new_n5272, new_n5273, new_n5274, new_n5275, new_n5276, new_n5277, new_n5278, new_n5279, new_n5280, new_n5281, new_n5282, new_n5283, new_n5284, new_n5285, new_n5286, new_n5287, new_n5288, new_n5289, new_n5290, new_n5291, new_n5292, new_n5293, new_n5294, new_n5295, new_n5296, new_n5297, new_n5298, new_n5299, new_n5300, new_n5301, new_n5302, new_n5303, new_n5304, new_n5305, new_n5306, new_n5307, new_n5308, new_n5309, new_n5310, new_n5311, new_n5312, new_n5313, new_n5314, new_n5315, new_n5316, new_n5317, new_n5318, new_n5319, new_n5320, new_n5321, new_n5322, new_n5323, new_n5324, new_n5325, new_n5326, new_n5327, new_n5328, new_n5329, new_n5330, new_n5331, new_n5332, new_n5333, new_n5334, new_n5335, new_n5336, new_n5337, new_n5338, new_n5339, new_n5340, new_n5341, new_n5342, new_n5343, new_n5344, new_n5345, new_n5346, new_n5347, new_n5348, new_n5349, new_n5350, new_n5351, new_n5352, new_n5353, new_n5354, new_n5355, new_n5356, new_n5357, new_n5358, new_n5359, new_n5360, new_n5361, new_n5362, new_n5363, new_n5364, new_n5365, new_n5366, new_n5367, new_n5368, new_n5369, new_n5370, new_n5371, new_n5372, new_n5373, new_n5374, new_n5375, new_n5376, new_n5377, new_n5378, new_n5379, new_n5380, new_n5381, new_n5382, new_n5383, new_n5384, new_n5385, new_n5386, new_n5387, new_n5388, new_n5389, new_n5390, new_n5391, new_n5392, new_n5393, new_n5394, new_n5395, new_n5396, new_n5397, new_n5398, new_n5399, new_n5400, new_n5401, new_n5402, new_n5403, new_n5404, new_n5405, new_n5406, new_n5407, new_n5408, new_n5409, new_n5410, new_n5411, new_n5412, new_n5413, new_n5414, new_n5415, new_n5416, new_n5417, new_n5418, new_n5419, new_n5420, new_n5421, new_n5422, new_n5423, new_n5424, new_n5425, new_n5426, new_n5427, new_n5428, new_n5429, new_n5430, new_n5431, new_n5432, new_n5433, new_n5434, new_n5435, new_n5436, new_n5437, new_n5438, new_n5439, new_n5440, new_n5441, new_n5442, new_n5443, new_n5444, new_n5445, new_n5446, new_n5447, new_n5448, new_n5449, new_n5450, new_n5451, new_n5452, new_n5453, new_n5454, new_n5455, new_n5456, new_n5457, new_n5458, new_n5459, new_n5460, new_n5461, new_n5462, new_n5463, new_n5464, new_n5465, new_n5466, new_n5467, new_n5468, new_n5469, new_n5470, new_n5471, new_n5472, new_n5473, new_n5474, new_n5475, new_n5476, new_n5477, new_n5478, new_n5479, new_n5480, new_n5481, new_n5482, new_n5483, new_n5484, new_n5485, new_n5486, new_n5487, new_n5488, new_n5489, new_n5490, new_n5491, new_n5492, new_n5493, new_n5494, new_n5495, new_n5496, new_n5497, new_n5498, new_n5499, new_n5500, new_n5501, new_n5502, new_n5503, new_n5504, new_n5505, new_n5506, new_n5507, new_n5508, new_n5509, new_n5510, new_n5511, new_n5512, new_n5513, new_n5514, new_n5515, new_n5516, new_n5517, new_n5518, new_n5519, new_n5520, new_n5521, new_n5522, new_n5523, new_n5524, new_n5525, new_n5526, new_n5527, new_n5528, new_n5529, new_n5530, new_n5531, new_n5532, new_n5533, new_n5534, new_n5535, new_n5536, new_n5537, new_n5538, new_n5539, new_n5540, new_n5541, new_n5542, new_n5543, new_n5544, new_n5545, new_n5546, new_n5547, new_n5548, new_n5549, new_n5550, new_n5551, new_n5552, new_n5553, new_n5554, new_n5555, new_n5556, new_n5557, new_n5558, new_n5559, new_n5560, new_n5561, new_n5562, new_n5563, new_n5564, new_n5565, new_n5566, new_n5567, new_n5568, new_n5569, new_n5570, new_n5571, new_n5572, new_n5573, new_n5574, new_n5575, new_n5576, new_n5577, new_n5578, new_n5579, new_n5580, new_n5581, new_n5582, new_n5583, new_n5584, new_n5585, new_n5586, new_n5587, new_n5588, new_n5589, new_n5590, new_n5591, new_n5592, new_n5593, new_n5594, new_n5595, new_n5596, new_n5597, new_n5598, new_n5599, new_n5600, new_n5601, new_n5602, new_n5603, new_n5604, new_n5605, new_n5606, new_n5607, new_n5608, new_n5609, new_n5610, new_n5611, new_n5612, new_n5613, new_n5614, new_n5615, new_n5616, new_n5617, new_n5618, new_n5619, new_n5620, new_n5621, new_n5622, new_n5623, new_n5624, new_n5625, new_n5626, new_n5627, new_n5628, new_n5629, new_n5630, new_n5631, new_n5632, new_n5633, new_n5634, new_n5635, new_n5636, new_n5637, new_n5638, new_n5639, new_n5640, new_n5641, new_n5642, new_n5643, new_n5644, new_n5645, new_n5646, new_n5647, new_n5648, new_n5649, new_n5650, new_n5651, new_n5652, new_n5653, new_n5654, new_n5655, new_n5656, new_n5657, new_n5658, new_n5659, new_n5660, new_n5661, new_n5662, new_n5663, new_n5664, new_n5665, new_n5666, new_n5667, new_n5668, new_n5669, new_n5670, new_n5671, new_n5672, new_n5673, new_n5674, new_n5675, new_n5676, new_n5677, new_n5678, new_n5679, new_n5680, new_n5681, new_n5682, new_n5683, new_n5684, new_n5685, new_n5686, new_n5687, new_n5688, new_n5689, new_n5690, new_n5691, new_n5692, new_n5693, new_n5694, new_n5695, new_n5696, new_n5697, new_n5698, new_n5699, new_n5700, new_n5701, new_n5702, new_n5703, new_n5704, new_n5705, new_n5706, new_n5707, new_n5708, new_n5709, new_n5710, new_n5711, new_n5712, new_n5713, new_n5714, new_n5715, new_n5716, new_n5717, new_n5718, new_n5719, new_n5720, new_n5721, new_n5722, new_n5723, new_n5724, new_n5725, new_n5726, new_n5727, new_n5728, new_n5729, new_n5730, new_n5731, new_n5732, new_n5733, new_n5734, new_n5735, new_n5736, new_n5737, new_n5738, new_n5739, new_n5740, new_n5741, new_n5742, new_n5743, new_n5744, new_n5745, new_n5746, new_n5747, new_n5748, new_n5749, new_n5750, new_n5751, new_n5752, new_n5753, new_n5754, new_n5755, new_n5756, new_n5757, new_n5758, new_n5759, new_n5760, new_n5761, new_n5762, new_n5763, new_n5764, new_n5765, new_n5766, new_n5767, new_n5768, new_n5769, new_n5770, new_n5771, new_n5772, new_n5773, new_n5774, new_n5775, new_n5776, new_n5777, new_n5778, new_n5779, new_n5780, new_n5781, new_n5782, new_n5783, new_n5784, new_n5785, new_n5786, new_n5787, new_n5788, new_n5789, new_n5790, new_n5791, new_n5792, new_n5793, new_n5794, new_n5795, new_n5796, new_n5797, new_n5798, new_n5799, new_n5800, new_n5801, new_n5802, new_n5803, new_n5804, new_n5805, new_n5806, new_n5807, new_n5808, new_n5809, new_n5810, new_n5811, new_n5812, new_n5813, new_n5814, new_n5815, new_n5816, new_n5817, new_n5818, new_n5819, new_n5820, new_n5821, new_n5822, new_n5823, new_n5824, new_n5825, new_n5826, new_n5827, new_n5828, new_n5829, new_n5830, new_n5831, new_n5832, new_n5833, new_n5834, new_n5835, new_n5836, new_n5837, new_n5838, new_n5839, new_n5840, new_n5841, new_n5842, new_n5843, new_n5844, new_n5845, new_n5846, new_n5847, new_n5848, new_n5849, new_n5850, new_n5851, new_n5852, new_n5853, new_n5854, new_n5855, new_n5856, new_n5857, new_n5858, new_n5859, new_n5860, new_n5861, new_n5862, new_n5863, new_n5864, new_n5865, new_n5866, new_n5867, new_n5868, new_n5869, new_n5870, new_n5871, new_n5872, new_n5873, new_n5874, new_n5875, new_n5876, new_n5877, new_n5878, new_n5879, new_n5880, new_n5881, new_n5882, new_n5883, new_n5884, new_n5885, new_n5886, new_n5887, new_n5888, new_n5889, new_n5890, new_n5891, new_n5892, new_n5893, new_n5894, new_n5895, new_n5896, new_n5897, new_n5898, new_n5899, new_n5900, new_n5901, new_n5902, new_n5903, new_n5904, new_n5905, new_n5906, new_n5907, new_n5908, new_n5909, new_n5910, new_n5911, new_n5912, new_n5913, new_n5914, new_n5915, new_n5916, new_n5917, new_n5918, new_n5919, new_n5920, new_n5921, new_n5922, new_n5923, new_n5924, new_n5925, new_n5926, new_n5927, new_n5928, new_n5929, new_n5930, new_n5931, new_n5932, new_n5933, new_n5934, new_n5935, new_n5936, new_n5937, new_n5938, new_n5939, new_n5940, new_n5941, new_n5942, new_n5943, new_n5944, new_n5945, new_n5946, new_n5947, new_n5948, new_n5949, new_n5950, new_n5951, new_n5952, new_n5953, new_n5954, new_n5955, new_n5956, new_n5957, new_n5958, new_n5959, new_n5960, new_n5961, new_n5962, new_n5963, new_n5964, new_n5965, new_n5966, new_n5967, new_n5968, new_n5969, new_n5970, new_n5971, new_n5972, new_n5973, new_n5974, new_n5975, new_n5976, new_n5977, new_n5978, new_n5979, new_n5980, new_n5981, new_n5982, new_n5983, new_n5984, new_n5985, new_n5986, new_n5987, new_n5988, new_n5989, new_n5990, new_n5991, new_n5992, new_n5993, new_n5994, new_n5995, new_n5996, new_n5997, new_n5998, new_n5999, new_n6000, new_n6001, new_n6002, new_n6003, new_n6004, new_n6005, new_n6006, new_n6007, new_n6008, new_n6009, new_n6010, new_n6011, new_n6012, new_n6013, new_n6014, new_n6015, new_n6016, new_n6017, new_n6018, new_n6019, new_n6020, new_n6021, new_n6022, new_n6023, new_n6024, new_n6025, new_n6026, new_n6027, new_n6028, new_n6029, new_n6030, new_n6031, new_n6032, new_n6033, new_n6034, new_n6035, new_n6036, new_n6037, new_n6038, new_n6039, new_n6040, new_n6041, new_n6042, new_n6043, new_n6044, new_n6045, new_n6046, new_n6047, new_n6048, new_n6049, new_n6050, new_n6051, new_n6052, new_n6053, new_n6054, new_n6055, new_n6056, new_n6057, new_n6058, new_n6059, new_n6060, new_n6061, new_n6062, new_n6063, new_n6064, new_n6065, new_n6066, new_n6067, new_n6068, new_n6069, new_n6070, new_n6071, new_n6072, new_n6073, new_n6074, new_n6075, new_n6076, new_n6077, new_n6078, new_n6079, new_n6080, new_n6081, new_n6082, new_n6083, new_n6084, new_n6085, new_n6086, new_n6087, new_n6088, new_n6089, new_n6090, new_n6091, new_n6092, new_n6093, new_n6094, new_n6095, new_n6096, new_n6097, new_n6098, new_n6099, new_n6100, new_n6101, new_n6102, new_n6103, new_n6104, new_n6105, new_n6106, new_n6107, new_n6108, new_n6109, new_n6110, new_n6111, new_n6112, new_n6113, new_n6114, new_n6115, new_n6116, new_n6117, new_n6118, new_n6119, new_n6120, new_n6121, new_n6122, new_n6123, new_n6124, new_n6125, new_n6126, new_n6127, new_n6128, new_n6129, new_n6130, new_n6131, new_n6132, new_n6133, new_n6134, new_n6135, new_n6136, new_n6137, new_n6138, new_n6139, new_n6140, new_n6141, new_n6142, new_n6143, new_n6144, new_n6145, new_n6146, new_n6147, new_n6148, new_n6149, new_n6150, new_n6151, new_n6152, new_n6153, new_n6154, new_n6155, new_n6156, new_n6157, new_n6158, new_n6159, new_n6160, new_n6161, new_n6162, new_n6163, new_n6164, new_n6165, new_n6166, new_n6167, new_n6168, new_n6169, new_n6170, new_n6171, new_n6172, new_n6173, new_n6174, new_n6175, new_n6176, new_n6177, new_n6178, new_n6179, new_n6180, new_n6181, new_n6182, new_n6183, new_n6184, new_n6185, new_n6186, new_n6187, new_n6188, new_n6189, new_n6190, new_n6191, new_n6192, new_n6193, new_n6194, new_n6195, new_n6196, new_n6197, new_n6198, new_n6199, new_n6200, new_n6201, new_n6202, new_n6203, new_n6204, new_n6205, new_n6206, new_n6207, new_n6208, new_n6209, new_n6210, new_n6211, new_n6212, new_n6213, new_n6214, new_n6215, new_n6216, new_n6217, new_n6218, new_n6219, new_n6220, new_n6221, new_n6222, new_n6223, new_n6224, new_n6225, new_n6226, new_n6227, new_n6228, new_n6229, new_n6230, new_n6231, new_n6232, new_n6233, new_n6234, new_n6235, new_n6236, new_n6237, new_n6238, new_n6239, new_n6240, new_n6241, new_n6242, new_n6243, new_n6244, new_n6245, new_n6246, new_n6247, new_n6248, new_n6249, new_n6250, new_n6251, new_n6252, new_n6253, new_n6254, new_n6255, new_n6256, new_n6257, new_n6258, new_n6259, new_n6260, new_n6261, new_n6262, new_n6263, new_n6264, new_n6265, new_n6266, new_n6267, new_n6268, new_n6269, new_n6270, new_n6271, new_n6272, new_n6273, new_n6274, new_n6275, new_n6276, new_n6277, new_n6278, new_n6279, new_n6280, new_n6281, new_n6282, new_n6283, new_n6284, new_n6285, new_n6286, new_n6287, new_n6288, new_n6289, new_n6290, new_n6291, new_n6292, new_n6293, new_n6294, new_n6295, new_n6296, new_n6297, new_n6298, new_n6299, new_n6300, new_n6301, new_n6302, new_n6303, new_n6304, new_n6305, new_n6306, new_n6307, new_n6308, new_n6309, new_n6310, new_n6311, new_n6312, new_n6313, new_n6314, new_n6315, new_n6316, new_n6317, new_n6318, new_n6319, new_n6320, new_n6321, new_n6322, new_n6323, new_n6324, new_n6325, new_n6326, new_n6327, new_n6328, new_n6329, new_n6330, new_n6331, new_n6332, new_n6333, new_n6334, new_n6335, new_n6336, new_n6337, new_n6338, new_n6339, new_n6340, new_n6341, new_n6342, new_n6343, new_n6344, new_n6345, new_n6346, new_n6347, new_n6348, new_n6349, new_n6350, new_n6351, new_n6352, new_n6353, new_n6354, new_n6355, new_n6356, new_n6357, new_n6358, new_n6359, new_n6360, new_n6361, new_n6362, new_n6363, new_n6364, new_n6365, new_n6366, new_n6367, new_n6368, new_n6369, new_n6370, new_n6371, new_n6372, new_n6373, new_n6374, new_n6375, new_n6376, new_n6377, new_n6378, new_n6379, new_n6380, new_n6381, new_n6382, new_n6383, new_n6384, new_n6385, new_n6386, new_n6387, new_n6388, new_n6389, new_n6390, new_n6391, new_n6392, new_n6393, new_n6394, new_n6395, new_n6396, new_n6397, new_n6398, new_n6399, new_n6400, new_n6401, new_n6402, new_n6403, new_n6404, new_n6405, new_n6406, new_n6407, new_n6408, new_n6409, new_n6410, new_n6411, new_n6412, new_n6413, new_n6414, new_n6415, new_n6416, new_n6417, new_n6418, new_n6419, new_n6420, new_n6421, new_n6422, new_n6423, new_n6424, new_n6425, new_n6426, new_n6427, new_n6428, new_n6429, new_n6430, new_n6431, new_n6432, new_n6433, new_n6434, new_n6435, new_n6436, new_n6437, new_n6438, new_n6439, new_n6440, new_n6441, new_n6442, new_n6443, new_n6444, new_n6445, new_n6446, new_n6447, new_n6448, new_n6449, new_n6450, new_n6451, new_n6452, new_n6453, new_n6454, new_n6455, new_n6456, new_n6457, new_n6458, new_n6459, new_n6460, new_n6461, new_n6462, new_n6463, new_n6464, new_n6465, new_n6466, new_n6467, new_n6468, new_n6469, new_n6470, new_n6471, new_n6472, new_n6473, new_n6474, new_n6475, new_n6476, new_n6477, new_n6478, new_n6479, new_n6480, new_n6481, new_n6482, new_n6483, new_n6484, new_n6485, new_n6486, new_n6487, new_n6488, new_n6489, new_n6490, new_n6491, new_n6492, new_n6493, new_n6494, new_n6495, new_n6496, new_n6497, new_n6498, new_n6499, new_n6500, new_n6501, new_n6502, new_n6503, new_n6504, new_n6505, new_n6506, new_n6507, new_n6508, new_n6509, new_n6510, new_n6511, new_n6512, new_n6513, new_n6514, new_n6515, new_n6516, new_n6517, new_n6518, new_n6519, new_n6520, new_n6521, new_n6522, new_n6523, new_n6524, new_n6525, new_n6526, new_n6527, new_n6528, new_n6529, new_n6530, new_n6531, new_n6532, new_n6533, new_n6534, new_n6535, new_n6536, new_n6537, new_n6538, new_n6539, new_n6540, new_n6541, new_n6542, new_n6543, new_n6544, new_n6545, new_n6546, new_n6547, new_n6548, new_n6549, new_n6550, new_n6551, new_n6552, new_n6553, new_n6554, new_n6555, new_n6556, new_n6557, new_n6558, new_n6559, new_n6560, new_n6561, new_n6562, new_n6563, new_n6564, new_n6565, new_n6566, new_n6567, new_n6568, new_n6569, new_n6570, new_n6571, new_n6572, new_n6573, new_n6574, new_n6575, new_n6576, new_n6577, new_n6578, new_n6579, new_n6580, new_n6581, new_n6582, new_n6583, new_n6584, new_n6585, new_n6586, new_n6587, new_n6588, new_n6589, new_n6590, new_n6591, new_n6592, new_n6593, new_n6594, new_n6595, new_n6596, new_n6597, new_n6598, new_n6599, new_n6600, new_n6601, new_n6602, new_n6603, new_n6604, new_n6605, new_n6606, new_n6607, new_n6608, new_n6609, new_n6610, new_n6611, new_n6612, new_n6613, new_n6614, new_n6615, new_n6616, new_n6617, new_n6618, new_n6619, new_n6620, new_n6621, new_n6622, new_n6623, new_n6624, new_n6625, new_n6626, new_n6627, new_n6628, new_n6629, new_n6630, new_n6631, new_n6632, new_n6633, new_n6634, new_n6635, new_n6636, new_n6637, new_n6638, new_n6639, new_n6640, new_n6641, new_n6642, new_n6643, new_n6644, new_n6645, new_n6646, new_n6647, new_n6648, new_n6649, new_n6650, new_n6651, new_n6652, new_n6653, new_n6654, new_n6655, new_n6656, new_n6657, new_n6658, new_n6659, new_n6660, new_n6661, new_n6662, new_n6663, new_n6664, new_n6665, new_n6666, new_n6667, new_n6668, new_n6669, new_n6670, new_n6671, new_n6672, new_n6673, new_n6674, new_n6675, new_n6676, new_n6677, new_n6678, new_n6679, new_n6680, new_n6681, new_n6682, new_n6683, new_n6684, new_n6685, new_n6686, new_n6687, new_n6688, new_n6689, new_n6690, new_n6691, new_n6692, new_n6693, new_n6694, new_n6695, new_n6696, new_n6697, new_n6698, new_n6699, new_n6700, new_n6701, new_n6702, new_n6703, new_n6704, new_n6705, new_n6706, new_n6707, new_n6708, new_n6709, new_n6710, new_n6711, new_n6712, new_n6713, new_n6714, new_n6715, new_n6716, new_n6717, new_n6718, new_n6719, new_n6720, new_n6721, new_n6722, new_n6723, new_n6724, new_n6725, new_n6726, new_n6727, new_n6728, new_n6729, new_n6730, new_n6731, new_n6732, new_n6733, new_n6734, new_n6735, new_n6736, new_n6737, new_n6738, new_n6739, new_n6740, new_n6741, new_n6742, new_n6743, new_n6744, new_n6745, new_n6746, new_n6747, new_n6748, new_n6749, new_n6750, new_n6751, new_n6752, new_n6753, new_n6754, new_n6755, new_n6756, new_n6757, new_n6758, new_n6759, new_n6760, new_n6761, new_n6762, new_n6763, new_n6764, new_n6765, new_n6766, new_n6767, new_n6768, new_n6769, new_n6770, new_n6771, new_n6772, new_n6773, new_n6774, new_n6775, new_n6776, new_n6777, new_n6778, new_n6779, new_n6780, new_n6781, new_n6782, new_n6783, new_n6784, new_n6785, new_n6786, new_n6787, new_n6788, new_n6789, new_n6790, new_n6791, new_n6792, new_n6793, new_n6794, new_n6795, new_n6796, new_n6797, new_n6798, new_n6799, new_n6800, new_n6801, new_n6802, new_n6803, new_n6804, new_n6805, new_n6806, new_n6807, new_n6808, new_n6809, new_n6810, new_n6811, new_n6812, new_n6813, new_n6814, new_n6815, new_n6816, new_n6817, new_n6818, new_n6819, new_n6820, new_n6821, new_n6822, new_n6823, new_n6824, new_n6825, new_n6826, new_n6827, new_n6828, new_n6829, new_n6830, new_n6831, new_n6832, new_n6833, new_n6834, new_n6835, new_n6836, new_n6837, new_n6838, new_n6839, new_n6840, new_n6841, new_n6842, new_n6843, new_n6844, new_n6845, new_n6846, new_n6847, new_n6848, new_n6849, new_n6850, new_n6851, new_n6852, new_n6853, new_n6854, new_n6855, new_n6856, new_n6857, new_n6858, new_n6859, new_n6860, new_n6861, new_n6862, new_n6863, new_n6864, new_n6865, new_n6866, new_n6867, new_n6868, new_n6869, new_n6870, new_n6871, new_n6872, new_n6873, new_n6874, new_n6875, new_n6876, new_n6877, new_n6878, new_n6879, new_n6880, new_n6881, new_n6882, new_n6883, new_n6884, new_n6885, new_n6886, new_n6887, new_n6888, new_n6889, new_n6890, new_n6891, new_n6892, new_n6893, new_n6894, new_n6895, new_n6896, new_n6897, new_n6898, new_n6899, new_n6900, new_n6901, new_n6902, new_n6903, new_n6904, new_n6905, new_n6906, new_n6907, new_n6908, new_n6909, new_n6910, new_n6911, new_n6912, new_n6913, new_n6914, new_n6915, new_n6916, new_n6917, new_n6918, new_n6919, new_n6920, new_n6921, new_n6922, new_n6923, new_n6924, new_n6925, new_n6926, new_n6927, new_n6928, new_n6929, new_n6930, new_n6931, new_n6932, new_n6933, new_n6934, new_n6935, new_n6936, new_n6937, new_n6938, new_n6939, new_n6940, new_n6941, new_n6942, new_n6943, new_n6944, new_n6945, new_n6946, new_n6947, new_n6948, new_n6949, new_n6950, new_n6951, new_n6952, new_n6953, new_n6954, new_n6955, new_n6956, new_n6957, new_n6958, new_n6959, new_n6960, new_n6961, new_n6962, new_n6963, new_n6964, new_n6965, new_n6966, new_n6967, new_n6968, new_n6969, new_n6970, new_n6971, new_n6972, new_n6973, new_n6974, new_n6975, new_n6976, new_n6977, new_n6978, new_n6979, new_n6980, new_n6981, new_n6982, new_n6983, new_n6984, new_n6985, new_n6986, new_n6987, new_n6988, new_n6989, new_n6990, new_n6991, new_n6992, new_n6993, new_n6994, new_n6995, new_n6996, new_n6997, new_n6998, new_n6999, new_n7000, new_n7001, new_n7002, new_n7003, new_n7004, new_n7005, new_n7006, new_n7007, new_n7008, new_n7009, new_n7010, new_n7011, new_n7012, new_n7013, new_n7014, new_n7015, new_n7016, new_n7017, new_n7018, new_n7019, new_n7020, new_n7021, new_n7022, new_n7023, new_n7024, new_n7025, new_n7026, new_n7027, new_n7028, new_n7029, new_n7030, new_n7031, new_n7032, new_n7033, new_n7034, new_n7035, new_n7036, new_n7037, new_n7038, new_n7039, new_n7040, new_n7041, new_n7042, new_n7043, new_n7044, new_n7045, new_n7046, new_n7047, new_n7048, new_n7049, new_n7050, new_n7051, new_n7052, new_n7053, new_n7054, new_n7055, new_n7056, new_n7057, new_n7058, new_n7059, new_n7060, new_n7061, new_n7062, new_n7063, new_n7064, new_n7065, new_n7066, new_n7067, new_n7068, new_n7069, new_n7070, new_n7071, new_n7072, new_n7073, new_n7074, new_n7075, new_n7076, new_n7077, new_n7078, new_n7079, new_n7080, new_n7081, new_n7082, new_n7083, new_n7084, new_n7085, new_n7086, new_n7087, new_n7088, new_n7089, new_n7090, new_n7091, new_n7092, new_n7093, new_n7094, new_n7095, new_n7096, new_n7097, new_n7098, new_n7099, new_n7100, new_n7101, new_n7102, new_n7103, new_n7104, new_n7105, new_n7106, new_n7107, new_n7108, new_n7109, new_n7110, new_n7111, new_n7112, new_n7113, new_n7114, new_n7115, new_n7116, new_n7117, new_n7118, new_n7119, new_n7120, new_n7121, new_n7122, new_n7123, new_n7124, new_n7125, new_n7126, new_n7127, new_n7128, new_n7129, new_n7130, new_n7131, new_n7132, new_n7133, new_n7134, new_n7135, new_n7136, new_n7137, new_n7138, new_n7139, new_n7140, new_n7141, new_n7142, new_n7143, new_n7144, new_n7145, new_n7146, new_n7147, new_n7148, new_n7149, new_n7150, new_n7151, new_n7152, new_n7153, new_n7154, new_n7155, new_n7156, new_n7157, new_n7158, new_n7159, new_n7160, new_n7161, new_n7162, new_n7163, new_n7164, new_n7165, new_n7166, new_n7167, new_n7168, new_n7169, new_n7170, new_n7171, new_n7172, new_n7173, new_n7174, new_n7175, new_n7176, new_n7177, new_n7178, new_n7179, new_n7180, new_n7181, new_n7182, new_n7183, new_n7184, new_n7185, new_n7186, new_n7187, new_n7188, new_n7189, new_n7190, new_n7191, new_n7192, new_n7193, new_n7194, new_n7195, new_n7196, new_n7197, new_n7198, new_n7199, new_n7200, new_n7201, new_n7202, new_n7203, new_n7204, new_n7205, new_n7206, new_n7207, new_n7208, new_n7209, new_n7210, new_n7211, new_n7212, new_n7213, new_n7214, new_n7215, new_n7216, new_n7217, new_n7218, new_n7219, new_n7220, new_n7221, new_n7222, new_n7223, new_n7224, new_n7225, new_n7226, new_n7227, new_n7228, new_n7229, new_n7230, new_n7231, new_n7232, new_n7233, new_n7234, new_n7235, new_n7236, new_n7237, new_n7238, new_n7239, new_n7240, new_n7241, new_n7242, new_n7243, new_n7244, new_n7245, new_n7246, new_n7247, new_n7248, new_n7249, new_n7250, new_n7251, new_n7252, new_n7253, new_n7254, new_n7255, new_n7256, new_n7257, new_n7258, new_n7259, new_n7260, new_n7261, new_n7262, new_n7263, new_n7264, new_n7265, new_n7266, new_n7267, new_n7268, new_n7269, new_n7270, new_n7271, new_n7272, new_n7273, new_n7274, new_n7275, new_n7276, new_n7277, new_n7278, new_n7279, new_n7280, new_n7281, new_n7282, new_n7283, new_n7284, new_n7285, new_n7286, new_n7287, new_n7288, new_n7289, new_n7290, new_n7291, new_n7292, new_n7293, new_n7294, new_n7295, new_n7296, new_n7297, new_n7298, new_n7299, new_n7300, new_n7301, new_n7302, new_n7303, new_n7304, new_n7305, new_n7306, new_n7307, new_n7308, new_n7309, new_n7310, new_n7311, new_n7312, new_n7313, new_n7314, new_n7315, new_n7316, new_n7317, new_n7318, new_n7319, new_n7320, new_n7321, new_n7322, new_n7323, new_n7324, new_n7325, new_n7326, new_n7327, new_n7328, new_n7329, new_n7330, new_n7331, new_n7332, new_n7333, new_n7334, new_n7335, new_n7336, new_n7337, new_n7338, new_n7339, new_n7340, new_n7341, new_n7342, new_n7343, new_n7344, new_n7345, new_n7346, new_n7347, new_n7348, new_n7349, new_n7350, new_n7351, new_n7352, new_n7353, new_n7354, new_n7355, new_n7356, new_n7357, new_n7358, new_n7359, new_n7360, new_n7361, new_n7362, new_n7363, new_n7364, new_n7365, new_n7366, new_n7367, new_n7368, new_n7369, new_n7370, new_n7371, new_n7372, new_n7373, new_n7374, new_n7375, new_n7376, new_n7377, new_n7378, new_n7379, new_n7380, new_n7381, new_n7382, new_n7383, new_n7384, new_n7385, new_n7386, new_n7387, new_n7388, new_n7389, new_n7390, new_n7391, new_n7392, new_n7393, new_n7394, new_n7395, new_n7396, new_n7397, new_n7398, new_n7399, new_n7400, new_n7401, new_n7402, new_n7403, new_n7404, new_n7405, new_n7406, new_n7407, new_n7408, new_n7409, new_n7410, new_n7411, new_n7412, new_n7413, new_n7414, new_n7415, new_n7416, new_n7417, new_n7418, new_n7419, new_n7420, new_n7421, new_n7422, new_n7423, new_n7424, new_n7425, new_n7426, new_n7427, new_n7428, new_n7429, new_n7430, new_n7431, new_n7432, new_n7433, new_n7434, new_n7435, new_n7436, new_n7437, new_n7438, new_n7439, new_n7440, new_n7441, new_n7442, new_n7443, new_n7444, new_n7445, new_n7446, new_n7447, new_n7448, new_n7449, new_n7450, new_n7451, new_n7452, new_n7453, new_n7454, new_n7455, new_n7456, new_n7457, new_n7458, new_n7459, new_n7460, new_n7461, new_n7462, new_n7463, new_n7464, new_n7465, new_n7466, new_n7467, new_n7468, new_n7469, new_n7470, new_n7471, new_n7472, new_n7473, new_n7474, new_n7475, new_n7476, new_n7477, new_n7478, new_n7479, new_n7480, new_n7481, new_n7482, new_n7483, new_n7484, new_n7485, new_n7486, new_n7487, new_n7488, new_n7489, new_n7490, new_n7491, new_n7492, new_n7493, new_n7494, new_n7495, new_n7496, new_n7497, new_n7498, new_n7499, new_n7500, new_n7501, new_n7502, new_n7503, new_n7504, new_n7505, new_n7506, new_n7507, new_n7508, new_n7509, new_n7510, new_n7511, new_n7512, new_n7513, new_n7514, new_n7515, new_n7516, new_n7517, new_n7518, new_n7519, new_n7520, new_n7521, new_n7522, new_n7523, new_n7524, new_n7525, new_n7526, new_n7527, new_n7528, new_n7529, new_n7530, new_n7531, new_n7532, new_n7533, new_n7534, new_n7535, new_n7536, new_n7537, new_n7538, new_n7539, new_n7540, new_n7541, new_n7542, new_n7543, new_n7544, new_n7545, new_n7546, new_n7547, new_n7548, new_n7549, new_n7550, new_n7551, new_n7552, new_n7553, new_n7554, new_n7555, new_n7556, new_n7557, new_n7558, new_n7559, new_n7560, new_n7561, new_n7562, new_n7563, new_n7564, new_n7565, new_n7566, new_n7567, new_n7568, new_n7569, new_n7570, new_n7571, new_n7572, new_n7573, new_n7574, new_n7575, new_n7576, new_n7577, new_n7578, new_n7579, new_n7580, new_n7581, new_n7582, new_n7583, new_n7584, new_n7585, new_n7586, new_n7587, new_n7588, new_n7589, new_n7590, new_n7591, new_n7592, new_n7593, new_n7594, new_n7595, new_n7596, new_n7597, new_n7598, new_n7599, new_n7600, new_n7601, new_n7602, new_n7603, new_n7604, new_n7605, new_n7606, new_n7607, new_n7608, new_n7609, new_n7610, new_n7611, new_n7612, new_n7613, new_n7614, new_n7615, new_n7616, new_n7617, new_n7618, new_n7619, new_n7620, new_n7621, new_n7622, new_n7623, new_n7624, new_n7625, new_n7626, new_n7627, new_n7628, new_n7629, new_n7630, new_n7631, new_n7632, new_n7633, new_n7634, new_n7635, new_n7636, new_n7637, new_n7638, new_n7639, new_n7640, new_n7641, new_n7642, new_n7643, new_n7644, new_n7645, new_n7646, new_n7647, new_n7648, new_n7649, new_n7650, new_n7651, new_n7652, new_n7653, new_n7654, new_n7655, new_n7656, new_n7657, new_n7658, new_n7659, new_n7660, new_n7661, new_n7662, new_n7663, new_n7664, new_n7665, new_n7666, new_n7667, new_n7668, new_n7669, new_n7670, new_n7671, new_n7672, new_n7673, new_n7674, new_n7675, new_n7676, new_n7677, new_n7678, new_n7679, new_n7680, new_n7681, new_n7682, new_n7683, new_n7684, new_n7685, new_n7686, new_n7687, new_n7688, new_n7689, new_n7690, new_n7691, new_n7692, new_n7693, new_n7694, new_n7695, new_n7696, new_n7697, new_n7698, new_n7699, new_n7700, new_n7701, new_n7702, new_n7703, new_n7704, new_n7705, new_n7706, new_n7707, new_n7708, new_n7709, new_n7710, new_n7711, new_n7712, new_n7713, new_n7714, new_n7715, new_n7716, new_n7717, new_n7718, new_n7719, new_n7720, new_n7721, new_n7722, new_n7723, new_n7724, new_n7725, new_n7726, new_n7727, new_n7728, new_n7729, new_n7730, new_n7731, new_n7732, new_n7733, new_n7734, new_n7735, new_n7736, new_n7737, new_n7738, new_n7739, new_n7740, new_n7741, new_n7742, new_n7743, new_n7744, new_n7745, new_n7746, new_n7747, new_n7748, new_n7749, new_n7750, new_n7751, new_n7752, new_n7753, new_n7754, new_n7755, new_n7756, new_n7757, new_n7758, new_n7759, new_n7760, new_n7761, new_n7762, new_n7763, new_n7764, new_n7765, new_n7766, new_n7767, new_n7768, new_n7769, new_n7770, new_n7771, new_n7772, new_n7773, new_n7774, new_n7775, new_n7776, new_n7777, new_n7778, new_n7779, new_n7780, new_n7781, new_n7782, new_n7783, new_n7784, new_n7785, new_n7786, new_n7787, new_n7788, new_n7789, new_n7790, new_n7791, new_n7792, new_n7793, new_n7794, new_n7795, new_n7796, new_n7797, new_n7798, new_n7799, new_n7800, new_n7801, new_n7802, new_n7803, new_n7804, new_n7805, new_n7806, new_n7807, new_n7808, new_n7809, new_n7810, new_n7811, new_n7812, new_n7813, new_n7814, new_n7815, new_n7816, new_n7817, new_n7818, new_n7819, new_n7820, new_n7821, new_n7822, new_n7823, new_n7824, new_n7825, new_n7826, new_n7827, new_n7828, new_n7829, new_n7830, new_n7831, new_n7832, new_n7833, new_n7834, new_n7835, new_n7836, new_n7837, new_n7838, new_n7839, new_n7840, new_n7841, new_n7842, new_n7843, new_n7844, new_n7845, new_n7846, new_n7847, new_n7848, new_n7849, new_n7850, new_n7851, new_n7852, new_n7853, new_n7854, new_n7855, new_n7856, new_n7857, new_n7858, new_n7859, new_n7860, new_n7861, new_n7862, new_n7863, new_n7864, new_n7865, new_n7866, new_n7867, new_n7868, new_n7869, new_n7870, new_n7871, new_n7872, new_n7873, new_n7874, new_n7875, new_n7876, new_n7877, new_n7878, new_n7879, new_n7880, new_n7881, new_n7882, new_n7883, new_n7884, new_n7885, new_n7886, new_n7887, new_n7888, new_n7889, new_n7890, new_n7891, new_n7892, new_n7893, new_n7894, new_n7895, new_n7896, new_n7897, new_n7898, new_n7899, new_n7900, new_n7901, new_n7902, new_n7903, new_n7904, new_n7905, new_n7906, new_n7907, new_n7908, new_n7909, new_n7910, new_n7911, new_n7912, new_n7913, new_n7914, new_n7915, new_n7916, new_n7917, new_n7918, new_n7919, new_n7920, new_n7921, new_n7922, new_n7923, new_n7924, new_n7925, new_n7926, new_n7927, new_n7928, new_n7929, new_n7930, new_n7931, new_n7932, new_n7933, new_n7934, new_n7935, new_n7936, new_n7937, new_n7938, new_n7939, new_n7940, new_n7941, new_n7942, new_n7943, new_n7944, new_n7945, new_n7946, new_n7947, new_n7948, new_n7949, new_n7950, new_n7951, new_n7952, new_n7953, new_n7954, new_n7955, new_n7956, new_n7957, new_n7958, new_n7959, new_n7960, new_n7961, new_n7962, new_n7963, new_n7964, new_n7965, new_n7966, new_n7967, new_n7968, new_n7969, new_n7970, new_n7971, new_n7972, new_n7973, new_n7974, new_n7975, new_n7976, new_n7977, new_n7978, new_n7979, new_n7980, new_n7981, new_n7982, new_n7983, new_n7984, new_n7985, new_n7986, new_n7987, new_n7988, new_n7989, new_n7990, new_n7991, new_n7992, new_n7993, new_n7994, new_n7995, new_n7996, new_n7997, new_n7998, new_n7999, new_n8000, new_n8001, new_n8002, new_n8003, new_n8004, new_n8005, new_n8006, new_n8007, new_n8008, new_n8009, new_n8010, new_n8011, new_n8012, new_n8013, new_n8014, new_n8015, new_n8016, new_n8017, new_n8018, new_n8019, new_n8020, new_n8021, new_n8022, new_n8023, new_n8024, new_n8025, new_n8026, new_n8027, new_n8028, new_n8029, new_n8030, new_n8031, new_n8032, new_n8033, new_n8034, new_n8035, new_n8036, new_n8037, new_n8038, new_n8039, new_n8040, new_n8041, new_n8042, new_n8043, new_n8044, new_n8045, new_n8046, new_n8047, new_n8048, new_n8049, new_n8050, new_n8051, new_n8052, new_n8053, new_n8054, new_n8055, new_n8056, new_n8057, new_n8058, new_n8059, new_n8060, new_n8061, new_n8062, new_n8063, new_n8064, new_n8065, new_n8066, new_n8067, new_n8068, new_n8069, new_n8070, new_n8071, new_n8072, new_n8073, new_n8074, new_n8075, new_n8076, new_n8077, new_n8078, new_n8079, new_n8080, new_n8081, new_n8082, new_n8083, new_n8084, new_n8085, new_n8086, new_n8087, new_n8088, new_n8089, new_n8090, new_n8091, new_n8092, new_n8093, new_n8094, new_n8095, new_n8096, new_n8097, new_n8098, new_n8099, new_n8100, new_n8101, new_n8102, new_n8103, new_n8104, new_n8105, new_n8106, new_n8107, new_n8108, new_n8109, new_n8110, new_n8111, new_n8112, new_n8113, new_n8114, new_n8115, new_n8116, new_n8117, new_n8118, new_n8119, new_n8120, new_n8121, new_n8122, new_n8123, new_n8124, new_n8125, new_n8126, new_n8127, new_n8128, new_n8129, new_n8130, new_n8131, new_n8132, new_n8133, new_n8134, new_n8135, new_n8136, new_n8137, new_n8138, new_n8139, new_n8140, new_n8141, new_n8142, new_n8143, new_n8144, new_n8145, new_n8146, new_n8147, new_n8148, new_n8149, new_n8150, new_n8151, new_n8152, new_n8153, new_n8154, new_n8155, new_n8156, new_n8157, new_n8158, new_n8159, new_n8160, new_n8161, new_n8162, new_n8163, new_n8164, new_n8165, new_n8166, new_n8167, new_n8168, new_n8169, new_n8170, new_n8171, new_n8172, new_n8173, new_n8174, new_n8175, new_n8176, new_n8177, new_n8178, new_n8179, new_n8180, new_n8181, new_n8182, new_n8183, new_n8184, new_n8185, new_n8186, new_n8187, new_n8188, new_n8189, new_n8190, new_n8191, new_n8192, new_n8193, new_n8194, new_n8195, new_n8196, new_n8197, new_n8198, new_n8199, new_n8200, new_n8201, new_n8202, new_n8203, new_n8204, new_n8205, new_n8206, new_n8207, new_n8208, new_n8209, new_n8210, new_n8211, new_n8212, new_n8213, new_n8214, new_n8215, new_n8216, new_n8217, new_n8218, new_n8219, new_n8220, new_n8221, new_n8222, new_n8223, new_n8224, new_n8225, new_n8226, new_n8227, new_n8228, new_n8229, new_n8230, new_n8231, new_n8232, new_n8233, new_n8234, new_n8235, new_n8236, new_n8237, new_n8238, new_n8239, new_n8240, new_n8241, new_n8242, new_n8243, new_n8244, new_n8245, new_n8246, new_n8247, new_n8248, new_n8249, new_n8250, new_n8251, new_n8252, new_n8253, new_n8254, new_n8255, new_n8256, new_n8257, new_n8258, new_n8259, new_n8260, new_n8261, new_n8262, new_n8263, new_n8264, new_n8265, new_n8266, new_n8267, new_n8268, new_n8269, new_n8270, new_n8271, new_n8272, new_n8273, new_n8274, new_n8275, new_n8276, new_n8277, new_n8278, new_n8279, new_n8280, new_n8281, new_n8282, new_n8283, new_n8284, new_n8285, new_n8286, new_n8287, new_n8288, new_n8289, new_n8290, new_n8291, new_n8292, new_n8293, new_n8294, new_n8295, new_n8296, new_n8297, new_n8298, new_n8299, new_n8300, new_n8301, new_n8302, new_n8303, new_n8304, new_n8305, new_n8306, new_n8307, new_n8308, new_n8309, new_n8310, new_n8311, new_n8312, new_n8313, new_n8314, new_n8315, new_n8316, new_n8317, new_n8318, new_n8319, new_n8320, new_n8321, new_n8322, new_n8323, new_n8324, new_n8325, new_n8326, new_n8327, new_n8328, new_n8329, new_n8330, new_n8331, new_n8332, new_n8333, new_n8334, new_n8335, new_n8336, new_n8337, new_n8338, new_n8339, new_n8340, new_n8341, new_n8342, new_n8343, new_n8344, new_n8345, new_n8346, new_n8347, new_n8348, new_n8349, new_n8350, new_n8351, new_n8352, new_n8353, new_n8354, new_n8355, new_n8356, new_n8357, new_n8358, new_n8359, new_n8360, new_n8361, new_n8362, new_n8363, new_n8364, new_n8365, new_n8366, new_n8367, new_n8368, new_n8369, new_n8370, new_n8371, new_n8372, new_n8373, new_n8374, new_n8375, new_n8376, new_n8377, new_n8378, new_n8379, new_n8380, new_n8381, new_n8382, new_n8383, new_n8384, new_n8385, new_n8386, new_n8387, new_n8388, new_n8389, new_n8390, new_n8391, new_n8392, new_n8393, new_n8394, new_n8395, new_n8396, new_n8397, new_n8398, new_n8399, new_n8400, new_n8401, new_n8402, new_n8403, new_n8404, new_n8405, new_n8406, new_n8407, new_n8408, new_n8409, new_n8410, new_n8411, new_n8412, new_n8413, new_n8414, new_n8415, new_n8416, new_n8417, new_n8418, new_n8419, new_n8420, new_n8421, new_n8422, new_n8423, new_n8424, new_n8425, new_n8426, new_n8427, new_n8428, new_n8429, new_n8430, new_n8431, new_n8432, new_n8433, new_n8434, new_n8435, new_n8436, new_n8437, new_n8438, new_n8439, new_n8440, new_n8441, new_n8442, new_n8443, new_n8444, new_n8445, new_n8446, new_n8447, new_n8448, new_n8449, new_n8450, new_n8451, new_n8452, new_n8453, new_n8454, new_n8455, new_n8456, new_n8457, new_n8458, new_n8459, new_n8460, new_n8461, new_n8462, new_n8463, new_n8464, new_n8465, new_n8466, new_n8467, new_n8468, new_n8469, new_n8470, new_n8471, new_n8472, new_n8473, new_n8474, new_n8475, new_n8476, new_n8477, new_n8478, new_n8479, new_n8480, new_n8481, new_n8482, new_n8483, new_n8484, new_n8485, new_n8486, new_n8487, new_n8488, new_n8489, new_n8490, new_n8491, new_n8492, new_n8493, new_n8494, new_n8495, new_n8496, new_n8497, new_n8498, new_n8499, new_n8500, new_n8501, new_n8502, new_n8503, new_n8504, new_n8505, new_n8506, new_n8507, new_n8508, new_n8509, new_n8510, new_n8511, new_n8512, new_n8513, new_n8514, new_n8515, new_n8516, new_n8517, new_n8518, new_n8519, new_n8520, new_n8521, new_n8522, new_n8523, new_n8524, new_n8525, new_n8526, new_n8527, new_n8528, new_n8529, new_n8530, new_n8531, new_n8532, new_n8533, new_n8534, new_n8535, new_n8536, new_n8537, new_n8538, new_n8539, new_n8540, new_n8541, new_n8542, new_n8543, new_n8544, new_n8545, new_n8546, new_n8547, new_n8548, new_n8549, new_n8550, new_n8551, new_n8552, new_n8553, new_n8554, new_n8555, new_n8556, new_n8557, new_n8558, new_n8559, new_n8560, new_n8561, new_n8562, new_n8563, new_n8564, new_n8565, new_n8566, new_n8567, new_n8568, new_n8569, new_n8570, new_n8571, new_n8572, new_n8573, new_n8574, new_n8575, new_n8576, new_n8577, new_n8578, new_n8579, new_n8580, new_n8581, new_n8582, new_n8583, new_n8584, new_n8585, new_n8586, new_n8587, new_n8588, new_n8589, new_n8590, new_n8591, new_n8592, new_n8593, new_n8594, new_n8595, new_n8596, new_n8597, new_n8598, new_n8599, new_n8600, new_n8601, new_n8602, new_n8603, new_n8604, new_n8605, new_n8606, new_n8607, new_n8608, new_n8609, new_n8610, new_n8611, new_n8612, new_n8613, new_n8614, new_n8615, new_n8616, new_n8617, new_n8618, new_n8619, new_n8620, new_n8621, new_n8622, new_n8623, new_n8624, new_n8625, new_n8626, new_n8627, new_n8628, new_n8629, new_n8630, new_n8631, new_n8632, new_n8633, new_n8634, new_n8635, new_n8636, new_n8637, new_n8638, new_n8639, new_n8640, new_n8641, new_n8642, new_n8643, new_n8644, new_n8645, new_n8646, new_n8647, new_n8648, new_n8649, new_n8650, new_n8651, new_n8652, new_n8653, new_n8654, new_n8655, new_n8656, new_n8657, new_n8658, new_n8659, new_n8660, new_n8661, new_n8662, new_n8663, new_n8664, new_n8665, new_n8666, new_n8667, new_n8668, new_n8669, new_n8670, new_n8671, new_n8672, new_n8673, new_n8674, new_n8675, new_n8676, new_n8677, new_n8678, new_n8679, new_n8680, new_n8681, new_n8682, new_n8683, new_n8684, new_n8685, new_n8686, new_n8687, new_n8688, new_n8689, new_n8690, new_n8691, new_n8692, new_n8693, new_n8694, new_n8695, new_n8696, new_n8697, new_n8698, new_n8699, new_n8700, new_n8701, new_n8702, new_n8703, new_n8704, new_n8705, new_n8706, new_n8707, new_n8708, new_n8709, new_n8710, new_n8711, new_n8712, new_n8713, new_n8714, new_n8715, new_n8716, new_n8717, new_n8718, new_n8719, new_n8720, new_n8721, new_n8722, new_n8723, new_n8724, new_n8725, new_n8726, new_n8727, new_n8728, new_n8729, new_n8730, new_n8731, new_n8732, new_n8733, new_n8734, new_n8735, new_n8736, new_n8737, new_n8738, new_n8739, new_n8740, new_n8741, new_n8742, new_n8743, new_n8744, new_n8745, new_n8746, new_n8747, new_n8748, new_n8749, new_n8750, new_n8751, new_n8752, new_n8753, new_n8754, new_n8755, new_n8756, new_n8757, new_n8758, new_n8759, new_n8760, new_n8761, new_n8762, new_n8763, new_n8764, new_n8765, new_n8766, new_n8767, new_n8768, new_n8769, new_n8770, new_n8771, new_n8772, new_n8773, new_n8774, new_n8775, new_n8776, new_n8777, new_n8778, new_n8779, new_n8780, new_n8781, new_n8782, new_n8783, new_n8784, new_n8785, new_n8786, new_n8787, new_n8788, new_n8789, new_n8790, new_n8791, new_n8792, new_n8793, new_n8794, new_n8795, new_n8796, new_n8797, new_n8798, new_n8799, new_n8800, new_n8801, new_n8802, new_n8803, new_n8804, new_n8805, new_n8806, new_n8807, new_n8808, new_n8809, new_n8810, new_n8811, new_n8812, new_n8813, new_n8814, new_n8815, new_n8816, new_n8817, new_n8818, new_n8819, new_n8820, new_n8821, new_n8822, new_n8823, new_n8824, new_n8825, new_n8826, new_n8827, new_n8828, new_n8829, new_n8830, new_n8831, new_n8832, new_n8833, new_n8834, new_n8835, new_n8836, new_n8837, new_n8838, new_n8839, new_n8840, new_n8841, new_n8842, new_n8843, new_n8844, new_n8845, new_n8846, new_n8847, new_n8848, new_n8849, new_n8850, new_n8851, new_n8852, new_n8853, new_n8854, new_n8855, new_n8856, new_n8857, new_n8858, new_n8859, new_n8860, new_n8861, new_n8862, new_n8863, new_n8864, new_n8865, new_n8866, new_n8867, new_n8868, new_n8869, new_n8870, new_n8871, new_n8872, new_n8873, new_n8874, new_n8875, new_n8876, new_n8877, new_n8878, new_n8879, new_n8880, new_n8881, new_n8882, new_n8883, new_n8884, new_n8885, new_n8886, new_n8887, new_n8888, new_n8889, new_n8890, new_n8891, new_n8892, new_n8893, new_n8894, new_n8895, new_n8896, new_n8897, new_n8898, new_n8899, new_n8900, new_n8901, new_n8902, new_n8903, new_n8904, new_n8905, new_n8906, new_n8907, new_n8908, new_n8909, new_n8910, new_n8911, new_n8912, new_n8913, new_n8914, new_n8915, new_n8916, new_n8917, new_n8918, new_n8919, new_n8920, new_n8921, new_n8922, new_n8923, new_n8924, new_n8925, new_n8926, new_n8927, new_n8928, new_n8929, new_n8930, new_n8931, new_n8932, new_n8933, new_n8934, new_n8935, new_n8936, new_n8937, new_n8938, new_n8939, new_n8940, new_n8941, new_n8942, new_n8943, new_n8944, new_n8945, new_n8946, new_n8947, new_n8948, new_n8949, new_n8950, new_n8951, new_n8952, new_n8953, new_n8954, new_n8955, new_n8956, new_n8957, new_n8958, new_n8959, new_n8960, new_n8961, new_n8962, new_n8963, new_n8964, new_n8965, new_n8966, new_n8967, new_n8968, new_n8969, new_n8970, new_n8971, new_n8972, new_n8973, new_n8974, new_n8975, new_n8976, new_n8977, new_n8978, new_n8979, new_n8980, new_n8981, new_n8982, new_n8983, new_n8984, new_n8985, new_n8986, new_n8987, new_n8988, new_n8989, new_n8990, new_n8991, new_n8992, new_n8993, new_n8994, new_n8995, new_n8996, new_n8997, new_n8998, new_n8999, new_n9000, new_n9001, new_n9002, new_n9003, new_n9004, new_n9005, new_n9006, new_n9007, new_n9008, new_n9009, new_n9010, new_n9011, new_n9012, new_n9013, new_n9014, new_n9015, new_n9016, new_n9017, new_n9018, new_n9019, new_n9020, new_n9021, new_n9022, new_n9023, new_n9024, new_n9025, new_n9026, new_n9027, new_n9028, new_n9029, new_n9030, new_n9031, new_n9032, new_n9033, new_n9034, new_n9035, new_n9036, new_n9037, new_n9038, new_n9039, new_n9040, new_n9041, new_n9042, new_n9043, new_n9044, new_n9045, new_n9046, new_n9047, new_n9048, new_n9049, new_n9050, new_n9051, new_n9052, new_n9053, new_n9054, new_n9055, new_n9056, new_n9057, new_n9058, new_n9059, new_n9060, new_n9061, new_n9062, new_n9063, new_n9064, new_n9065, new_n9066, new_n9067, new_n9068, new_n9069, new_n9070, new_n9071, new_n9072, new_n9073, new_n9074, new_n9075, new_n9076, new_n9077, new_n9078, new_n9079, new_n9080, new_n9081, new_n9082, new_n9083, new_n9084, new_n9085, new_n9086, new_n9087, new_n9088, new_n9089, new_n9090, new_n9091, new_n9092, new_n9093, new_n9094, new_n9095, new_n9096, new_n9097, new_n9098, new_n9099, new_n9100, new_n9101, new_n9102, new_n9103, new_n9104, new_n9105, new_n9106, new_n9107, new_n9108, new_n9109, new_n9110, new_n9111, new_n9112, new_n9113, new_n9114, new_n9115, new_n9116, new_n9117, new_n9118, new_n9119, new_n9120, new_n9121, new_n9122, new_n9123, new_n9124, new_n9125, new_n9126, new_n9127, new_n9128, new_n9129, new_n9130, new_n9131, new_n9132, new_n9133, new_n9134, new_n9135, new_n9136, new_n9137, new_n9138, new_n9139, new_n9140, new_n9141, new_n9142, new_n9143, new_n9144, new_n9145, new_n9146, new_n9147, new_n9148, new_n9149, new_n9150, new_n9151, new_n9152, new_n9153, new_n9154, new_n9155, new_n9156, new_n9157, new_n9158, new_n9159, new_n9160, new_n9161, new_n9162, new_n9163, new_n9164, new_n9165, new_n9166, new_n9167, new_n9168, new_n9169, new_n9170, new_n9171, new_n9172, new_n9173, new_n9174, new_n9175, new_n9176, new_n9177, new_n9178, new_n9179, new_n9180, new_n9181, new_n9182, new_n9183, new_n9184, new_n9185, new_n9186, new_n9187, new_n9188, new_n9189, new_n9190, new_n9191, new_n9192, new_n9193, new_n9194, new_n9195, new_n9196, new_n9197, new_n9198, new_n9199, new_n9200, new_n9201, new_n9202, new_n9203, new_n9204, new_n9205, new_n9206, new_n9207, new_n9208, new_n9209, new_n9210, new_n9211, new_n9212, new_n9213, new_n9214, new_n9215, new_n9216, new_n9217, new_n9218, new_n9219, new_n9220, new_n9221, new_n9222, new_n9223, new_n9224, new_n9225, new_n9226, new_n9227, new_n9228, new_n9229, new_n9230, new_n9231, new_n9232, new_n9233, new_n9234, new_n9235, new_n9236, new_n9237, new_n9238, new_n9239, new_n9240, new_n9241, new_n9242, new_n9243, new_n9244, new_n9245, new_n9246, new_n9247, new_n9248, new_n9249, new_n9250, new_n9251, new_n9252, new_n9253, new_n9254, new_n9255, new_n9256, new_n9257, new_n9258, new_n9259, new_n9260, new_n9261, new_n9262, new_n9263, new_n9264, new_n9265, new_n9266, new_n9267, new_n9268, new_n9269, new_n9270, new_n9271, new_n9272, new_n9273, new_n9274, new_n9275, new_n9276, new_n9277, new_n9278, new_n9279, new_n9280, new_n9281, new_n9282, new_n9283, new_n9284, new_n9285, new_n9286, new_n9287, new_n9288, new_n9289, new_n9290, new_n9291, new_n9292, new_n9293, new_n9294, new_n9295, new_n9296, new_n9297, new_n9298, new_n9299, new_n9300, new_n9301, new_n9302, new_n9303, new_n9304, new_n9305, new_n9306, new_n9307, new_n9308, new_n9309, new_n9310, new_n9311, new_n9312, new_n9313, new_n9314, new_n9315, new_n9316, new_n9317, new_n9318, new_n9319, new_n9320, new_n9321, new_n9322, new_n9323, new_n9324, new_n9325, new_n9326, new_n9327, new_n9328, new_n9329, new_n9330, new_n9331, new_n9332, new_n9333, new_n9334, new_n9335, new_n9336, new_n9337, new_n9338, new_n9339, new_n9340, new_n9341, new_n9342, new_n9343, new_n9344, new_n9345, new_n9346, new_n9347, new_n9348, new_n9349, new_n9350, new_n9351, new_n9352, new_n9353, new_n9354, new_n9355, new_n9356, new_n9357, new_n9358, new_n9359, new_n9360, new_n9361, new_n9362, new_n9363, new_n9364, new_n9365, new_n9366, new_n9367, new_n9368, new_n9369, new_n9370, new_n9371, new_n9372, new_n9373, new_n9374, new_n9375, new_n9376, new_n9377, new_n9378, new_n9379, new_n9380, new_n9381, new_n9382, new_n9383, new_n9384, new_n9385, new_n9386, new_n9387, new_n9388, new_n9389, new_n9390, new_n9391, new_n9392, new_n9393, new_n9394, new_n9395, new_n9396, new_n9397, new_n9398, new_n9399, new_n9400, new_n9401, new_n9402, new_n9403, new_n9404, new_n9405, new_n9406, new_n9407, new_n9408, new_n9409, new_n9410, new_n9411, new_n9412, new_n9413, new_n9414, new_n9415, new_n9416, new_n9417, new_n9418, new_n9419, new_n9420, new_n9421, new_n9422, new_n9423, new_n9424, new_n9425, new_n9426, new_n9427, new_n9428, new_n9429, new_n9430, new_n9431, new_n9432, new_n9433, new_n9434, new_n9435, new_n9436, new_n9437, new_n9438, new_n9439, new_n9440, new_n9441, new_n9442, new_n9443, new_n9444, new_n9445, new_n9446, new_n9447, new_n9448, new_n9449, new_n9450, new_n9451, new_n9452, new_n9453, new_n9454, new_n9455, new_n9456, new_n9457, new_n9458, new_n9459, new_n9460, new_n9461, new_n9462, new_n9463, new_n9464, new_n9465, new_n9466, new_n9467, new_n9468, new_n9469, new_n9470, new_n9471, new_n9472, new_n9473, new_n9474, new_n9475, new_n9476, new_n9477, new_n9478, new_n9479, new_n9480, new_n9481, new_n9482, new_n9483, new_n9484, new_n9485, new_n9486, new_n9487, new_n9488, new_n9489, new_n9490, new_n9491, new_n9492, new_n9493, new_n9494, new_n9495, new_n9496, new_n9497, new_n9498, new_n9499, new_n9500, new_n9501, new_n9502, new_n9503, new_n9504, new_n9505, new_n9506, new_n9507, new_n9508, new_n9509, new_n9510, new_n9511, new_n9512, new_n9513, new_n9514, new_n9515, new_n9516, new_n9517, new_n9518, new_n9519, new_n9520, new_n9521, new_n9522, new_n9523, new_n9524, new_n9525, new_n9526, new_n9527, new_n9528, new_n9529, new_n9530, new_n9531, new_n9532, new_n9533, new_n9534, new_n9535, new_n9536, new_n9537, new_n9538, new_n9539, new_n9540, new_n9541, new_n9542, new_n9543, new_n9544, new_n9545, new_n9546, new_n9547, new_n9548, new_n9549, new_n9550, new_n9551, new_n9552, new_n9553, new_n9554, new_n9555, new_n9556, new_n9557, new_n9558, new_n9559, new_n9560, new_n9561, new_n9562, new_n9563, new_n9564, new_n9565, new_n9566, new_n9567, new_n9568, new_n9569, new_n9570, new_n9571, new_n9572, new_n9573, new_n9574, new_n9575, new_n9576, new_n9577, new_n9578, new_n9579, new_n9580, new_n9581, new_n9582, new_n9583, new_n9584, new_n9585, new_n9586, new_n9587, new_n9588, new_n9589, new_n9590, new_n9591, new_n9592, new_n9593, new_n9594, new_n9595, new_n9596, new_n9597, new_n9598, new_n9599, new_n9600, new_n9601, new_n9602, new_n9603, new_n9604, new_n9605, new_n9606, new_n9607, new_n9608, new_n9609, new_n9610, new_n9611, new_n9612, new_n9613, new_n9614, new_n9615, new_n9616, new_n9617, new_n9618, new_n9619, new_n9620, new_n9621, new_n9622, new_n9623, new_n9624, new_n9625, new_n9626, new_n9627, new_n9628, new_n9629, new_n9630, new_n9631, new_n9632, new_n9633, new_n9634, new_n9635, new_n9636, new_n9637, new_n9638, new_n9639, new_n9640, new_n9641, new_n9642, new_n9643, new_n9644, new_n9645, new_n9646, new_n9647, new_n9648, new_n9649, new_n9650, new_n9651, new_n9652, new_n9653, new_n9654, new_n9655, new_n9656, new_n9657, new_n9658, new_n9659, new_n9660, new_n9661, new_n9662, new_n9663, new_n9664, new_n9665, new_n9666, new_n9667, new_n9668, new_n9669, new_n9670, new_n9671, new_n9672, new_n9673, new_n9674, new_n9675, new_n9676, new_n9677, new_n9678, new_n9679, new_n9680, new_n9681, new_n9682, new_n9683, new_n9684, new_n9685, new_n9686, new_n9687, new_n9688, new_n9689, new_n9690, new_n9691, new_n9692, new_n9693, new_n9694, new_n9695, new_n9696, new_n9697, new_n9698, new_n9699, new_n9700, new_n9701, new_n9702, new_n9703, new_n9704, new_n9705, new_n9706, new_n9707, new_n9708, new_n9709, new_n9710, new_n9711, new_n9712, new_n9713, new_n9714, new_n9715, new_n9716, new_n9717, new_n9718, new_n9719, new_n9720, new_n9721, new_n9722, new_n9723, new_n9724, new_n9725, new_n9726, new_n9727, new_n9728, new_n9729, new_n9730, new_n9731, new_n9732, new_n9733, new_n9734, new_n9735, new_n9736, new_n9737, new_n9738, new_n9739, new_n9740, new_n9741, new_n9742, new_n9743, new_n9744, new_n9745, new_n9746, new_n9747, new_n9748, new_n9749, new_n9750, new_n9751, new_n9752, new_n9753, new_n9754, new_n9755, new_n9756, new_n9757, new_n9758, new_n9759, new_n9760, new_n9761, new_n9762, new_n9763, new_n9764, new_n9765, new_n9766, new_n9767, new_n9768, new_n9769, new_n9770, new_n9771, new_n9772, new_n9773, new_n9774, new_n9775, new_n9776, new_n9777, new_n9778, new_n9779, new_n9780, new_n9781, new_n9782, new_n9783, new_n9784, new_n9785, new_n9786, new_n9787, new_n9788, new_n9789, new_n9790, new_n9791, new_n9792, new_n9793, new_n9794, new_n9795, new_n9796, new_n9797, new_n9798, new_n9799, new_n9800, new_n9801, new_n9802, new_n9803, new_n9804, new_n9805, new_n9806, new_n9807, new_n9808, new_n9809, new_n9810, new_n9811, new_n9812, new_n9813, new_n9814, new_n9815, new_n9816, new_n9817, new_n9818, new_n9819, new_n9820, new_n9821, new_n9822, new_n9823, new_n9824, new_n9825, new_n9826, new_n9827, new_n9828, new_n9829, new_n9830, new_n9831, new_n9832, new_n9833, new_n9834, new_n9835, new_n9836, new_n9837, new_n9838, new_n9839, new_n9840, new_n9841, new_n9842, new_n9843, new_n9844, new_n9845, new_n9846, new_n9847, new_n9848, new_n9849, new_n9850, new_n9851, new_n9852, new_n9853, new_n9854, new_n9855, new_n9856, new_n9857, new_n9858, new_n9859, new_n9860, new_n9861, new_n9862, new_n9863, new_n9864, new_n9865, new_n9866, new_n9867, new_n9868, new_n9869, new_n9870, new_n9871, new_n9872, new_n9873, new_n9874, new_n9875, new_n9876, new_n9877, new_n9878, new_n9879, new_n9880, new_n9881, new_n9882, new_n9883, new_n9884, new_n9885, new_n9886, new_n9887, new_n9888, new_n9889, new_n9890, new_n9891, new_n9892, new_n9893, new_n9894, new_n9895, new_n9896, new_n9897, new_n9898, new_n9899, new_n9900, new_n9901, new_n9902, new_n9903, new_n9904, new_n9905, new_n9906, new_n9907, new_n9908, new_n9909, new_n9910, new_n9911, new_n9912, new_n9913, new_n9914, new_n9915, new_n9916, new_n9917, new_n9918, new_n9919, new_n9920, new_n9921, new_n9922, new_n9923, new_n9924, new_n9925, new_n9926, new_n9927, new_n9928, new_n9929, new_n9930, new_n9931, new_n9932, new_n9933, new_n9934, new_n9935, new_n9936, new_n9937, new_n9938, new_n9939, new_n9940, new_n9941, new_n9942, new_n9943, new_n9944, new_n9945, new_n9946, new_n9947, new_n9948, new_n9949, new_n9950, new_n9951, new_n9952, new_n9953, new_n9954, new_n9955, new_n9956, new_n9957, new_n9958, new_n9959, new_n9960, new_n9961, new_n9962, new_n9963, new_n9964, new_n9965, new_n9966, new_n9967, new_n9968, new_n9969, new_n9970, new_n9971, new_n9972, new_n9973, new_n9974, new_n9975, new_n9976, new_n9977, new_n9978, new_n9979, new_n9980, new_n9981, new_n9982, new_n9983, new_n9984, new_n9985, new_n9986, new_n9987, new_n9988, new_n9989, new_n9990, new_n9991, new_n9992, new_n9993, new_n9994, new_n9995, new_n9996, new_n9997, new_n9998, new_n9999, new_n10000, new_n10001, new_n10002, new_n10003, new_n10004, new_n10005, new_n10006, new_n10007, new_n10008, new_n10009, new_n10010, new_n10011, new_n10012, new_n10013, new_n10014, new_n10015, new_n10016, new_n10017, new_n10018, new_n10019, new_n10020, new_n10021, new_n10022, new_n10023, new_n10024, new_n10025, new_n10026, new_n10027, new_n10028, new_n10029, new_n10030, new_n10031, new_n10032, new_n10033, new_n10034, new_n10035, new_n10036, new_n10037, new_n10038, new_n10039, new_n10040, new_n10041, new_n10042, new_n10043, new_n10044, new_n10045, new_n10046, new_n10047, new_n10048, new_n10049, new_n10050, new_n10051, new_n10052, new_n10053, new_n10054, new_n10055, new_n10056, new_n10057, new_n10058, new_n10059, new_n10060, new_n10061, new_n10062, new_n10063, new_n10064, new_n10065, new_n10066, new_n10067, new_n10068, new_n10069, new_n10070, new_n10071, new_n10072, new_n10073, new_n10074, new_n10075, new_n10076, new_n10077, new_n10078, new_n10079, new_n10080, new_n10081, new_n10082, new_n10083, new_n10084, new_n10085, new_n10086, new_n10087, new_n10088, new_n10089, new_n10090, new_n10091, new_n10092, new_n10093, new_n10094, new_n10095, new_n10096, new_n10097, new_n10098, new_n10099, new_n10100, new_n10101, new_n10102, new_n10103, new_n10104, new_n10105, new_n10106, new_n10107, new_n10108, new_n10109, new_n10110, new_n10111, new_n10112, new_n10113, new_n10114, new_n10115, new_n10116, new_n10117, new_n10118, new_n10119, new_n10120, new_n10121, new_n10122, new_n10123, new_n10124, new_n10125, new_n10126, new_n10127, new_n10128, new_n10129, new_n10130, new_n10131, new_n10132, new_n10133, new_n10134, new_n10135, new_n10136, new_n10137, new_n10138, new_n10139, new_n10140, new_n10141, new_n10142, new_n10143, new_n10144, new_n10145, new_n10146, new_n10147, new_n10148, new_n10149, new_n10150, new_n10151, new_n10152, new_n10153, new_n10154, new_n10155, new_n10156, new_n10157, new_n10158, new_n10159, new_n10160, new_n10161, new_n10162, new_n10163, new_n10164, new_n10165, new_n10166, new_n10167, new_n10168, new_n10169, new_n10170, new_n10171, new_n10172, new_n10173, new_n10174, new_n10175, new_n10176, new_n10177, new_n10178, new_n10179, new_n10180, new_n10181, new_n10182, new_n10183, new_n10184, new_n10185, new_n10186, new_n10187, new_n10188, new_n10189, new_n10190, new_n10191, new_n10192, new_n10193, new_n10194, new_n10195, new_n10196, new_n10197, new_n10198, new_n10199, new_n10200, new_n10201, new_n10202, new_n10203, new_n10204, new_n10205, new_n10206, new_n10207, new_n10208, new_n10209, new_n10210, new_n10211, new_n10212, new_n10213, new_n10214, new_n10215, new_n10216, new_n10217, new_n10218, new_n10219, new_n10220, new_n10221, new_n10222, new_n10223, new_n10224, new_n10225, new_n10226, new_n10227, new_n10228, new_n10229, new_n10230, new_n10231, new_n10232, new_n10233, new_n10234, new_n10235, new_n10236, new_n10237, new_n10238, new_n10239, new_n10240, new_n10241, new_n10242, new_n10243, new_n10244, new_n10245, new_n10246, new_n10247, new_n10248, new_n10249, new_n10250, new_n10251, new_n10252, new_n10253, new_n10254, new_n10255, new_n10256, new_n10257, new_n10258, new_n10259, new_n10260, new_n10261, new_n10262, new_n10263, new_n10264, new_n10265, new_n10266, new_n10267, new_n10268, new_n10269, new_n10270, new_n10271, new_n10272, new_n10273, new_n10274, new_n10275, new_n10276, new_n10277, new_n10278, new_n10279, new_n10280, new_n10281, new_n10282, new_n10283, new_n10284, new_n10285, new_n10286, new_n10287, new_n10288, new_n10289, new_n10290, new_n10291, new_n10292, new_n10293, new_n10294, new_n10295, new_n10296, new_n10297, new_n10298, new_n10299, new_n10300, new_n10301, new_n10302, new_n10303, new_n10304, new_n10305, new_n10306, new_n10307, new_n10308, new_n10309, new_n10310, new_n10311, new_n10312, new_n10313, new_n10314, new_n10315, new_n10316, new_n10317, new_n10318, new_n10319, new_n10320, new_n10321, new_n10322, new_n10323, new_n10324, new_n10325, new_n10326, new_n10327, new_n10328, new_n10329, new_n10330, new_n10331, new_n10332, new_n10333, new_n10334, new_n10335, new_n10336, new_n10337, new_n10338, new_n10339, new_n10340, new_n10341, new_n10342, new_n10343, new_n10344, new_n10345, new_n10346, new_n10347, new_n10348, new_n10349, new_n10350, new_n10351, new_n10352, new_n10353, new_n10354, new_n10355, new_n10356, new_n10357, new_n10358, new_n10359, new_n10360, new_n10361, new_n10362, new_n10363, new_n10364, new_n10365, new_n10366, new_n10367, new_n10368, new_n10369, new_n10370, new_n10371, new_n10372, new_n10373, new_n10374, new_n10375, new_n10376, new_n10377, new_n10378, new_n10379, new_n10380, new_n10381, new_n10382, new_n10383, new_n10384, new_n10385, new_n10386, new_n10387, new_n10388, new_n10389, new_n10390, new_n10391, new_n10392, new_n10393, new_n10394, new_n10395, new_n10396, new_n10397, new_n10398, new_n10399, new_n10400, new_n10401, new_n10402, new_n10403, new_n10404, new_n10405, new_n10406, new_n10407, new_n10408, new_n10409, new_n10410, new_n10411, new_n10412, new_n10413, new_n10414, new_n10415, new_n10416, new_n10417, new_n10418, new_n10419, new_n10420, new_n10421, new_n10422, new_n10423, new_n10424, new_n10425, new_n10426, new_n10427, new_n10428, new_n10429, new_n10430, new_n10431, new_n10432, new_n10433, new_n10434, new_n10435, new_n10436, new_n10437, new_n10438, new_n10439, new_n10440, new_n10441, new_n10442, new_n10443, new_n10444, new_n10445, new_n10446, new_n10447, new_n10448, new_n10449, new_n10450, new_n10451, new_n10452, new_n10453, new_n10454, new_n10455, new_n10456, new_n10457, new_n10458, new_n10459, new_n10460, new_n10461, new_n10462, new_n10463, new_n10464, new_n10465, new_n10466, new_n10467, new_n10468, new_n10469, new_n10470, new_n10471, new_n10472, new_n10473, new_n10474, new_n10475, new_n10476, new_n10477, new_n10478, new_n10479, new_n10480, new_n10481, new_n10482, new_n10483, new_n10484, new_n10485, new_n10486, new_n10487, new_n10488, new_n10489, new_n10490, new_n10491, new_n10492, new_n10493, new_n10494, new_n10495, new_n10496, new_n10497, new_n10498, new_n10499, new_n10500, new_n10501, new_n10502, new_n10503, new_n10504, new_n10505, new_n10506, new_n10507, new_n10508, new_n10509, new_n10510, new_n10511, new_n10512, new_n10513, new_n10514, new_n10515, new_n10516, new_n10517, new_n10518, new_n10519, new_n10520, new_n10521, new_n10522, new_n10523, new_n10524, new_n10525, new_n10526, new_n10527, new_n10528, new_n10529, new_n10530, new_n10531, new_n10532, new_n10533, new_n10534, new_n10535, new_n10536, new_n10537, new_n10538, new_n10539, new_n10540, new_n10541, new_n10542, new_n10543, new_n10544, new_n10545, new_n10546, new_n10547, new_n10548, new_n10549, new_n10550, new_n10551, new_n10552, new_n10553, new_n10554, new_n10555, new_n10556, new_n10557, new_n10558, new_n10559, new_n10560, new_n10561, new_n10562, new_n10563, new_n10564, new_n10565, new_n10566, new_n10567, new_n10568, new_n10569, new_n10570, new_n10571, new_n10572, new_n10573, new_n10574, new_n10575, new_n10576, new_n10577, new_n10578, new_n10579, new_n10580, new_n10581, new_n10582, new_n10583, new_n10584, new_n10585, new_n10586, new_n10587, new_n10588, new_n10589, new_n10590, new_n10591, new_n10592, new_n10593, new_n10594, new_n10595, new_n10596, new_n10597, new_n10598, new_n10599, new_n10600, new_n10601, new_n10602, new_n10603, new_n10604, new_n10605, new_n10606, new_n10607, new_n10608, new_n10609, new_n10610, new_n10611, new_n10612, new_n10613, new_n10614, new_n10615, new_n10616, new_n10617, new_n10618, new_n10619, new_n10620, new_n10621, new_n10622, new_n10623, new_n10624, new_n10625, new_n10626, new_n10627, new_n10628, new_n10629, new_n10630, new_n10631, new_n10632, new_n10633, new_n10634, new_n10635, new_n10636, new_n10637, new_n10638, new_n10639, new_n10640, new_n10641, new_n10642, new_n10643, new_n10644, new_n10645, new_n10646, new_n10647, new_n10648, new_n10649, new_n10650, new_n10651, new_n10652, new_n10653, new_n10654, new_n10655, new_n10656, new_n10657, new_n10658, new_n10659, new_n10660, new_n10661, new_n10662, new_n10663, new_n10664, new_n10665, new_n10666, new_n10667, new_n10668, new_n10669, new_n10670, new_n10671, new_n10672, new_n10673, new_n10674, new_n10675, new_n10676, new_n10677, new_n10678, new_n10679, new_n10680, new_n10681, new_n10682, new_n10683, new_n10684, new_n10685, new_n10686, new_n10687, new_n10688, new_n10689, new_n10690, new_n10691, new_n10692, new_n10693, new_n10694, new_n10695, new_n10696, new_n10697, new_n10698, new_n10699, new_n10700, new_n10701, new_n10702, new_n10703, new_n10704, new_n10705, new_n10706, new_n10707, new_n10708, new_n10709, new_n10710, new_n10711, new_n10712, new_n10713, new_n10714, new_n10715, new_n10716, new_n10717, new_n10718, new_n10719, new_n10720, new_n10721, new_n10722, new_n10723, new_n10724, new_n10725, new_n10726, new_n10727, new_n10728, new_n10729, new_n10730, new_n10731, new_n10732, new_n10733, new_n10734, new_n10735, new_n10736, new_n10737, new_n10738, new_n10739, new_n10740, new_n10741, new_n10742, new_n10743, new_n10744, new_n10745, new_n10746, new_n10747, new_n10748, new_n10749, new_n10750, new_n10751, new_n10752, new_n10753, new_n10754, new_n10755, new_n10756, new_n10757, new_n10758, new_n10759, new_n10760, new_n10761, new_n10762, new_n10763, new_n10764, new_n10765, new_n10766, new_n10767, new_n10768, new_n10769, new_n10770, new_n10771, new_n10772, new_n10773, new_n10774, new_n10775, new_n10776, new_n10777, new_n10778, new_n10779, new_n10780, new_n10781, new_n10782, new_n10783, new_n10784, new_n10785, new_n10786, new_n10787, new_n10788, new_n10789, new_n10790, new_n10791, new_n10792, new_n10793, new_n10794, new_n10795, new_n10796, new_n10797, new_n10798, new_n10799, new_n10800, new_n10801, new_n10802, new_n10803, new_n10804, new_n10805, new_n10806, new_n10807, new_n10808, new_n10809, new_n10810, new_n10811, new_n10812, new_n10813, new_n10814, new_n10815, new_n10816, new_n10817, new_n10818, new_n10819, new_n10820, new_n10821, new_n10822, new_n10823, new_n10824, new_n10825, new_n10826, new_n10827, new_n10828, new_n10829, new_n10830, new_n10831, new_n10832, new_n10833, new_n10834, new_n10835, new_n10836, new_n10837, new_n10838, new_n10839, new_n10840, new_n10841, new_n10842, new_n10843, new_n10844, new_n10845, new_n10846, new_n10847, new_n10848, new_n10849, new_n10850, new_n10851, new_n10852, new_n10853, new_n10854, new_n10855, new_n10856, new_n10857, new_n10858, new_n10859, new_n10860, new_n10861, new_n10862, new_n10863, new_n10864, new_n10865, new_n10866, new_n10867, new_n10868, new_n10869, new_n10870, new_n10871, new_n10872, new_n10873, new_n10874, new_n10875, new_n10876, new_n10877, new_n10878, new_n10879, new_n10880, new_n10881, new_n10882, new_n10883, new_n10884, new_n10885, new_n10886, new_n10887, new_n10888, new_n10889, new_n10890, new_n10891, new_n10892, new_n10893, new_n10894, new_n10895, new_n10896, new_n10897, new_n10898, new_n10899, new_n10900, new_n10901, new_n10902, new_n10903, new_n10904, new_n10905, new_n10906, new_n10907, new_n10908, new_n10909, new_n10910, new_n10911, new_n10912, new_n10913, new_n10914, new_n10915, new_n10916, new_n10917, new_n10918, new_n10919, new_n10920, new_n10921, new_n10922, new_n10923, new_n10924, new_n10925, new_n10926, new_n10927, new_n10928, new_n10929, new_n10930, new_n10931, new_n10932, new_n10933, new_n10934, new_n10935, new_n10936, new_n10937, new_n10938, new_n10939, new_n10940, new_n10941, new_n10942, new_n10943, new_n10944, new_n10945, new_n10946, new_n10947, new_n10948, new_n10949, new_n10950, new_n10951, new_n10952, new_n10953, new_n10954, new_n10955, new_n10956, new_n10957, new_n10958, new_n10959, new_n10960, new_n10961, new_n10962, new_n10963, new_n10964, new_n10965, new_n10966, new_n10967, new_n10968, new_n10969, new_n10970, new_n10971, new_n10972, new_n10973, new_n10974, new_n10975, new_n10976, new_n10977, new_n10978, new_n10979, new_n10980, new_n10981, new_n10982, new_n10983, new_n10984, new_n10985, new_n10986, new_n10987, new_n10988, new_n10989, new_n10990, new_n10991, new_n10992, new_n10993, new_n10994, new_n10995, new_n10996, new_n10997, new_n10998, new_n10999, new_n11000, new_n11001, new_n11002, new_n11003, new_n11004, new_n11005, new_n11006, new_n11007, new_n11008, new_n11009, new_n11010, new_n11011, new_n11012, new_n11013, new_n11014, new_n11015, new_n11016, new_n11017, new_n11018, new_n11019, new_n11020, new_n11021, new_n11022, new_n11023, new_n11024, new_n11025, new_n11026, new_n11027, new_n11028, new_n11029, new_n11030, new_n11031, new_n11032, new_n11033, new_n11034, new_n11035, new_n11036, new_n11037, new_n11038, new_n11039, new_n11040, new_n11041, new_n11042, new_n11043, new_n11044, new_n11045, new_n11046, new_n11047, new_n11048, new_n11049, new_n11050, new_n11051, new_n11052, new_n11053, new_n11054, new_n11055, new_n11056, new_n11057, new_n11058, new_n11059, new_n11060, new_n11061, new_n11062, new_n11063, new_n11064, new_n11065, new_n11066, new_n11067, new_n11068, new_n11069, new_n11070, new_n11071, new_n11072, new_n11073, new_n11074, new_n11075, new_n11076, new_n11077, new_n11078, new_n11079, new_n11080, new_n11081, new_n11082, new_n11083, new_n11084, new_n11085, new_n11086, new_n11087, new_n11088, new_n11089, new_n11090, new_n11091, new_n11092, new_n11093, new_n11094, new_n11095, new_n11096, new_n11097, new_n11098, new_n11099, new_n11100, new_n11101, new_n11102, new_n11103, new_n11104, new_n11105, new_n11106, new_n11107, new_n11108, new_n11109, new_n11110, new_n11111, new_n11112, new_n11113, new_n11114, new_n11115, new_n11116, new_n11117, new_n11118, new_n11119, new_n11120, new_n11121, new_n11122, new_n11123, new_n11124, new_n11125, new_n11126, new_n11127, new_n11128, new_n11129, new_n11130, new_n11131, new_n11132, new_n11133, new_n11134, new_n11135, new_n11136, new_n11137, new_n11138, new_n11139, new_n11140, new_n11141, new_n11142, new_n11143, new_n11144, new_n11145, new_n11146, new_n11147, new_n11148, new_n11149, new_n11150, new_n11151, new_n11152, new_n11153, new_n11154, new_n11155, new_n11156, new_n11157, new_n11158, new_n11159, new_n11160, new_n11161, new_n11162, new_n11163, new_n11164, new_n11165, new_n11166, new_n11167, new_n11168, new_n11169, new_n11170, new_n11171, new_n11172, new_n11173, new_n11174, new_n11175, new_n11176, new_n11177, new_n11178, new_n11179, new_n11180, new_n11181, new_n11182, new_n11183, new_n11184, new_n11185, new_n11186, new_n11187, new_n11188, new_n11189, new_n11190, new_n11191, new_n11192, new_n11193, new_n11194, new_n11195, new_n11196, new_n11197, new_n11198, new_n11199, new_n11200, new_n11201, new_n11202, new_n11203, new_n11204, new_n11205, new_n11206, new_n11207, new_n11208, new_n11209, new_n11210, new_n11211, new_n11212, new_n11213, new_n11214, new_n11215, new_n11216, new_n11217, new_n11218, new_n11219, new_n11220, new_n11221, new_n11222, new_n11223, new_n11224, new_n11225, new_n11226, new_n11227, new_n11228, new_n11229, new_n11230, new_n11231, new_n11232, new_n11233, new_n11234, new_n11235, new_n11236, new_n11237, new_n11238, new_n11239, new_n11240, new_n11241, new_n11242, new_n11243, new_n11244, new_n11245, new_n11246, new_n11247, new_n11248, new_n11249, new_n11250, new_n11251, new_n11252, new_n11253, new_n11254, new_n11255, new_n11256, new_n11257, new_n11258, new_n11259, new_n11260, new_n11261, new_n11262, new_n11263, new_n11264, new_n11265, new_n11266, new_n11267, new_n11268, new_n11269, new_n11270, new_n11271, new_n11272, new_n11273, new_n11274, new_n11275, new_n11276, new_n11277, new_n11278, new_n11279, new_n11280, new_n11281, new_n11282, new_n11283, new_n11284, new_n11285, new_n11286, new_n11287, new_n11288, new_n11289, new_n11290, new_n11291, new_n11292, new_n11293, new_n11294, new_n11295, new_n11296, new_n11297, new_n11298, new_n11299, new_n11300, new_n11301, new_n11302, new_n11303, new_n11304, new_n11305, new_n11306, new_n11307, new_n11308, new_n11309, new_n11310, new_n11311, new_n11312, new_n11313, new_n11314, new_n11315, new_n11316, new_n11317, new_n11318, new_n11319, new_n11320, new_n11321, new_n11322, new_n11323, new_n11324, new_n11325, new_n11326, new_n11327, new_n11328, new_n11329, new_n11330, new_n11331, new_n11332, new_n11333, new_n11334, new_n11335, new_n11336, new_n11337, new_n11338, new_n11339, new_n11340, new_n11341, new_n11342, new_n11343, new_n11344, new_n11345, new_n11346, new_n11347, new_n11348, new_n11349, new_n11350, new_n11351, new_n11352, new_n11353, new_n11354, new_n11355, new_n11356, new_n11357, new_n11358, new_n11359, new_n11360, new_n11361, new_n11362, new_n11363, new_n11364, new_n11365, new_n11366, new_n11367, new_n11368, new_n11369, new_n11370, new_n11371, new_n11372, new_n11373, new_n11374, new_n11375, new_n11376, new_n11377, new_n11378, new_n11379, new_n11380, new_n11381, new_n11382, new_n11383, new_n11384, new_n11385, new_n11386, new_n11387, new_n11388, new_n11389, new_n11390, new_n11391, new_n11392, new_n11393, new_n11394, new_n11395, new_n11396, new_n11397, new_n11398, new_n11399, new_n11400, new_n11401, new_n11402, new_n11403, new_n11404, new_n11405, new_n11406, new_n11407, new_n11408, new_n11409, new_n11410, new_n11411, new_n11412, new_n11413, new_n11414, new_n11415, new_n11416, new_n11417, new_n11418, new_n11419, new_n11420, new_n11421, new_n11422, new_n11423, new_n11424, new_n11425, new_n11426, new_n11427, new_n11428, new_n11429, new_n11430, new_n11431, new_n11432, new_n11433, new_n11434, new_n11435, new_n11436, new_n11437, new_n11438, new_n11439, new_n11440, new_n11441, new_n11442, new_n11443, new_n11444, new_n11445, new_n11446, new_n11447, new_n11448, new_n11449, new_n11450, new_n11451, new_n11452, new_n11453, new_n11454, new_n11455, new_n11456, new_n11457, new_n11458, new_n11459, new_n11460, new_n11461, new_n11462, new_n11463, new_n11464, new_n11465, new_n11466, new_n11467, new_n11468, new_n11469, new_n11470, new_n11471, new_n11472, new_n11473, new_n11474, new_n11475, new_n11476, new_n11477, new_n11478, new_n11479, new_n11480, new_n11481, new_n11482, new_n11483, new_n11484, new_n11485, new_n11486, new_n11487, new_n11488, new_n11489, new_n11490, new_n11491, new_n11492, new_n11493, new_n11494, new_n11495, new_n11496, new_n11497, new_n11498, new_n11499, new_n11500, new_n11501, new_n11502, new_n11503, new_n11504, new_n11505, new_n11506, new_n11507, new_n11508, new_n11509, new_n11510, new_n11511, new_n11512, new_n11513, new_n11514, new_n11515, new_n11516, new_n11517, new_n11518, new_n11519, new_n11520, new_n11521, new_n11522, new_n11523, new_n11524, new_n11525, new_n11526, new_n11527, new_n11528, new_n11529, new_n11530, new_n11531, new_n11532, new_n11533, new_n11534, new_n11535, new_n11536, new_n11537, new_n11538, new_n11539, new_n11540, new_n11541, new_n11542, new_n11543, new_n11544, new_n11545, new_n11546, new_n11547, new_n11548, new_n11549, new_n11550, new_n11551, new_n11552, new_n11553, new_n11554, new_n11555, new_n11556, new_n11557, new_n11558, new_n11559, new_n11560, new_n11561, new_n11562, new_n11563, new_n11564, new_n11565, new_n11566, new_n11567, new_n11568, new_n11569, new_n11570, new_n11571, new_n11572, new_n11573, new_n11574, new_n11575, new_n11576, new_n11577, new_n11578, new_n11579, new_n11580, new_n11581, new_n11582, new_n11583, new_n11584, new_n11585, new_n11586, new_n11587, new_n11588, new_n11589, new_n11590, new_n11591, new_n11592, new_n11593, new_n11594, new_n11595, new_n11596, new_n11597, new_n11598, new_n11599, new_n11600, new_n11601, new_n11602, new_n11603, new_n11604, new_n11605, new_n11606, new_n11607, new_n11608, new_n11609, new_n11610, new_n11611, new_n11612, new_n11613, new_n11614, new_n11615, new_n11616, new_n11617, new_n11618, new_n11619, new_n11620, new_n11621, new_n11622, new_n11623, new_n11624, new_n11625, new_n11626, new_n11627, new_n11628, new_n11629, new_n11630, new_n11631, new_n11632, new_n11633, new_n11634, new_n11635, new_n11636, new_n11637, new_n11638, new_n11639, new_n11640, new_n11641, new_n11642, new_n11643, new_n11644, new_n11645, new_n11646, new_n11647, new_n11648, new_n11649, new_n11650, new_n11651, new_n11652, new_n11653, new_n11654, new_n11655, new_n11656, new_n11657, new_n11658, new_n11659, new_n11660, new_n11661, new_n11662, new_n11663, new_n11664, new_n11665, new_n11666, new_n11667, new_n11668, new_n11669, new_n11670, new_n11671, new_n11672, new_n11673, new_n11674, new_n11675, new_n11676, new_n11677, new_n11678, new_n11679, new_n11680, new_n11681, new_n11682, new_n11683, new_n11684, new_n11685, new_n11686, new_n11687, new_n11688, new_n11689, new_n11690, new_n11691, new_n11692, new_n11693, new_n11694, new_n11695, new_n11696, new_n11697, new_n11698, new_n11699, new_n11700, new_n11701, new_n11702, new_n11703, new_n11704, new_n11705, new_n11706, new_n11707, new_n11708, new_n11709, new_n11710, new_n11711, new_n11712, new_n11713, new_n11714, new_n11715, new_n11716, new_n11717, new_n11718, new_n11719, new_n11720, new_n11721, new_n11722, new_n11723, new_n11724, new_n11725, new_n11726, new_n11727, new_n11728, new_n11729, new_n11730, new_n11731, new_n11732, new_n11733, new_n11734, new_n11735, new_n11736, new_n11737, new_n11738, new_n11739, new_n11740, new_n11741, new_n11742, new_n11743, new_n11744, new_n11745, new_n11746, new_n11747, new_n11748, new_n11749, new_n11750, new_n11751, new_n11752, new_n11753, new_n11754, new_n11755, new_n11756, new_n11757, new_n11758, new_n11759, new_n11760, new_n11761, new_n11762, new_n11763, new_n11764, new_n11765, new_n11766, new_n11767, new_n11768, new_n11769, new_n11770, new_n11771, new_n11772, new_n11773, new_n11774, new_n11775, new_n11776, new_n11777, new_n11778, new_n11779, new_n11780, new_n11781, new_n11782, new_n11783, new_n11784, new_n11785, new_n11786, new_n11787, new_n11788, new_n11789, new_n11790, new_n11791, new_n11792, new_n11793, new_n11794, new_n11795, new_n11796, new_n11797, new_n11798, new_n11799, new_n11800, new_n11801, new_n11802, new_n11803, new_n11804, new_n11805, new_n11806, new_n11807, new_n11808, new_n11809, new_n11810, new_n11811, new_n11812, new_n11813, new_n11814, new_n11815, new_n11816, new_n11817, new_n11818, new_n11819, new_n11820, new_n11821, new_n11822, new_n11823, new_n11824, new_n11825, new_n11826, new_n11827, new_n11828, new_n11829, new_n11830, new_n11831, new_n11832, new_n11833, new_n11834, new_n11835, new_n11836, new_n11837, new_n11838, new_n11839, new_n11840, new_n11841, new_n11842, new_n11843, new_n11844, new_n11845, new_n11846, new_n11847, new_n11848, new_n11849, new_n11850, new_n11851, new_n11852, new_n11853, new_n11854, new_n11855, new_n11856, new_n11857, new_n11858, new_n11859, new_n11860, new_n11861, new_n11862, new_n11863, new_n11864, new_n11865, new_n11866, new_n11867, new_n11868, new_n11869, new_n11870, new_n11871, new_n11872, new_n11873, new_n11874, new_n11875, new_n11876, new_n11877, new_n11878, new_n11879, new_n11880, new_n11881, new_n11882, new_n11883, new_n11884, new_n11885, new_n11886, new_n11887, new_n11888, new_n11889, new_n11890, new_n11891, new_n11892, new_n11893, new_n11894, new_n11895, new_n11896, new_n11897, new_n11898, new_n11899, new_n11900, new_n11901, new_n11902, new_n11903, new_n11904, new_n11905, new_n11906, new_n11907, new_n11908, new_n11909, new_n11910, new_n11911, new_n11912, new_n11913, new_n11914, new_n11915, new_n11916, new_n11917, new_n11918, new_n11919, new_n11920, new_n11921, new_n11922, new_n11923, new_n11924, new_n11925, new_n11926, new_n11927, new_n11928, new_n11929, new_n11930, new_n11931, new_n11932, new_n11933, new_n11934, new_n11935, new_n11936, new_n11937, new_n11938, new_n11939, new_n11940, new_n11941, new_n11942, new_n11943, new_n11944, new_n11945, new_n11946, new_n11947, new_n11948, new_n11949, new_n11950, new_n11951, new_n11952, new_n11953, new_n11954, new_n11955, new_n11956, new_n11957, new_n11958, new_n11959, new_n11960, new_n11961, new_n11962, new_n11963, new_n11964, new_n11965, new_n11966, new_n11967, new_n11968, new_n11969, new_n11970, new_n11971, new_n11972, new_n11973, new_n11974, new_n11975, new_n11976, new_n11977, new_n11978, new_n11979, new_n11980, new_n11981, new_n11982, new_n11983, new_n11984, new_n11985, new_n11986, new_n11987, new_n11988, new_n11989, new_n11990, new_n11991, new_n11992, new_n11993, new_n11994, new_n11995, new_n11996, new_n11997, new_n11998, new_n11999, new_n12000, new_n12001, new_n12002, new_n12003, new_n12004, new_n12005, new_n12006, new_n12007, new_n12008, new_n12009, new_n12010, new_n12011, new_n12012, new_n12013, new_n12014, new_n12015, new_n12016, new_n12017, new_n12018, new_n12019, new_n12020, new_n12021, new_n12022, new_n12023, new_n12024, new_n12025, new_n12026, new_n12027, new_n12028, new_n12029, new_n12030, new_n12031, new_n12032, new_n12033, new_n12034, new_n12035, new_n12036, new_n12037, new_n12038, new_n12039, new_n12040, new_n12041, new_n12042, new_n12043, new_n12044, new_n12045, new_n12046, new_n12047, new_n12048, new_n12049, new_n12050, new_n12051, new_n12052, new_n12053, new_n12054, new_n12055, new_n12056, new_n12057, new_n12058, new_n12059, new_n12060, new_n12061, new_n12062, new_n12063, new_n12064, new_n12065, new_n12066, new_n12067, new_n12068, new_n12069, new_n12070, new_n12071, new_n12072, new_n12073, new_n12074, new_n12075, new_n12076, new_n12077, new_n12078, new_n12079, new_n12080, new_n12081, new_n12082, new_n12083, new_n12084, new_n12085, new_n12086, new_n12087, new_n12088, new_n12089, new_n12090, new_n12091, new_n12092, new_n12093, new_n12094, new_n12095, new_n12096, new_n12097, new_n12098, new_n12099, new_n12100, new_n12101, new_n12102, new_n12103, new_n12104, new_n12105, new_n12106, new_n12107, new_n12108, new_n12109, new_n12110, new_n12111, new_n12112, new_n12113, new_n12114, new_n12115, new_n12116, new_n12117, new_n12118, new_n12119, new_n12120, new_n12121, new_n12122, new_n12123, new_n12124, new_n12125, new_n12126, new_n12127, new_n12128, new_n12129, new_n12130, new_n12131, new_n12132, new_n12133, new_n12134, new_n12135, new_n12136, new_n12137, new_n12138, new_n12139, new_n12140, new_n12141, new_n12142, new_n12143, new_n12144, new_n12145, new_n12146, new_n12147, new_n12148, new_n12149, new_n12150, new_n12151, new_n12152, new_n12153, new_n12154, new_n12155, new_n12156, new_n12157, new_n12158, new_n12159, new_n12160, new_n12161, new_n12162, new_n12163, new_n12164, new_n12165, new_n12166, new_n12167, new_n12168, new_n12169, new_n12170, new_n12171, new_n12172, new_n12173, new_n12174, new_n12175, new_n12176, new_n12177, new_n12178, new_n12179, new_n12180, new_n12181, new_n12182, new_n12183, new_n12184, new_n12185, new_n12186, new_n12187, new_n12188, new_n12189, new_n12190, new_n12191, new_n12192, new_n12193, new_n12194, new_n12195, new_n12196, new_n12197, new_n12198, new_n12199, new_n12200, new_n12201, new_n12202, new_n12203, new_n12204, new_n12205, new_n12206, new_n12207, new_n12208, new_n12209, new_n12210, new_n12211, new_n12212, new_n12213, new_n12214, new_n12215, new_n12216, new_n12217, new_n12218, new_n12219, new_n12220, new_n12221, new_n12222, new_n12223, new_n12224, new_n12225, new_n12226, new_n12227, new_n12228, new_n12229, new_n12230, new_n12231, new_n12232, new_n12233, new_n12234, new_n12235, new_n12236, new_n12237, new_n12238, new_n12239, new_n12240, new_n12241, new_n12242, new_n12243, new_n12244, new_n12245, new_n12246, new_n12247, new_n12248, new_n12249, new_n12250, new_n12251, new_n12252, new_n12253, new_n12254, new_n12255, new_n12256, new_n12257, new_n12258, new_n12259, new_n12260, new_n12261, new_n12262, new_n12263, new_n12264, new_n12265, new_n12266, new_n12267, new_n12268, new_n12269, new_n12270, new_n12271, new_n12272, new_n12273, new_n12274, new_n12275, new_n12276, new_n12277, new_n12278, new_n12279, new_n12280, new_n12281, new_n12282, new_n12283, new_n12284, new_n12285, new_n12286, new_n12287, new_n12288, new_n12289, new_n12290, new_n12291, new_n12292, new_n12293, new_n12294, new_n12295, new_n12296, new_n12297, new_n12298, new_n12299, new_n12300, new_n12301, new_n12302, new_n12303, new_n12304, new_n12305, new_n12306, new_n12307, new_n12308, new_n12309, new_n12310, new_n12311, new_n12312, new_n12313, new_n12314, new_n12315, new_n12316, new_n12317, new_n12318, new_n12319, new_n12320, new_n12321, new_n12322, new_n12323, new_n12324, new_n12325, new_n12326, new_n12327, new_n12328, new_n12329, new_n12330, new_n12331, new_n12332, new_n12333, new_n12334, new_n12335, new_n12336, new_n12337, new_n12338, new_n12339, new_n12340, new_n12341, new_n12342, new_n12343, new_n12344, new_n12345, new_n12346, new_n12347, new_n12348, new_n12349, new_n12350, new_n12351, new_n12352, new_n12353, new_n12354, new_n12355, new_n12356, new_n12357, new_n12358, new_n12359, new_n12360, new_n12361, new_n12362, new_n12363, new_n12364, new_n12365, new_n12366, new_n12367, new_n12368, new_n12369, new_n12370, new_n12371, new_n12372, new_n12373, new_n12374, new_n12375, new_n12376, new_n12377, new_n12378, new_n12379, new_n12380, new_n12381, new_n12382, new_n12383, new_n12384, new_n12385, new_n12386, new_n12387, new_n12388, new_n12389, new_n12390, new_n12391, new_n12392, new_n12393, new_n12394, new_n12395, new_n12396, new_n12397, new_n12398, new_n12399, new_n12400, new_n12401, new_n12402, new_n12403, new_n12404, new_n12405, new_n12406, new_n12407, new_n12408, new_n12409, new_n12410, new_n12411, new_n12412, new_n12413, new_n12414, new_n12415, new_n12416, new_n12417, new_n12418, new_n12419, new_n12420, new_n12421, new_n12422, new_n12423, new_n12424, new_n12425, new_n12426, new_n12427, new_n12428, new_n12429, new_n12430, new_n12431, new_n12432, new_n12433, new_n12434, new_n12435, new_n12436, new_n12437, new_n12438, new_n12439, new_n12440, new_n12441, new_n12442, new_n12443, new_n12444, new_n12445, new_n12446, new_n12447, new_n12448, new_n12449, new_n12450, new_n12451, new_n12452, new_n12453, new_n12454, new_n12455, new_n12456, new_n12457, new_n12458, new_n12459, new_n12460, new_n12461, new_n12462, new_n12463, new_n12464, new_n12465, new_n12466, new_n12467, new_n12468, new_n12469, new_n12470, new_n12471, new_n12472, new_n12473, new_n12474, new_n12475, new_n12476, new_n12477, new_n12478, new_n12479, new_n12480, new_n12481, new_n12482, new_n12483, new_n12484, new_n12485, new_n12486, new_n12487, new_n12488, new_n12489, new_n12490, new_n12491, new_n12492, new_n12493, new_n12494, new_n12495, new_n12496, new_n12497, new_n12498, new_n12499, new_n12500, new_n12501, new_n12502, new_n12503, new_n12504, new_n12505, new_n12506, new_n12507, new_n12508, new_n12509, new_n12510, new_n12511, new_n12512, new_n12513, new_n12514, new_n12515, new_n12516, new_n12517, new_n12518, new_n12519, new_n12520, new_n12521, new_n12522, new_n12523, new_n12524, new_n12525, new_n12526, new_n12527, new_n12528, new_n12529, new_n12530, new_n12531, new_n12532, new_n12533, new_n12534, new_n12535, new_n12536, new_n12537, new_n12538, new_n12539, new_n12540, new_n12541, new_n12542, new_n12543, new_n12544, new_n12545, new_n12546, new_n12547, new_n12548, new_n12549, new_n12550, new_n12551, new_n12552, new_n12553, new_n12554, new_n12555, new_n12556, new_n12557, new_n12558, new_n12559, new_n12560, new_n12561, new_n12562, new_n12563, new_n12564, new_n12565, new_n12566, new_n12567, new_n12568, new_n12569, new_n12570, new_n12571, new_n12572, new_n12573, new_n12574, new_n12575, new_n12576, new_n12577, new_n12578, new_n12579, new_n12580, new_n12581, new_n12582, new_n12583, new_n12584, new_n12585, new_n12586, new_n12587, new_n12588, new_n12589, new_n12590, new_n12591, new_n12592, new_n12593, new_n12594, new_n12595, new_n12596, new_n12597, new_n12598, new_n12599, new_n12600, new_n12601, new_n12602, new_n12603, new_n12604, new_n12605, new_n12606, new_n12607, new_n12608, new_n12609, new_n12610, new_n12611, new_n12612, new_n12613, new_n12614, new_n12615, new_n12616, new_n12617, new_n12618, new_n12619, new_n12620, new_n12621, new_n12622, new_n12623, new_n12624, new_n12625, new_n12626, new_n12627, new_n12628, new_n12629, new_n12630, new_n12631, new_n12632, new_n12633, new_n12634, new_n12635, new_n12636, new_n12637, new_n12638, new_n12639, new_n12640, new_n12641, new_n12642, new_n12643, new_n12644, new_n12645, new_n12646, new_n12647, new_n12648, new_n12649, new_n12650, new_n12651, new_n12652, new_n12653, new_n12654, new_n12655, new_n12656, new_n12657, new_n12658, new_n12659, new_n12660, new_n12661, new_n12662, new_n12663, new_n12664, new_n12665, new_n12666, new_n12667, new_n12668, new_n12669, new_n12670, new_n12671, new_n12672, new_n12673, new_n12674, new_n12675, new_n12676, new_n12677, new_n12678, new_n12679, new_n12680, new_n12681, new_n12682, new_n12683, new_n12684, new_n12685, new_n12686, new_n12687, new_n12688, new_n12689, new_n12690, new_n12691, new_n12692, new_n12693, new_n12694, new_n12695, new_n12696, new_n12697, new_n12698, new_n12699, new_n12700, new_n12701, new_n12702, new_n12703, new_n12704, new_n12705, new_n12706, new_n12707, new_n12708, new_n12709, new_n12710, new_n12711, new_n12712, new_n12713, new_n12714, new_n12715, new_n12716, new_n12717, new_n12718, new_n12719, new_n12720, new_n12721, new_n12722, new_n12723, new_n12724, new_n12725, new_n12726, new_n12727, new_n12728, new_n12729, new_n12730, new_n12731, new_n12732, new_n12733, new_n12734, new_n12735, new_n12736, new_n12737, new_n12738, new_n12739, new_n12740, new_n12741, new_n12742, new_n12743, new_n12744, new_n12745, new_n12746, new_n12747, new_n12748, new_n12749, new_n12750, new_n12751, new_n12752, new_n12753, new_n12754, new_n12755, new_n12756, new_n12757, new_n12758, new_n12759, new_n12760, new_n12761, new_n12762, new_n12763, new_n12764, new_n12765, new_n12766, new_n12767, new_n12768, new_n12769, new_n12770, new_n12771, new_n12772, new_n12773, new_n12774, new_n12775, new_n12776, new_n12777, new_n12778, new_n12779, new_n12780, new_n12781, new_n12782, new_n12783, new_n12784, new_n12785, new_n12786, new_n12787, new_n12788, new_n12789, new_n12790, new_n12791, new_n12792, new_n12793, new_n12794, new_n12795, new_n12796, new_n12797, new_n12798, new_n12799, new_n12800, new_n12801, new_n12802, new_n12803, new_n12804, new_n12805, new_n12806, new_n12807, new_n12808, new_n12809, new_n12810, new_n12811, new_n12812, new_n12813, new_n12814, new_n12815, new_n12816, new_n12817, new_n12818, new_n12819, new_n12820, new_n12821, new_n12822, new_n12823, new_n12824, new_n12825, new_n12826, new_n12827, new_n12828, new_n12829, new_n12830, new_n12831, new_n12832, new_n12833, new_n12834, new_n12835, new_n12836, new_n12837, new_n12838, new_n12839, new_n12840, new_n12841, new_n12842, new_n12843, new_n12844, new_n12845, new_n12846, new_n12847, new_n12848, new_n12849, new_n12850, new_n12851, new_n12852, new_n12853, new_n12854, new_n12855, new_n12856, new_n12857, new_n12858, new_n12859, new_n12860, new_n12861, new_n12862, new_n12863, new_n12864, new_n12865, new_n12866, new_n12867, new_n12868, new_n12869, new_n12870, new_n12871, new_n12872, new_n12873, new_n12874, new_n12875, new_n12876, new_n12877, new_n12878, new_n12879, new_n12880, new_n12881, new_n12882, new_n12883, new_n12884, new_n12885, new_n12886, new_n12887, new_n12888, new_n12889, new_n12890, new_n12891, new_n12892, new_n12893, new_n12894, new_n12895, new_n12896, new_n12897, new_n12898, new_n12899, new_n12900, new_n12901, new_n12902, new_n12903, new_n12904, new_n12905, new_n12906, new_n12907, new_n12908, new_n12909, new_n12910, new_n12911, new_n12912, new_n12913, new_n12914, new_n12915, new_n12916, new_n12917, new_n12918, new_n12919, new_n12920, new_n12921, new_n12922, new_n12923, new_n12924, new_n12925, new_n12926, new_n12927, new_n12928, new_n12929, new_n12930, new_n12931, new_n12932, new_n12933, new_n12934, new_n12935, new_n12936, new_n12937, new_n12938, new_n12939, new_n12940, new_n12941, new_n12942, new_n12943, new_n12944, new_n12945, new_n12946, new_n12947, new_n12948, new_n12949, new_n12950, new_n12951, new_n12952, new_n12953, new_n12954, new_n12955, new_n12956, new_n12957, new_n12958, new_n12959, new_n12960, new_n12961, new_n12962, new_n12963, new_n12964, new_n12965, new_n12966, new_n12967, new_n12968, new_n12969, new_n12970, new_n12971, new_n12972, new_n12973, new_n12974, new_n12975, new_n12976, new_n12977, new_n12978, new_n12979, new_n12980, new_n12981, new_n12982, new_n12983, new_n12984, new_n12985, new_n12986, new_n12987, new_n12988, new_n12989, new_n12990, new_n12991, new_n12992, new_n12993, new_n12994, new_n12995, new_n12996, new_n12997, new_n12998, new_n12999, new_n13000, new_n13001, new_n13002, new_n13003, new_n13004, new_n13005, new_n13006, new_n13007, new_n13008, new_n13009, new_n13010, new_n13011, new_n13012, new_n13013, new_n13014, new_n13015, new_n13016, new_n13017, new_n13018, new_n13019, new_n13020, new_n13021, new_n13022, new_n13023, new_n13024, new_n13025, new_n13026, new_n13027, new_n13028, new_n13029, new_n13030, new_n13031, new_n13032, new_n13033, new_n13034, new_n13035, new_n13036, new_n13037, new_n13038, new_n13039, new_n13040, new_n13041, new_n13042, new_n13043, new_n13044, new_n13045, new_n13046, new_n13047, new_n13048, new_n13049, new_n13050, new_n13051, new_n13052, new_n13053, new_n13054, new_n13055, new_n13056, new_n13057, new_n13058, new_n13059, new_n13060, new_n13061, new_n13062, new_n13063, new_n13064, new_n13065, new_n13066, new_n13067, new_n13068, new_n13069, new_n13070, new_n13071, new_n13072, new_n13073, new_n13074, new_n13075, new_n13076, new_n13077, new_n13078, new_n13079, new_n13080, new_n13081, new_n13082, new_n13083, new_n13084, new_n13085, new_n13086, new_n13087, new_n13088, new_n13089, new_n13090, new_n13091, new_n13092, new_n13093, new_n13094, new_n13095, new_n13096, new_n13097, new_n13098, new_n13099, new_n13100, new_n13101, new_n13102, new_n13103, new_n13104, new_n13105, new_n13106, new_n13107, new_n13108, new_n13109, new_n13110, new_n13111, new_n13112, new_n13113, new_n13114, new_n13115, new_n13116, new_n13117, new_n13118, new_n13119, new_n13120, new_n13121, new_n13122, new_n13123, new_n13124, new_n13125, new_n13126, new_n13127, new_n13128, new_n13129, new_n13130, new_n13131, new_n13132, new_n13133, new_n13134, new_n13135, new_n13136, new_n13137, new_n13138, new_n13139, new_n13140, new_n13141, new_n13142, new_n13143, new_n13144, new_n13145, new_n13146, new_n13147, new_n13148, new_n13149, new_n13150, new_n13151, new_n13152, new_n13153, new_n13154, new_n13155, new_n13156, new_n13157, new_n13158, new_n13159, new_n13160, new_n13161, new_n13162, new_n13163, new_n13164, new_n13165, new_n13166, new_n13167, new_n13168, new_n13169, new_n13170, new_n13171, new_n13172, new_n13173, new_n13174, new_n13175, new_n13176, new_n13177, new_n13178, new_n13179, new_n13180, new_n13181, new_n13182, new_n13183, new_n13184, new_n13185, new_n13186, new_n13187, new_n13188, new_n13189, new_n13190, new_n13191, new_n13192, new_n13193, new_n13194, new_n13195, new_n13196, new_n13197, new_n13198, new_n13199, new_n13200, new_n13201, new_n13202, new_n13203, new_n13204, new_n13205, new_n13206, new_n13207, new_n13208, new_n13209, new_n13210, new_n13211, new_n13212, new_n13213, new_n13214, new_n13215, new_n13216, new_n13217, new_n13218, new_n13219, new_n13220, new_n13221, new_n13222, new_n13223, new_n13224, new_n13225, new_n13226, new_n13227, new_n13228, new_n13229, new_n13230, new_n13231, new_n13232, new_n13233, new_n13234, new_n13235, new_n13236, new_n13237, new_n13238, new_n13239, new_n13240, new_n13241, new_n13242, new_n13243, new_n13244, new_n13245, new_n13246, new_n13247, new_n13248, new_n13249, new_n13250, new_n13251, new_n13252, new_n13253, new_n13254, new_n13255, new_n13256, new_n13257, new_n13258, new_n13259, new_n13260, new_n13261, new_n13262, new_n13263, new_n13264, new_n13265, new_n13266, new_n13267, new_n13268, new_n13269, new_n13270, new_n13271, new_n13272, new_n13273, new_n13274, new_n13275, new_n13276, new_n13277, new_n13278, new_n13279, new_n13280, new_n13281, new_n13282, new_n13283, new_n13284, new_n13285, new_n13286, new_n13287, new_n13288, new_n13289, new_n13290, new_n13291, new_n13292, new_n13293, new_n13294, new_n13295, new_n13296, new_n13297, new_n13298, new_n13299, new_n13300, new_n13301, new_n13302, new_n13303, new_n13304, new_n13305, new_n13306, new_n13307, new_n13308, new_n13309, new_n13310, new_n13311, new_n13312, new_n13313, new_n13314, new_n13315, new_n13316, new_n13317, new_n13318, new_n13319, new_n13320, new_n13321, new_n13322, new_n13323, new_n13324, new_n13325, new_n13326, new_n13327, new_n13328, new_n13329, new_n13330, new_n13331, new_n13332, new_n13333, new_n13334, new_n13335, new_n13336, new_n13337, new_n13338, new_n13339, new_n13340, new_n13341, new_n13342, new_n13343, new_n13344, new_n13345, new_n13346, new_n13347, new_n13348, new_n13349, new_n13350, new_n13351, new_n13352, new_n13353, new_n13354, new_n13355, new_n13356, new_n13357, new_n13358, new_n13359, new_n13360, new_n13361, new_n13362, new_n13363, new_n13364, new_n13365, new_n13366, new_n13367, new_n13368, new_n13369, new_n13370, new_n13371, new_n13372, new_n13373, new_n13374, new_n13375, new_n13376, new_n13377, new_n13378, new_n13379, new_n13380, new_n13381, new_n13382, new_n13383, new_n13384, new_n13385, new_n13386, new_n13387, new_n13388, new_n13389, new_n13390, new_n13391, new_n13392, new_n13393, new_n13394, new_n13395, new_n13396, new_n13397, new_n13398, new_n13399, new_n13400, new_n13401, new_n13402, new_n13403, new_n13404, new_n13405, new_n13406, new_n13407, new_n13408, new_n13409, new_n13410, new_n13411, new_n13412, new_n13413, new_n13414, new_n13415, new_n13416, new_n13417, new_n13418, new_n13419, new_n13420, new_n13421, new_n13422, new_n13423, new_n13424, new_n13425, new_n13426, new_n13427, new_n13428, new_n13429, new_n13430, new_n13431, new_n13432, new_n13433, new_n13434, new_n13435, new_n13436, new_n13437, new_n13438, new_n13439, new_n13440, new_n13441, new_n13442, new_n13443, new_n13444, new_n13445, new_n13446, new_n13447, new_n13448, new_n13449, new_n13450, new_n13451, new_n13452, new_n13453, new_n13454, new_n13455, new_n13456, new_n13457, new_n13458, new_n13459, new_n13460, new_n13461, new_n13462, new_n13463, new_n13464, new_n13465, new_n13466, new_n13467, new_n13468, new_n13469, new_n13470, new_n13471, new_n13472, new_n13473, new_n13474, new_n13475, new_n13476, new_n13477, new_n13478, new_n13479, new_n13480, new_n13481, new_n13482, new_n13483, new_n13484, new_n13485, new_n13486, new_n13487, new_n13488, new_n13489, new_n13490, new_n13491, new_n13492, new_n13493, new_n13494, new_n13495, new_n13496, new_n13497, new_n13498, new_n13499, new_n13500, new_n13501, new_n13502, new_n13503, new_n13504, new_n13505, new_n13506, new_n13507, new_n13508, new_n13509, new_n13510, new_n13511, new_n13512, new_n13513, new_n13514, new_n13515, new_n13516, new_n13517, new_n13518, new_n13519, new_n13520, new_n13521, new_n13522, new_n13523, new_n13524, new_n13525, new_n13526, new_n13527, new_n13528, new_n13529, new_n13530, new_n13531, new_n13532, new_n13533, new_n13534, new_n13535, new_n13536, new_n13537, new_n13538, new_n13539, new_n13540, new_n13541, new_n13542, new_n13543, new_n13544, new_n13545, new_n13546, new_n13547, new_n13548, new_n13549, new_n13550, new_n13551, new_n13552, new_n13553, new_n13554, new_n13555, new_n13556, new_n13557, new_n13558, new_n13559, new_n13560, new_n13561, new_n13562, new_n13563, new_n13564, new_n13565, new_n13566, new_n13567, new_n13568, new_n13569, new_n13570, new_n13571, new_n13572, new_n13573, new_n13574, new_n13575, new_n13576, new_n13577, new_n13578, new_n13579, new_n13580, new_n13581, new_n13582, new_n13583, new_n13584, new_n13585, new_n13586, new_n13587, new_n13588, new_n13589, new_n13590, new_n13591, new_n13592, new_n13593, new_n13594, new_n13595, new_n13596, new_n13597, new_n13598, new_n13599, new_n13600, new_n13601, new_n13602, new_n13603, new_n13604, new_n13605, new_n13606, new_n13607, new_n13608, new_n13609, new_n13610, new_n13611, new_n13612, new_n13613, new_n13614, new_n13615, new_n13616, new_n13617, new_n13618, new_n13619, new_n13620, new_n13621, new_n13622, new_n13623, new_n13624, new_n13625, new_n13626, new_n13627, new_n13628, new_n13629, new_n13630, new_n13631, new_n13632, new_n13633, new_n13634, new_n13635, new_n13636, new_n13637, new_n13638, new_n13639, new_n13640, new_n13641, new_n13642, new_n13643, new_n13644, new_n13645, new_n13646, new_n13647, new_n13648, new_n13649, new_n13650, new_n13651, new_n13652, new_n13653, new_n13654, new_n13655, new_n13656, new_n13657, new_n13658, new_n13659, new_n13660, new_n13661, new_n13662, new_n13663, new_n13664, new_n13665, new_n13666, new_n13667, new_n13668, new_n13669, new_n13670, new_n13671, new_n13672, new_n13673, new_n13674, new_n13675, new_n13676, new_n13677, new_n13678, new_n13679, new_n13680, new_n13681, new_n13682, new_n13683, new_n13684, new_n13685, new_n13686, new_n13687, new_n13688, new_n13689, new_n13690, new_n13691, new_n13692, new_n13693, new_n13694, new_n13695, new_n13696, new_n13697, new_n13698, new_n13699, new_n13700, new_n13701, new_n13702, new_n13703, new_n13704, new_n13705, new_n13706, new_n13707, new_n13708, new_n13709, new_n13710, new_n13711, new_n13712, new_n13713, new_n13714, new_n13715, new_n13716, new_n13717, new_n13718, new_n13719, new_n13720, new_n13721, new_n13722, new_n13723, new_n13724, new_n13725, new_n13726, new_n13727, new_n13728, new_n13729, new_n13730, new_n13731, new_n13732, new_n13733, new_n13734, new_n13735, new_n13736, new_n13737, new_n13738, new_n13739, new_n13740, new_n13741, new_n13742, new_n13743, new_n13744, new_n13745, new_n13746, new_n13747, new_n13748, new_n13749, new_n13750, new_n13751, new_n13752, new_n13753, new_n13754, new_n13755, new_n13756, new_n13757, new_n13758, new_n13759, new_n13760, new_n13761, new_n13762, new_n13763, new_n13764, new_n13765, new_n13766, new_n13767, new_n13768, new_n13769, new_n13770, new_n13771, new_n13772, new_n13773, new_n13774, new_n13775, new_n13776, new_n13777, new_n13778, new_n13779, new_n13780, new_n13781, new_n13782, new_n13783, new_n13784, new_n13785, new_n13786, new_n13787, new_n13788, new_n13789, new_n13790, new_n13791, new_n13792, new_n13793, new_n13794, new_n13795, new_n13796, new_n13797, new_n13798, new_n13799, new_n13800, new_n13801, new_n13802, new_n13803, new_n13804, new_n13805, new_n13806, new_n13807, new_n13808, new_n13809, new_n13810, new_n13811, new_n13812, new_n13813, new_n13814, new_n13815, new_n13816, new_n13817, new_n13818, new_n13819, new_n13820, new_n13821, new_n13822, new_n13823, new_n13824, new_n13825, new_n13826, new_n13827, new_n13828, new_n13829, new_n13830, new_n13831, new_n13832, new_n13833, new_n13834, new_n13835, new_n13836, new_n13837, new_n13838, new_n13839, new_n13840, new_n13841, new_n13842, new_n13843, new_n13844, new_n13845, new_n13846, new_n13847, new_n13848, new_n13849, new_n13850, new_n13851, new_n13852, new_n13853, new_n13854, new_n13855, new_n13856, new_n13857, new_n13858, new_n13859, new_n13860, new_n13861, new_n13862, new_n13863, new_n13864, new_n13865, new_n13866, new_n13867, new_n13868, new_n13869, new_n13870, new_n13871, new_n13872, new_n13873, new_n13874, new_n13875, new_n13876, new_n13877, new_n13878, new_n13879, new_n13880, new_n13881, new_n13882, new_n13883, new_n13884, new_n13885, new_n13886, new_n13887, new_n13888, new_n13889, new_n13890, new_n13891, new_n13892, new_n13893, new_n13894, new_n13895, new_n13896, new_n13897, new_n13898, new_n13899, new_n13900, new_n13901, new_n13902, new_n13903, new_n13904, new_n13905, new_n13906, new_n13907, new_n13908, new_n13909, new_n13910, new_n13911, new_n13912, new_n13913, new_n13914, new_n13915, new_n13916, new_n13917, new_n13918, new_n13919, new_n13920, new_n13921, new_n13922, new_n13923, new_n13924, new_n13925, new_n13926, new_n13927, new_n13928, new_n13929, new_n13930, new_n13931, new_n13932, new_n13933, new_n13934, new_n13935, new_n13936, new_n13937, new_n13938, new_n13939, new_n13940, new_n13941, new_n13942, new_n13943, new_n13944, new_n13945, new_n13946, new_n13947, new_n13948, new_n13949, new_n13950, new_n13951, new_n13952, new_n13953, new_n13954, new_n13955, new_n13956, new_n13957, new_n13958, new_n13959, new_n13960, new_n13961, new_n13962, new_n13963, new_n13964, new_n13965, new_n13966, new_n13967, new_n13968, new_n13969, new_n13970, new_n13971, new_n13972, new_n13973, new_n13974, new_n13975, new_n13976, new_n13977, new_n13978, new_n13979, new_n13980, new_n13981, new_n13982, new_n13983, new_n13984, new_n13985, new_n13986, new_n13987, new_n13988, new_n13989, new_n13990, new_n13991, new_n13992, new_n13993, new_n13994, new_n13995, new_n13996, new_n13997, new_n13998, new_n13999, new_n14000, new_n14001, new_n14002, new_n14003, new_n14004, new_n14005, new_n14006, new_n14007, new_n14008, new_n14009, new_n14010, new_n14011, new_n14012, new_n14013, new_n14014, new_n14015, new_n14016, new_n14017, new_n14018, new_n14019, new_n14020, new_n14021, new_n14022, new_n14023, new_n14024, new_n14025, new_n14026, new_n14027, new_n14028, new_n14029, new_n14030, new_n14031, new_n14032, new_n14033, new_n14034, new_n14035, new_n14036, new_n14037, new_n14038, new_n14039, new_n14040, new_n14041, new_n14042, new_n14043, new_n14044, new_n14045, new_n14046, new_n14047, new_n14048, new_n14049, new_n14050, new_n14051, new_n14052, new_n14053, new_n14054, new_n14055, new_n14056, new_n14057, new_n14058, new_n14059, new_n14060, new_n14061, new_n14062, new_n14063, new_n14064, new_n14065, new_n14066, new_n14067, new_n14068, new_n14069, new_n14070, new_n14071, new_n14072, new_n14073, new_n14074, new_n14075, new_n14076, new_n14077, new_n14078, new_n14079, new_n14080, new_n14081, new_n14082, new_n14083, new_n14084, new_n14085, new_n14086, new_n14087, new_n14088, new_n14089, new_n14090, new_n14091, new_n14092, new_n14093, new_n14094, new_n14095, new_n14096, new_n14097, new_n14098, new_n14099, new_n14100, new_n14101, new_n14102, new_n14103, new_n14104, new_n14105, new_n14106, new_n14107, new_n14108, new_n14109, new_n14110, new_n14111, new_n14112, new_n14113, new_n14114, new_n14115, new_n14116, new_n14117, new_n14118, new_n14119, new_n14120, new_n14121, new_n14122, new_n14123, new_n14124, new_n14125, new_n14126, new_n14127, new_n14128, new_n14129, new_n14130, new_n14131, new_n14132, new_n14133, new_n14134, new_n14135, new_n14136, new_n14137, new_n14138, new_n14139, new_n14140, new_n14141, new_n14142, new_n14143, new_n14144, new_n14145, new_n14146, new_n14147, new_n14148, new_n14149, new_n14150, new_n14151, new_n14152, new_n14153, new_n14154, new_n14155, new_n14156, new_n14157, new_n14158, new_n14159, new_n14160, new_n14161, new_n14162, new_n14163, new_n14164, new_n14165, new_n14166, new_n14167, new_n14168, new_n14169, new_n14170, new_n14171, new_n14172, new_n14173, new_n14174, new_n14175, new_n14176, new_n14177, new_n14178, new_n14179, new_n14180, new_n14181, new_n14182, new_n14183, new_n14184, new_n14185, new_n14186, new_n14187, new_n14188, new_n14189, new_n14190, new_n14191, new_n14192, new_n14193, new_n14194, new_n14195, new_n14196, new_n14197, new_n14198, new_n14199, new_n14200, new_n14201, new_n14202, new_n14203, new_n14204, new_n14205, new_n14206, new_n14207, new_n14208, new_n14209, new_n14210, new_n14211, new_n14212, new_n14213, new_n14214, new_n14215, new_n14216, new_n14217, new_n14218, new_n14219, new_n14220, new_n14221, new_n14222, new_n14223, new_n14224, new_n14225, new_n14226, new_n14227, new_n14228, new_n14229, new_n14230, new_n14231, new_n14232, new_n14233, new_n14234, new_n14235, new_n14236, new_n14237, new_n14238, new_n14239, new_n14240, new_n14241, new_n14242, new_n14243, new_n14244, new_n14245, new_n14246, new_n14247, new_n14248, new_n14249, new_n14250, new_n14251, new_n14252, new_n14253, new_n14254, new_n14255, new_n14256, new_n14257, new_n14258, new_n14259, new_n14260, new_n14261, new_n14262, new_n14263, new_n14264, new_n14265, new_n14266, new_n14267, new_n14268, new_n14269, new_n14270, new_n14271, new_n14272, new_n14273, new_n14274, new_n14275, new_n14276, new_n14277, new_n14278, new_n14279, new_n14280, new_n14281, new_n14282, new_n14283, new_n14284, new_n14285, new_n14286, new_n14287, new_n14288, new_n14289, new_n14290, new_n14291, new_n14292, new_n14293, new_n14294, new_n14295, new_n14296, new_n14297, new_n14298, new_n14299, new_n14300, new_n14301, new_n14302, new_n14303, new_n14304, new_n14305, new_n14306, new_n14307, new_n14308, new_n14309, new_n14310, new_n14311, new_n14312, new_n14313, new_n14314, new_n14315, new_n14316, new_n14317, new_n14318, new_n14319, new_n14320, new_n14321, new_n14322, new_n14323, new_n14324, new_n14325, new_n14326, new_n14327, new_n14328, new_n14329, new_n14330, new_n14331, new_n14332, new_n14333, new_n14334, new_n14335, new_n14336, new_n14337, new_n14338, new_n14339, new_n14340, new_n14341, new_n14342, new_n14343, new_n14344, new_n14345, new_n14346, new_n14347, new_n14348, new_n14349, new_n14350, new_n14351, new_n14352, new_n14353, new_n14354, new_n14355, new_n14356, new_n14357, new_n14358, new_n14359, new_n14360, new_n14361, new_n14362, new_n14363, new_n14364, new_n14365, new_n14366, new_n14367, new_n14368, new_n14369, new_n14370, new_n14371, new_n14372, new_n14373, new_n14374, new_n14375, new_n14376, new_n14377, new_n14378, new_n14379, new_n14380, new_n14381, new_n14382, new_n14383, new_n14384, new_n14385, new_n14386, new_n14387, new_n14388, new_n14389, new_n14390, new_n14391, new_n14392, new_n14393, new_n14394, new_n14395, new_n14396, new_n14397, new_n14398, new_n14399, new_n14400, new_n14401, new_n14402, new_n14403, new_n14404, new_n14405, new_n14406, new_n14407, new_n14408, new_n14409, new_n14410, new_n14411, new_n14412, new_n14413, new_n14414, new_n14415, new_n14416, new_n14417, new_n14418, new_n14419, new_n14420, new_n14421, new_n14422, new_n14423, new_n14424, new_n14425, new_n14426, new_n14427, new_n14428, new_n14429, new_n14430, new_n14431, new_n14432, new_n14433, new_n14434, new_n14435, new_n14436, new_n14437, new_n14438, new_n14439, new_n14440, new_n14441, new_n14442, new_n14443, new_n14444, new_n14445, new_n14446, new_n14447, new_n14448, new_n14449, new_n14450, new_n14451, new_n14452, new_n14453, new_n14454, new_n14455, new_n14456, new_n14457, new_n14458, new_n14459, new_n14460, new_n14461, new_n14462, new_n14463, new_n14464, new_n14465, new_n14466, new_n14467, new_n14468, new_n14469, new_n14470, new_n14471, new_n14472, new_n14473, new_n14474, new_n14475, new_n14476, new_n14477, new_n14478, new_n14479, new_n14480, new_n14481, new_n14482, new_n14483, new_n14484, new_n14485, new_n14486, new_n14487, new_n14488, new_n14489, new_n14490, new_n14491, new_n14492, new_n14493, new_n14494, new_n14495, new_n14496, new_n14497, new_n14498, new_n14499, new_n14500, new_n14501, new_n14502, new_n14503, new_n14504, new_n14505, new_n14506, new_n14507, new_n14508, new_n14509, new_n14510, new_n14511, new_n14512, new_n14513, new_n14514, new_n14515, new_n14516, new_n14517, new_n14518, new_n14519, new_n14520, new_n14521, new_n14522, new_n14523, new_n14524, new_n14525, new_n14526, new_n14527, new_n14528, new_n14529, new_n14530, new_n14531, new_n14532, new_n14533, new_n14534, new_n14535, new_n14536, new_n14537, new_n14538, new_n14539, new_n14540, new_n14541, new_n14542, new_n14543, new_n14544, new_n14545, new_n14546, new_n14547, new_n14548, new_n14549, new_n14550, new_n14551, new_n14552, new_n14553, new_n14554, new_n14555, new_n14556, new_n14557, new_n14558, new_n14559, new_n14560, new_n14561, new_n14562, new_n14563, new_n14564, new_n14565, new_n14566, new_n14567, new_n14568, new_n14569, new_n14570, new_n14571, new_n14572, new_n14573, new_n14574, new_n14575, new_n14576, new_n14577, new_n14578, new_n14579, new_n14580, new_n14581, new_n14582, new_n14583, new_n14584, new_n14585, new_n14586, new_n14587, new_n14588, new_n14589, new_n14590, new_n14591, new_n14592, new_n14593, new_n14594, new_n14595, new_n14596, new_n14597, new_n14598, new_n14599, new_n14600, new_n14601, new_n14602, new_n14603, new_n14604, new_n14605, new_n14606, new_n14607, new_n14608, new_n14609, new_n14610, new_n14611, new_n14612, new_n14613, new_n14614, new_n14615, new_n14616, new_n14617, new_n14618, new_n14619, new_n14620, new_n14621, new_n14622, new_n14623, new_n14624, new_n14625, new_n14626, new_n14627, new_n14628, new_n14629, new_n14630, new_n14631, new_n14632, new_n14633, new_n14634, new_n14635, new_n14636, new_n14637, new_n14638, new_n14639, new_n14640, new_n14641, new_n14642, new_n14643, new_n14644, new_n14645, new_n14646, new_n14647, new_n14648, new_n14649, new_n14650, new_n14651, new_n14652, new_n14653, new_n14654, new_n14655, new_n14656, new_n14657, new_n14658, new_n14659, new_n14660, new_n14661, new_n14662, new_n14663, new_n14664, new_n14665, new_n14666, new_n14667, new_n14668, new_n14669, new_n14670, new_n14671, new_n14672, new_n14673, new_n14674, new_n14675, new_n14676, new_n14677, new_n14678, new_n14679, new_n14680, new_n14681, new_n14682, new_n14683, new_n14684, new_n14685, new_n14686, new_n14687, new_n14688, new_n14689, new_n14690, new_n14691, new_n14692, new_n14693, new_n14694, new_n14695, new_n14696, new_n14697, new_n14698, new_n14699, new_n14700, new_n14701, new_n14702, new_n14703, new_n14704, new_n14705, new_n14706, new_n14707, new_n14708, new_n14709, new_n14710, new_n14711, new_n14712, new_n14713, new_n14714, new_n14715, new_n14716, new_n14717, new_n14718, new_n14719, new_n14720, new_n14721, new_n14722, new_n14723, new_n14724, new_n14725, new_n14726, new_n14727, new_n14728, new_n14729, new_n14730, new_n14731, new_n14732, new_n14733, new_n14734, new_n14735, new_n14736, new_n14737, new_n14738, new_n14739, new_n14740, new_n14741, new_n14742, new_n14743, new_n14744, new_n14745, new_n14746, new_n14747, new_n14748, new_n14749, new_n14750, new_n14751, new_n14752, new_n14753, new_n14754, new_n14755, new_n14756, new_n14757, new_n14758, new_n14759, new_n14760, new_n14761, new_n14762, new_n14763, new_n14764, new_n14765, new_n14766, new_n14767, new_n14768, new_n14769, new_n14770, new_n14771, new_n14772, new_n14773, new_n14774, new_n14775, new_n14776, new_n14777, new_n14778, new_n14779, new_n14780, new_n14781, new_n14782, new_n14783, new_n14784, new_n14785, new_n14786, new_n14787, new_n14788, new_n14789, new_n14790, new_n14791, new_n14792, new_n14793, new_n14794, new_n14795, new_n14796, new_n14797, new_n14798, new_n14799, new_n14800, new_n14801, new_n14802, new_n14803, new_n14804, new_n14805, new_n14806, new_n14807, new_n14808, new_n14809, new_n14810, new_n14811, new_n14812, new_n14813, new_n14814, new_n14815, new_n14816, new_n14817, new_n14818, new_n14819, new_n14820, new_n14821, new_n14822, new_n14823, new_n14824, new_n14825, new_n14826, new_n14827, new_n14828, new_n14829, new_n14830, new_n14831, new_n14832, new_n14833, new_n14834, new_n14835, new_n14836, new_n14837, new_n14838, new_n14839, new_n14840, new_n14841, new_n14842, new_n14843, new_n14844, new_n14845, new_n14846, new_n14847, new_n14848, new_n14849, new_n14850, new_n14851, new_n14852, new_n14853, new_n14854, new_n14855, new_n14856, new_n14857, new_n14858, new_n14859, new_n14860, new_n14861, new_n14862, new_n14863, new_n14864, new_n14865, new_n14866, new_n14867, new_n14868, new_n14869, new_n14870, new_n14871, new_n14872, new_n14873, new_n14874, new_n14875, new_n14876, new_n14877, new_n14878, new_n14879, new_n14880, new_n14881, new_n14882, new_n14883, new_n14884, new_n14885, new_n14886, new_n14887, new_n14888, new_n14889, new_n14890, new_n14891, new_n14892, new_n14893, new_n14894, new_n14895, new_n14896, new_n14897, new_n14898, new_n14899, new_n14900, new_n14901, new_n14902, new_n14903, new_n14904, new_n14905, new_n14906, new_n14907, new_n14908, new_n14909, new_n14910, new_n14911, new_n14912, new_n14913, new_n14914, new_n14915, new_n14916, new_n14917, new_n14918, new_n14919, new_n14920, new_n14921, new_n14922, new_n14923, new_n14924, new_n14925, new_n14926, new_n14927, new_n14928, new_n14929, new_n14930, new_n14931, new_n14932, new_n14933, new_n14934, new_n14935, new_n14936, new_n14937, new_n14938, new_n14939, new_n14940, new_n14941, new_n14942, new_n14943, new_n14944, new_n14945, new_n14946, new_n14947, new_n14948, new_n14949, new_n14950, new_n14951, new_n14952, new_n14953, new_n14954, new_n14955, new_n14956, new_n14957, new_n14958, new_n14959, new_n14960, new_n14961, new_n14962, new_n14963, new_n14964, new_n14965, new_n14966, new_n14967, new_n14968, new_n14969, new_n14970, new_n14971, new_n14972, new_n14973, new_n14974, new_n14975, new_n14976, new_n14977, new_n14978, new_n14979, new_n14980, new_n14981, new_n14982, new_n14983, new_n14984, new_n14985, new_n14986, new_n14987, new_n14988, new_n14989, new_n14990, new_n14991, new_n14992, new_n14993, new_n14994, new_n14995, new_n14996, new_n14997, new_n14998, new_n14999, new_n15000, new_n15001, new_n15002, new_n15003, new_n15004, new_n15005, new_n15006, new_n15007, new_n15008, new_n15009, new_n15010, new_n15011, new_n15012, new_n15013, new_n15014, new_n15015, new_n15016, new_n15017, new_n15018, new_n15019, new_n15020, new_n15021, new_n15022, new_n15023, new_n15024, new_n15025, new_n15026, new_n15027, new_n15028, new_n15029, new_n15030, new_n15031, new_n15032, new_n15033, new_n15034, new_n15035, new_n15036, new_n15037, new_n15038, new_n15039, new_n15040, new_n15041, new_n15042, new_n15043, new_n15044, new_n15045, new_n15046, new_n15047, new_n15048, new_n15049, new_n15050, new_n15051, new_n15052, new_n15053, new_n15054, new_n15055, new_n15056, new_n15057, new_n15058, new_n15059, new_n15060, new_n15061, new_n15062, new_n15063, new_n15064, new_n15065, new_n15066, new_n15067, new_n15068, new_n15069, new_n15070, new_n15071, new_n15072, new_n15073, new_n15074, new_n15075, new_n15076, new_n15077, new_n15078, new_n15079, new_n15080, new_n15081, new_n15082, new_n15083, new_n15084, new_n15085, new_n15086, new_n15087, new_n15088, new_n15089, new_n15090, new_n15091, new_n15092, new_n15093, new_n15094, new_n15095, new_n15096, new_n15097, new_n15098, new_n15099, new_n15100, new_n15101, new_n15102, new_n15103, new_n15104, new_n15105, new_n15106, new_n15107, new_n15108, new_n15109, new_n15110, new_n15111, new_n15112, new_n15113, new_n15114, new_n15115, new_n15116, new_n15117, new_n15118, new_n15119, new_n15120, new_n15121, new_n15122, new_n15123, new_n15124, new_n15125, new_n15126, new_n15127, new_n15128, new_n15129, new_n15130, new_n15131, new_n15132, new_n15133, new_n15134, new_n15135, new_n15136, new_n15137, new_n15138, new_n15139, new_n15140, new_n15141, new_n15142, new_n15143, new_n15144, new_n15145, new_n15146, new_n15147, new_n15148, new_n15149, new_n15150, new_n15151, new_n15152, new_n15153, new_n15154, new_n15155, new_n15156, new_n15157, new_n15158, new_n15159, new_n15160, new_n15161, new_n15162, new_n15163, new_n15164, new_n15165, new_n15166, new_n15167, new_n15168, new_n15169, new_n15170, new_n15171, new_n15172, new_n15173, new_n15174, new_n15175, new_n15176, new_n15177, new_n15178, new_n15179, new_n15180, new_n15181, new_n15182, new_n15183, new_n15184, new_n15185, new_n15186, new_n15187, new_n15188, new_n15189, new_n15190, new_n15191, new_n15192, new_n15193, new_n15194, new_n15195, new_n15196, new_n15197, new_n15198, new_n15199, new_n15200, new_n15201, new_n15202, new_n15203, new_n15204, new_n15205, new_n15206, new_n15207, new_n15208, new_n15209, new_n15210, new_n15211, new_n15212, new_n15213, new_n15214, new_n15215, new_n15216, new_n15217, new_n15218, new_n15219, new_n15220, new_n15221, new_n15222, new_n15223, new_n15224, new_n15225, new_n15226, new_n15227, new_n15228, new_n15229, new_n15230, new_n15231, new_n15232, new_n15233, new_n15234, new_n15235, new_n15236, new_n15237, new_n15238, new_n15239, new_n15240, new_n15241, new_n15242, new_n15243, new_n15244, new_n15245, new_n15246, new_n15247, new_n15248, new_n15249, new_n15250, new_n15251, new_n15252, new_n15253, new_n15254, new_n15255, new_n15256, new_n15257, new_n15258, new_n15259, new_n15260, new_n15261, new_n15262, new_n15263, new_n15264, new_n15265, new_n15266, new_n15267, new_n15268, new_n15269, new_n15270, new_n15271, new_n15272, new_n15273, new_n15274, new_n15275, new_n15276, new_n15277, new_n15278, new_n15279, new_n15280, new_n15281, new_n15282, new_n15283, new_n15284, new_n15285, new_n15286, new_n15287, new_n15288, new_n15289, new_n15290, new_n15291, new_n15292, new_n15293, new_n15294, new_n15295, new_n15296, new_n15297, new_n15298, new_n15299, new_n15300, new_n15301, new_n15302, new_n15303, new_n15304, new_n15305, new_n15306, new_n15307, new_n15308, new_n15309, new_n15310, new_n15311, new_n15312, new_n15313, new_n15314, new_n15315, new_n15316, new_n15317, new_n15318, new_n15319, new_n15320, new_n15321, new_n15322, new_n15323, new_n15324, new_n15325, new_n15326, new_n15327, new_n15328, new_n15329, new_n15330, new_n15331, new_n15332, new_n15333, new_n15334, new_n15335, new_n15336, new_n15337, new_n15338, new_n15339, new_n15340, new_n15341, new_n15342, new_n15343, new_n15344, new_n15345, new_n15346, new_n15347, new_n15348, new_n15349, new_n15350, new_n15351, new_n15352, new_n15353, new_n15354, new_n15355, new_n15356, new_n15357, new_n15358, new_n15359, new_n15360, new_n15361, new_n15362, new_n15363, new_n15364, new_n15365, new_n15366, new_n15367, new_n15368, new_n15369, new_n15370, new_n15371, new_n15372, new_n15373, new_n15374, new_n15375, new_n15376, new_n15377, new_n15378, new_n15379, new_n15380, new_n15381, new_n15382, new_n15383, new_n15384, new_n15385, new_n15386, new_n15387, new_n15388, new_n15389, new_n15390, new_n15391, new_n15392, new_n15393, new_n15394, new_n15395, new_n15396, new_n15397, new_n15398, new_n15399, new_n15400, new_n15401, new_n15402, new_n15403, new_n15404, new_n15405, new_n15406, new_n15407, new_n15408, new_n15409, new_n15410, new_n15411, new_n15412, new_n15413, new_n15414, new_n15415, new_n15416, new_n15417, new_n15418, new_n15419, new_n15420, new_n15421, new_n15422, new_n15423, new_n15424, new_n15425, new_n15426, new_n15427, new_n15428, new_n15429, new_n15430, new_n15431, new_n15432, new_n15433, new_n15434, new_n15435, new_n15436, new_n15437, new_n15438, new_n15439, new_n15440, new_n15441, new_n15442, new_n15443, new_n15444, new_n15445, new_n15446, new_n15447, new_n15448, new_n15449, new_n15450, new_n15451, new_n15452, new_n15453, new_n15454, new_n15455, new_n15456, new_n15457, new_n15458, new_n15459, new_n15460, new_n15461, new_n15462, new_n15463, new_n15464, new_n15465, new_n15466, new_n15467, new_n15468, new_n15469, new_n15470, new_n15471, new_n15472, new_n15473, new_n15474, new_n15475, new_n15476, new_n15477, new_n15478, new_n15479, new_n15480, new_n15481, new_n15482, new_n15483, new_n15484, new_n15485, new_n15486, new_n15487, new_n15488, new_n15489, new_n15490, new_n15491, new_n15492, new_n15493, new_n15494, new_n15495, new_n15496, new_n15497, new_n15498, new_n15499, new_n15500, new_n15501, new_n15502, new_n15503, new_n15504, new_n15505, new_n15506, new_n15507, new_n15508, new_n15509, new_n15510, new_n15511, new_n15512, new_n15513, new_n15514, new_n15515, new_n15516, new_n15517, new_n15518, new_n15519, new_n15520, new_n15521, new_n15522, new_n15523, new_n15524, new_n15525, new_n15526, new_n15527, new_n15528, new_n15529, new_n15530, new_n15531, new_n15532, new_n15533, new_n15534, new_n15535, new_n15536, new_n15537, new_n15538, new_n15539, new_n15540, new_n15541, new_n15542, new_n15543, new_n15544, new_n15545, new_n15546, new_n15547, new_n15548, new_n15549, new_n15550, new_n15551, new_n15552, new_n15553, new_n15554, new_n15555, new_n15556, new_n15557, new_n15558, new_n15559, new_n15560, new_n15561, new_n15562, new_n15563, new_n15564, new_n15565, new_n15566, new_n15567, new_n15568, new_n15569, new_n15570, new_n15571, new_n15572, new_n15573, new_n15574, new_n15575, new_n15576, new_n15577, new_n15578, new_n15579, new_n15580, new_n15581, new_n15582, new_n15583, new_n15584, new_n15585, new_n15586, new_n15587, new_n15588, new_n15589, new_n15590, new_n15591, new_n15592, new_n15593, new_n15594, new_n15595, new_n15596, new_n15597, new_n15598, new_n15599, new_n15600, new_n15601, new_n15602, new_n15603, new_n15604, new_n15605, new_n15606, new_n15607, new_n15608, new_n15609, new_n15610, new_n15611, new_n15612, new_n15613, new_n15614, new_n15615, new_n15616, new_n15617, new_n15618, new_n15619, new_n15620, new_n15621, new_n15622, new_n15623, new_n15624, new_n15625, new_n15626, new_n15627, new_n15628, new_n15629, new_n15630, new_n15631, new_n15632, new_n15633, new_n15634, new_n15635, new_n15636, new_n15637, new_n15638, new_n15639, new_n15640, new_n15641, new_n15642, new_n15643, new_n15644, new_n15645, new_n15646, new_n15647, new_n15648, new_n15649, new_n15650, new_n15651, new_n15652, new_n15653, new_n15654, new_n15655, new_n15656, new_n15657, new_n15658, new_n15659, new_n15660, new_n15661, new_n15662, new_n15663, new_n15664, new_n15665, new_n15666, new_n15667, new_n15668, new_n15669, new_n15670, new_n15671, new_n15672, new_n15673, new_n15674, new_n15675, new_n15676, new_n15677, new_n15678, new_n15679, new_n15680, new_n15681, new_n15682, new_n15683, new_n15684, new_n15685, new_n15686, new_n15687, new_n15688, new_n15689, new_n15690, new_n15691, new_n15692, new_n15693, new_n15694, new_n15695, new_n15696, new_n15697, new_n15698, new_n15699, new_n15700, new_n15701, new_n15702, new_n15703, new_n15704, new_n15705, new_n15706, new_n15707, new_n15708, new_n15709, new_n15710, new_n15711, new_n15712, new_n15713, new_n15714, new_n15715, new_n15716, new_n15717, new_n15718, new_n15719, new_n15720, new_n15721, new_n15722, new_n15723, new_n15724, new_n15725, new_n15726, new_n15727, new_n15728, new_n15729, new_n15730, new_n15731, new_n15732, new_n15733, new_n15734, new_n15735, new_n15736, new_n15737, new_n15738, new_n15739, new_n15740, new_n15741, new_n15742, new_n15743, new_n15744, new_n15745, new_n15746, new_n15747, new_n15748, new_n15749, new_n15750, new_n15751, new_n15752, new_n15753, new_n15754, new_n15755, new_n15756, new_n15757, new_n15758, new_n15759, new_n15760, new_n15761, new_n15762, new_n15763, new_n15764, new_n15765, new_n15766, new_n15767, new_n15768, new_n15769, new_n15770, new_n15771, new_n15772, new_n15773, new_n15774, new_n15775, new_n15776, new_n15777, new_n15778, new_n15779, new_n15780, new_n15781, new_n15782, new_n15783, new_n15784, new_n15785, new_n15786, new_n15787, new_n15788, new_n15789, new_n15790, new_n15791, new_n15792, new_n15793, new_n15794, new_n15795, new_n15796, new_n15797, new_n15798, new_n15799, new_n15800, new_n15801, new_n15802, new_n15803, new_n15804, new_n15805, new_n15806, new_n15807, new_n15808, new_n15809, new_n15810, new_n15811, new_n15812, new_n15813, new_n15814, new_n15815, new_n15816, new_n15817, new_n15818, new_n15819, new_n15820, new_n15821, new_n15822, new_n15823, new_n15824, new_n15825, new_n15826, new_n15827, new_n15828, new_n15829, new_n15830, new_n15831, new_n15832, new_n15833, new_n15834, new_n15835, new_n15836, new_n15837, new_n15838, new_n15839, new_n15840, new_n15841, new_n15842, new_n15843, new_n15844, new_n15845, new_n15846, new_n15847, new_n15848, new_n15849, new_n15850, new_n15851, new_n15852, new_n15853, new_n15854, new_n15855, new_n15856, new_n15857, new_n15858, new_n15859, new_n15860, new_n15861, new_n15862, new_n15863, new_n15864, new_n15865, new_n15866, new_n15867, new_n15868, new_n15869, new_n15870, new_n15871, new_n15872, new_n15873, new_n15874, new_n15875, new_n15876, new_n15877, new_n15878, new_n15879, new_n15880, new_n15881, new_n15882, new_n15883, new_n15884, new_n15885, new_n15886, new_n15887, new_n15888, new_n15889, new_n15890, new_n15891, new_n15892, new_n15893, new_n15894, new_n15895, new_n15896, new_n15897, new_n15898, new_n15899, new_n15900, new_n15901, new_n15902, new_n15903, new_n15904, new_n15905, new_n15906, new_n15907, new_n15908, new_n15909, new_n15910, new_n15911, new_n15912, new_n15913, new_n15914, new_n15915, new_n15916, new_n15917, new_n15918, new_n15919, new_n15920, new_n15921, new_n15922, new_n15923, new_n15924, new_n15925, new_n15926, new_n15927, new_n15928, new_n15929, new_n15930, new_n15931, new_n15932, new_n15933, new_n15934, new_n15935, new_n15936, new_n15937, new_n15938, new_n15939, new_n15940, new_n15941, new_n15942, new_n15943, new_n15944, new_n15945, new_n15946, new_n15947, new_n15948, new_n15949, new_n15950, new_n15951, new_n15952, new_n15953, new_n15954, new_n15955, new_n15956, new_n15957, new_n15958, new_n15959, new_n15960, new_n15961, new_n15962, new_n15963, new_n15964, new_n15965, new_n15966, new_n15967, new_n15968, new_n15969, new_n15970, new_n15971, new_n15972, new_n15973, new_n15974, new_n15975, new_n15976, new_n15977, new_n15978, new_n15979, new_n15980, new_n15981, new_n15982, new_n15983, new_n15984, new_n15985, new_n15986, new_n15987, new_n15988, new_n15989, new_n15990, new_n15991, new_n15992, new_n15993, new_n15994, new_n15995, new_n15996, new_n15997, new_n15998, new_n15999, new_n16000, new_n16001, new_n16002, new_n16003, new_n16004, new_n16005, new_n16006, new_n16007, new_n16008, new_n16009, new_n16010, new_n16011, new_n16012, new_n16013, new_n16014, new_n16015, new_n16016, new_n16017, new_n16018, new_n16019, new_n16020, new_n16021, new_n16022, new_n16023, new_n16024, new_n16025, new_n16026, new_n16027, new_n16028, new_n16029, new_n16030, new_n16031, new_n16032, new_n16033, new_n16034, new_n16035, new_n16036, new_n16037, new_n16038, new_n16039, new_n16040, new_n16041, new_n16042, new_n16043, new_n16044, new_n16045, new_n16046, new_n16047, new_n16048, new_n16049, new_n16050, new_n16051, new_n16052, new_n16053, new_n16054, new_n16055, new_n16056, new_n16057, new_n16058, new_n16059, new_n16060, new_n16061, new_n16062, new_n16063, new_n16064, new_n16065, new_n16066, new_n16067, new_n16068, new_n16069, new_n16070, new_n16071, new_n16072, new_n16073, new_n16074, new_n16075, new_n16076, new_n16077, new_n16078, new_n16079, new_n16080, new_n16081, new_n16082, new_n16083, new_n16084, new_n16085, new_n16086, new_n16087, new_n16088, new_n16089, new_n16090, new_n16091, new_n16092, new_n16093, new_n16094, new_n16095, new_n16096, new_n16097, new_n16098, new_n16099, new_n16100, new_n16101, new_n16102, new_n16103, new_n16104, new_n16105, new_n16106, new_n16107, new_n16108, new_n16109, new_n16110, new_n16111, new_n16112, new_n16113, new_n16114, new_n16115, new_n16116, new_n16117, new_n16118, new_n16119, new_n16120, new_n16121, new_n16122, new_n16123, new_n16124, new_n16125, new_n16126, new_n16127, new_n16128, new_n16129, new_n16130, new_n16131, new_n16132, new_n16133, new_n16134, new_n16135, new_n16136, new_n16137, new_n16138, new_n16139, new_n16140, new_n16141, new_n16142, new_n16143, new_n16144, new_n16145, new_n16146, new_n16147, new_n16148, new_n16149, new_n16150, new_n16151, new_n16152, new_n16153, new_n16154, new_n16155, new_n16156, new_n16157, new_n16158, new_n16159, new_n16160, new_n16161, new_n16162, new_n16163, new_n16164, new_n16165, new_n16166, new_n16167, new_n16168, new_n16169, new_n16170, new_n16171, new_n16172, new_n16173, new_n16174, new_n16175, new_n16176, new_n16177, new_n16178, new_n16179, new_n16180, new_n16181, new_n16182, new_n16183, new_n16184, new_n16185, new_n16186, new_n16187, new_n16188, new_n16189, new_n16190, new_n16191, new_n16192, new_n16193, new_n16194, new_n16195, new_n16196, new_n16197, new_n16198, new_n16199, new_n16200, new_n16201, new_n16202, new_n16203, new_n16204, new_n16205, new_n16206, new_n16207, new_n16208, new_n16209, new_n16210, new_n16211, new_n16212, new_n16213, new_n16214, new_n16215, new_n16216, new_n16217, new_n16218, new_n16219, new_n16220, new_n16221, new_n16222, new_n16223, new_n16224, new_n16225, new_n16226, new_n16227, new_n16228, new_n16229, new_n16230, new_n16231, new_n16232, new_n16233, new_n16234, new_n16235, new_n16236, new_n16237, new_n16238, new_n16239, new_n16240, new_n16241, new_n16242, new_n16243, new_n16244, new_n16245, new_n16246, new_n16247, new_n16248, new_n16249, new_n16250, new_n16251, new_n16252, new_n16253, new_n16254, new_n16255, new_n16256, new_n16257, new_n16258, new_n16259, new_n16260, new_n16261, new_n16262, new_n16263, new_n16264, new_n16265, new_n16266, new_n16267, new_n16268, new_n16269, new_n16270, new_n16271, new_n16272, new_n16273, new_n16274, new_n16275, new_n16276, new_n16277, new_n16278, new_n16279, new_n16280, new_n16281, new_n16282, new_n16283, new_n16284, new_n16285, new_n16286, new_n16287, new_n16288, new_n16289, new_n16290, new_n16291, new_n16292, new_n16293, new_n16294, new_n16295, new_n16296, new_n16297, new_n16298, new_n16299, new_n16300, new_n16301, new_n16302, new_n16303, new_n16304, new_n16305, new_n16306, new_n16307, new_n16308, new_n16309, new_n16310, new_n16311, new_n16312, new_n16313, new_n16314, new_n16315, new_n16316, new_n16317, new_n16318, new_n16319, new_n16320, new_n16321, new_n16322, new_n16323, new_n16324, new_n16325, new_n16326, new_n16327, new_n16328, new_n16329, new_n16330, new_n16331, new_n16332, new_n16333, new_n16334, new_n16335, new_n16336, new_n16337, new_n16338, new_n16339, new_n16340, new_n16341, new_n16342, new_n16343, new_n16344, new_n16345, new_n16346, new_n16347, new_n16348, new_n16349, new_n16350, new_n16351, new_n16352, new_n16353, new_n16354, new_n16355, new_n16356, new_n16357, new_n16358, new_n16359, new_n16360, new_n16361, new_n16362, new_n16363, new_n16364, new_n16365, new_n16366, new_n16367, new_n16368, new_n16369, new_n16370, new_n16371, new_n16372, new_n16373, new_n16374, new_n16375, new_n16376, new_n16377, new_n16378, new_n16379, new_n16380, new_n16381, new_n16382, new_n16383, new_n16384, new_n16385, new_n16386, new_n16387, new_n16388, new_n16389, new_n16390, new_n16391, new_n16392, new_n16393, new_n16394, new_n16395, new_n16396, new_n16397, new_n16398, new_n16399, new_n16400, new_n16401, new_n16402, new_n16403, new_n16404, new_n16405, new_n16406, new_n16407, new_n16408, new_n16409, new_n16410, new_n16411, new_n16412, new_n16413, new_n16414, new_n16415, new_n16416, new_n16417, new_n16418, new_n16419, new_n16420, new_n16421, new_n16422, new_n16423, new_n16424, new_n16425, new_n16426, new_n16427, new_n16428, new_n16429, new_n16430, new_n16431, new_n16432, new_n16433, new_n16434, new_n16435, new_n16436, new_n16437, new_n16438, new_n16439, new_n16440, new_n16441, new_n16442, new_n16443, new_n16444, new_n16445, new_n16446, new_n16447, new_n16448, new_n16449, new_n16450, new_n16451, new_n16452, new_n16453, new_n16454, new_n16455, new_n16456, new_n16457, new_n16458, new_n16459, new_n16460, new_n16461, new_n16462, new_n16463, new_n16464, new_n16465, new_n16466, new_n16467, new_n16468, new_n16469, new_n16470, new_n16471, new_n16472, new_n16473, new_n16474, new_n16475, new_n16476, new_n16477, new_n16478, new_n16479, new_n16480, new_n16481, new_n16482, new_n16483, new_n16484, new_n16485, new_n16486, new_n16487, new_n16488, new_n16489, new_n16490, new_n16491, new_n16492, new_n16493, new_n16494, new_n16495, new_n16496, new_n16497, new_n16498, new_n16499, new_n16500, new_n16501, new_n16502, new_n16503, new_n16504, new_n16505, new_n16506, new_n16507, new_n16508, new_n16509, new_n16510, new_n16511, new_n16512, new_n16513, new_n16514, new_n16515, new_n16516, new_n16517, new_n16518, new_n16519, new_n16520, new_n16521, new_n16522, new_n16523, new_n16524, new_n16525, new_n16526, new_n16527, new_n16528, new_n16529, new_n16530, new_n16531, new_n16532, new_n16533, new_n16534, new_n16535, new_n16536, new_n16537, new_n16538, new_n16539, new_n16540, new_n16541, new_n16542, new_n16543, new_n16544, new_n16545, new_n16546, new_n16547, new_n16548, new_n16549, new_n16550, new_n16551, new_n16552, new_n16553, new_n16554, new_n16555, new_n16556, new_n16557, new_n16558, new_n16559, new_n16560, new_n16561, new_n16562, new_n16563, new_n16564, new_n16565, new_n16566, new_n16567, new_n16568, new_n16569, new_n16570, new_n16571, new_n16572, new_n16573, new_n16574, new_n16575, new_n16576, new_n16577, new_n16578, new_n16579, new_n16580, new_n16581, new_n16582, new_n16583, new_n16584, new_n16585, new_n16586, new_n16587, new_n16588, new_n16589, new_n16590, new_n16591, new_n16592, new_n16593, new_n16594, new_n16595, new_n16596, new_n16597, new_n16598, new_n16599, new_n16600, new_n16601, new_n16602, new_n16603, new_n16604, new_n16605, new_n16606, new_n16607, new_n16608, new_n16609, new_n16610, new_n16611, new_n16612, new_n16613, new_n16614, new_n16615, new_n16616, new_n16617, new_n16618, new_n16619, new_n16620, new_n16621, new_n16622, new_n16623, new_n16624, new_n16625, new_n16626, new_n16627, new_n16628, new_n16629, new_n16630, new_n16631, new_n16632, new_n16633, new_n16634, new_n16635, new_n16636, new_n16637, new_n16638, new_n16639, new_n16640, new_n16641, new_n16642, new_n16643, new_n16644, new_n16645, new_n16646, new_n16647, new_n16648, new_n16649, new_n16650, new_n16651, new_n16652, new_n16653, new_n16654, new_n16655, new_n16656, new_n16657, new_n16658, new_n16659, new_n16660, new_n16661, new_n16662, new_n16663, new_n16664, new_n16665, new_n16666, new_n16667, new_n16668, new_n16669, new_n16670, new_n16671, new_n16672, new_n16673, new_n16674, new_n16675, new_n16676, new_n16677, new_n16678, new_n16679, new_n16680, new_n16681, new_n16682, new_n16683, new_n16684, new_n16685, new_n16686, new_n16687, new_n16688, new_n16689, new_n16690, new_n16691, new_n16692, new_n16693, new_n16694, new_n16695, new_n16696, new_n16697, new_n16698, new_n16699, new_n16700, new_n16701, new_n16702, new_n16703, new_n16704, new_n16705, new_n16706, new_n16707, new_n16708, new_n16709, new_n16710, new_n16711, new_n16712, new_n16713, new_n16714, new_n16715, new_n16716, new_n16717, new_n16718, new_n16719, new_n16720, new_n16721, new_n16722, new_n16723, new_n16724, new_n16725, new_n16726, new_n16727, new_n16728, new_n16729, new_n16730, new_n16731, new_n16732, new_n16733, new_n16734, new_n16735, new_n16736, new_n16737, new_n16738, new_n16739, new_n16740, new_n16741, new_n16742, new_n16743, new_n16744, new_n16745, new_n16746, new_n16747, new_n16748, new_n16749, new_n16750, new_n16751, new_n16752, new_n16753, new_n16754, new_n16755, new_n16756, new_n16757, new_n16758, new_n16759, new_n16760, new_n16761, new_n16762, new_n16763, new_n16764, new_n16765, new_n16766, new_n16767, new_n16768, new_n16769, new_n16770, new_n16771, new_n16772, new_n16773, new_n16774, new_n16775, new_n16776, new_n16777, new_n16778, new_n16779, new_n16780, new_n16781, new_n16782, new_n16783, new_n16784, new_n16785, new_n16786, new_n16787, new_n16788, new_n16789, new_n16790, new_n16791, new_n16792, new_n16793, new_n16794, new_n16795, new_n16796, new_n16797, new_n16798, new_n16799, new_n16800, new_n16801, new_n16802, new_n16803, new_n16804, new_n16805, new_n16806, new_n16807, new_n16808, new_n16809, new_n16810, new_n16811, new_n16812, new_n16813, new_n16814, new_n16815, new_n16816, new_n16817, new_n16818, new_n16819, new_n16820, new_n16821, new_n16822, new_n16823, new_n16824, new_n16825, new_n16826, new_n16827, new_n16828, new_n16829, new_n16830, new_n16831, new_n16832, new_n16833, new_n16834, new_n16835, new_n16836, new_n16837, new_n16838, new_n16839, new_n16840, new_n16841, new_n16842, new_n16843, new_n16844, new_n16845, new_n16846, new_n16847, new_n16848, new_n16849, new_n16850, new_n16851, new_n16852, new_n16853, new_n16854, new_n16855, new_n16856, new_n16857, new_n16858, new_n16859, new_n16860, new_n16861, new_n16862, new_n16863, new_n16864, new_n16865, new_n16866, new_n16867, new_n16868, new_n16869, new_n16870, new_n16871, new_n16872, new_n16873, new_n16874, new_n16875, new_n16876, new_n16877, new_n16878, new_n16879, new_n16880, new_n16881, new_n16882, new_n16883, new_n16884, new_n16885, new_n16886, new_n16887, new_n16888, new_n16889, new_n16890, new_n16891, new_n16892, new_n16893, new_n16894, new_n16895, new_n16896, new_n16897, new_n16898, new_n16899, new_n16900, new_n16901, new_n16902, new_n16903, new_n16904, new_n16905, new_n16906, new_n16907, new_n16908, new_n16909, new_n16910, new_n16911, new_n16912, new_n16913, new_n16914, new_n16915, new_n16916, new_n16917, new_n16918, new_n16919, new_n16920, new_n16921, new_n16922, new_n16923, new_n16924, new_n16925, new_n16926, new_n16927, new_n16928, new_n16929, new_n16930, new_n16931, new_n16932, new_n16933, new_n16934, new_n16935, new_n16936, new_n16937, new_n16938, new_n16939, new_n16940, new_n16941, new_n16942, new_n16943, new_n16944, new_n16945, new_n16946, new_n16947, new_n16948, new_n16949, new_n16950, new_n16951, new_n16952, new_n16953, new_n16954, new_n16955, new_n16956, new_n16957, new_n16958, new_n16959, new_n16960, new_n16961, new_n16962, new_n16963, new_n16964, new_n16965, new_n16966, new_n16967, new_n16968, new_n16969, new_n16970, new_n16971, new_n16972, new_n16973, new_n16974, new_n16975, new_n16976, new_n16977, new_n16978, new_n16979, new_n16980, new_n16981, new_n16982, new_n16983, new_n16984, new_n16985, new_n16986, new_n16987, new_n16988, new_n16989, new_n16990, new_n16991, new_n16992, new_n16993, new_n16994, new_n16995, new_n16996, new_n16997, new_n16998, new_n16999, new_n17000, new_n17001, new_n17002, new_n17003, new_n17004, new_n17005, new_n17006, new_n17007, new_n17008, new_n17009, new_n17010, new_n17011, new_n17012, new_n17013, new_n17014, new_n17015, new_n17016, new_n17017, new_n17018, new_n17019, new_n17020, new_n17021, new_n17022, new_n17023, new_n17024, new_n17025, new_n17026, new_n17027, new_n17028, new_n17029, new_n17030, new_n17031, new_n17032, new_n17033, new_n17034, new_n17035, new_n17036, new_n17037, new_n17038, new_n17039, new_n17040, new_n17041, new_n17042, new_n17043, new_n17044, new_n17045, new_n17046, new_n17047, new_n17048, new_n17049, new_n17050, new_n17051, new_n17052, new_n17053, new_n17054, new_n17055, new_n17056, new_n17057, new_n17058, new_n17059, new_n17060, new_n17061, new_n17062, new_n17063, new_n17064, new_n17065, new_n17066, new_n17067, new_n17068, new_n17069, new_n17070, new_n17071, new_n17072, new_n17073, new_n17074, new_n17075, new_n17076, new_n17077, new_n17078, new_n17079, new_n17080, new_n17081, new_n17082, new_n17083, new_n17084, new_n17085, new_n17086, new_n17087, new_n17088, new_n17089, new_n17090, new_n17091, new_n17092, new_n17093, new_n17094, new_n17095, new_n17096, new_n17097, new_n17098, new_n17099, new_n17100, new_n17101, new_n17102, new_n17103, new_n17104, new_n17105, new_n17106, new_n17107, new_n17108, new_n17109, new_n17110, new_n17111, new_n17112, new_n17113, new_n17114, new_n17115, new_n17116, new_n17117, new_n17118, new_n17119, new_n17120, new_n17121, new_n17122, new_n17123, new_n17124, new_n17125, new_n17126, new_n17127, new_n17128, new_n17129, new_n17130, new_n17131, new_n17132, new_n17133, new_n17134, new_n17135, new_n17136, new_n17137, new_n17138, new_n17139, new_n17140, new_n17141, new_n17142, new_n17143, new_n17144, new_n17145, new_n17146, new_n17147, new_n17148, new_n17149, new_n17150, new_n17151, new_n17152, new_n17153, new_n17154, new_n17155, new_n17156, new_n17157, new_n17158, new_n17159, new_n17160, new_n17161, new_n17162, new_n17163, new_n17164, new_n17165, new_n17166, new_n17167, new_n17168, new_n17169, new_n17170, new_n17171, new_n17172, new_n17173, new_n17174, new_n17175, new_n17176, new_n17177, new_n17178, new_n17179, new_n17180, new_n17181, new_n17182, new_n17183, new_n17184, new_n17185, new_n17186, new_n17187, new_n17188, new_n17189, new_n17190, new_n17191, new_n17192, new_n17193, new_n17194, new_n17195, new_n17196, new_n17197, new_n17198, new_n17199, new_n17200, new_n17201, new_n17202, new_n17203, new_n17204, new_n17205, new_n17206, new_n17207, new_n17208, new_n17209, new_n17210, new_n17211, new_n17212, new_n17213, new_n17214, new_n17215, new_n17216, new_n17217, new_n17218, new_n17219, new_n17220, new_n17221, new_n17222, new_n17223, new_n17224, new_n17225, new_n17226, new_n17227, new_n17228, new_n17229, new_n17230, new_n17231, new_n17232, new_n17233, new_n17234, new_n17235, new_n17236, new_n17237, new_n17238, new_n17239, new_n17240, new_n17241, new_n17242, new_n17243, new_n17244, new_n17245, new_n17246, new_n17247, new_n17248, new_n17249, new_n17250, new_n17251, new_n17252, new_n17253, new_n17254, new_n17255, new_n17256, new_n17257, new_n17258, new_n17259, new_n17260, new_n17261, new_n17262, new_n17263, new_n17264, new_n17265, new_n17266, new_n17267, new_n17268, new_n17269, new_n17270, new_n17271, new_n17272, new_n17273, new_n17274, new_n17275, new_n17276, new_n17277, new_n17278, new_n17279, new_n17280, new_n17281, new_n17282, new_n17283, new_n17284, new_n17285, new_n17286, new_n17287, new_n17288, new_n17289, new_n17290, new_n17291, new_n17292, new_n17293, new_n17294, new_n17295, new_n17296, new_n17297, new_n17298, new_n17299, new_n17300, new_n17301, new_n17302, new_n17303, new_n17304, new_n17305, new_n17306, new_n17307, new_n17308, new_n17309, new_n17310, new_n17311, new_n17312, new_n17313, new_n17314, new_n17315, new_n17316, new_n17317, new_n17318, new_n17319, new_n17320, new_n17321, new_n17322, new_n17323, new_n17324, new_n17325, new_n17326, new_n17327, new_n17328, new_n17329, new_n17330, new_n17331, new_n17332, new_n17333, new_n17334, new_n17335, new_n17336, new_n17337, new_n17338, new_n17339, new_n17340, new_n17341, new_n17342, new_n17343, new_n17344, new_n17345, new_n17346, new_n17347, new_n17348, new_n17349, new_n17350, new_n17351, new_n17352, new_n17353, new_n17354, new_n17355, new_n17356, new_n17357, new_n17358, new_n17359, new_n17360, new_n17361, new_n17362, new_n17363, new_n17364, new_n17365, new_n17366, new_n17367, new_n17368, new_n17369, new_n17370, new_n17371, new_n17372, new_n17373, new_n17374, new_n17375, new_n17376, new_n17377, new_n17378, new_n17379, new_n17380, new_n17381, new_n17382, new_n17383, new_n17384, new_n17385, new_n17386, new_n17387, new_n17388, new_n17389, new_n17390, new_n17391, new_n17392, new_n17393, new_n17394, new_n17395, new_n17396, new_n17397, new_n17398, new_n17399, new_n17400, new_n17401, new_n17402, new_n17403, new_n17404, new_n17405, new_n17406, new_n17407, new_n17408, new_n17409, new_n17410, new_n17411, new_n17412, new_n17413, new_n17414, new_n17415, new_n17416, new_n17417, new_n17418, new_n17419, new_n17420, new_n17421, new_n17422, new_n17423, new_n17424, new_n17425, new_n17426, new_n17427, new_n17428, new_n17429, new_n17430, new_n17431, new_n17432, new_n17433, new_n17434, new_n17435, new_n17436, new_n17437, new_n17438, new_n17439, new_n17440, new_n17441, new_n17442, new_n17443, new_n17444, new_n17445, new_n17446, new_n17447, new_n17448, new_n17449, new_n17450, new_n17451, new_n17452, new_n17453, new_n17454, new_n17455, new_n17456, new_n17457, new_n17458, new_n17459, new_n17460, new_n17461, new_n17462, new_n17463, new_n17464, new_n17465, new_n17466, new_n17467, new_n17468, new_n17469, new_n17470, new_n17471, new_n17472, new_n17473, new_n17474, new_n17475, new_n17476, new_n17477, new_n17478, new_n17479, new_n17480, new_n17481, new_n17482, new_n17483, new_n17484, new_n17485, new_n17486, new_n17487, new_n17488, new_n17489, new_n17490, new_n17491, new_n17492, new_n17493, new_n17494, new_n17495, new_n17496, new_n17497, new_n17498, new_n17499, new_n17500, new_n17501, new_n17502, new_n17503, new_n17504, new_n17505, new_n17506, new_n17507, new_n17508, new_n17509, new_n17510, new_n17511, new_n17512, new_n17513, new_n17514, new_n17515, new_n17516, new_n17517, new_n17518, new_n17519, new_n17520, new_n17521, new_n17522, new_n17523, new_n17524, new_n17525, new_n17526, new_n17527, new_n17528, new_n17529, new_n17530, new_n17531, new_n17532, new_n17533, new_n17534, new_n17535, new_n17536, new_n17537, new_n17538, new_n17539, new_n17540, new_n17541, new_n17542, new_n17543, new_n17544, new_n17545, new_n17546, new_n17547, new_n17548, new_n17549, new_n17550, new_n17551, new_n17552, new_n17553, new_n17554, new_n17555, new_n17556, new_n17557, new_n17558, new_n17559, new_n17560, new_n17561, new_n17562, new_n17563, new_n17564, new_n17565, new_n17566, new_n17567, new_n17568, new_n17569, new_n17570, new_n17571, new_n17572, new_n17573, new_n17574, new_n17575, new_n17576, new_n17577, new_n17578, new_n17579, new_n17580, new_n17581, new_n17582, new_n17583, new_n17584, new_n17585, new_n17586, new_n17587, new_n17588, new_n17589, new_n17590, new_n17591, new_n17592, new_n17593, new_n17594, new_n17595, new_n17596, new_n17597, new_n17598, new_n17599, new_n17600, new_n17601, new_n17602, new_n17603, new_n17604, new_n17605, new_n17606, new_n17607, new_n17608, new_n17609, new_n17610, new_n17611, new_n17612, new_n17613, new_n17614, new_n17615, new_n17616, new_n17617, new_n17618, new_n17619, new_n17620, new_n17621, new_n17622, new_n17623, new_n17624, new_n17625, new_n17626, new_n17627, new_n17628, new_n17629, new_n17630, new_n17631, new_n17632, new_n17633, new_n17634, new_n17635, new_n17636, new_n17637, new_n17638, new_n17639, new_n17640, new_n17641, new_n17642, new_n17643, new_n17644, new_n17645, new_n17646, new_n17647, new_n17648, new_n17649, new_n17650, new_n17651, new_n17652, new_n17653, new_n17654, new_n17655, new_n17656, new_n17657, new_n17658, new_n17659, new_n17660, new_n17661, new_n17662, new_n17663, new_n17664, new_n17665, new_n17666, new_n17667, new_n17668, new_n17669, new_n17670, new_n17671, new_n17672, new_n17673, new_n17674, new_n17675, new_n17676, new_n17677, new_n17678, new_n17679, new_n17680, new_n17681, new_n17682, new_n17683, new_n17684, new_n17685, new_n17686, new_n17687, new_n17688, new_n17689, new_n17690, new_n17691, new_n17692, new_n17693, new_n17694, new_n17695, new_n17696, new_n17697, new_n17698, new_n17699, new_n17700, new_n17701, new_n17702, new_n17703, new_n17704, new_n17705, new_n17706, new_n17707, new_n17708, new_n17709, new_n17710, new_n17711, new_n17712, new_n17713, new_n17714, new_n17715, new_n17716, new_n17717, new_n17718, new_n17719, new_n17720, new_n17721, new_n17722, new_n17723, new_n17724, new_n17725, new_n17726, new_n17727, new_n17728, new_n17729, new_n17730, new_n17731, new_n17732, new_n17733, new_n17734, new_n17735, new_n17736, new_n17737, new_n17738, new_n17739, new_n17740, new_n17741, new_n17742, new_n17743, new_n17744, new_n17745, new_n17746, new_n17747, new_n17748, new_n17749, new_n17750, new_n17751, new_n17752, new_n17753, new_n17754, new_n17755, new_n17756, new_n17757, new_n17758, new_n17759, new_n17760, new_n17761, new_n17762, new_n17763, new_n17764, new_n17765, new_n17766, new_n17767, new_n17768, new_n17769, new_n17770, new_n17771, new_n17772, new_n17773, new_n17774, new_n17775, new_n17776, new_n17777, new_n17778, new_n17779, new_n17780, new_n17781, new_n17782, new_n17783, new_n17784, new_n17785, new_n17786, new_n17787, new_n17788, new_n17789, new_n17790, new_n17791, new_n17792, new_n17793, new_n17794, new_n17795, new_n17796, new_n17797, new_n17798, new_n17799, new_n17800, new_n17801, new_n17802, new_n17803, new_n17804, new_n17805, new_n17806, new_n17807, new_n17808, new_n17809, new_n17810, new_n17811, new_n17812, new_n17813, new_n17814, new_n17815, new_n17816, new_n17817, new_n17818, new_n17819, new_n17820, new_n17821, new_n17822, new_n17823, new_n17824, new_n17825, new_n17826, new_n17827, new_n17828, new_n17829, new_n17830, new_n17831, new_n17832, new_n17833, new_n17834, new_n17835, new_n17836, new_n17837, new_n17838, new_n17839, new_n17840, new_n17841, new_n17842, new_n17843, new_n17844, new_n17845, new_n17846, new_n17847, new_n17848, new_n17849, new_n17850, new_n17851, new_n17852, new_n17853, new_n17854, new_n17855, new_n17856, new_n17857, new_n17858, new_n17859, new_n17860, new_n17861, new_n17862, new_n17863, new_n17864, new_n17865, new_n17866, new_n17867, new_n17868, new_n17869, new_n17870, new_n17871, new_n17872, new_n17873, new_n17874, new_n17875, new_n17876, new_n17877, new_n17878, new_n17879, new_n17880, new_n17881, new_n17882, new_n17883, new_n17884, new_n17885, new_n17886, new_n17887, new_n17888, new_n17889, new_n17890, new_n17891, new_n17892, new_n17893, new_n17894, new_n17895, new_n17896, new_n17897, new_n17898, new_n17899, new_n17900, new_n17901, new_n17902, new_n17903, new_n17904, new_n17905, new_n17906, new_n17907, new_n17908, new_n17909, new_n17910, new_n17911, new_n17912, new_n17913, new_n17914, new_n17915, new_n17916, new_n17917, new_n17918, new_n17919, new_n17920, new_n17921, new_n17922, new_n17923, new_n17924, new_n17925, new_n17926, new_n17927, new_n17928, new_n17929, new_n17930, new_n17931, new_n17932, new_n17933, new_n17934, new_n17935, new_n17936, new_n17937, new_n17938, new_n17939, new_n17940, new_n17941, new_n17942, new_n17943, new_n17944, new_n17945, new_n17946, new_n17947, new_n17948, new_n17949, new_n17950, new_n17951, new_n17952, new_n17953, new_n17954, new_n17955, new_n17956, new_n17957, new_n17958, new_n17959, new_n17960, new_n17961, new_n17962, new_n17963, new_n17964, new_n17965, new_n17966, new_n17967, new_n17968, new_n17969, new_n17970, new_n17971, new_n17972, new_n17973, new_n17974, new_n17975, new_n17976, new_n17977, new_n17978, new_n17979, new_n17980, new_n17981, new_n17982, new_n17983, new_n17984, new_n17985, new_n17986, new_n17987, new_n17988, new_n17989, new_n17990, new_n17991, new_n17992, new_n17993, new_n17994, new_n17995, new_n17996, new_n17997, new_n17998, new_n17999, new_n18000, new_n18001, new_n18002, new_n18003, new_n18004, new_n18005, new_n18006, new_n18007, new_n18008, new_n18009, new_n18010, new_n18011, new_n18012, new_n18013, new_n18014, new_n18015, new_n18016, new_n18017, new_n18018, new_n18019, new_n18020, new_n18021, new_n18022, new_n18023, new_n18024, new_n18025, new_n18026, new_n18027, new_n18028, new_n18029, new_n18030, new_n18031, new_n18032, new_n18033, new_n18034, new_n18035, new_n18036, new_n18037, new_n18038, new_n18039, new_n18040, new_n18041, new_n18042, new_n18043, new_n18044, new_n18045, new_n18046, new_n18047, new_n18048, new_n18049, new_n18050, new_n18051, new_n18052, new_n18053, new_n18054, new_n18055, new_n18056, new_n18057, new_n18058, new_n18059, new_n18060, new_n18061, new_n18062, new_n18063, new_n18064, new_n18065, new_n18066, new_n18067, new_n18068, new_n18069, new_n18070, new_n18071, new_n18072, new_n18073, new_n18074, new_n18075, new_n18076, new_n18077, new_n18078, new_n18079, new_n18080, new_n18081, new_n18082, new_n18083, new_n18084, new_n18085, new_n18086, new_n18087, new_n18088, new_n18089, new_n18090, new_n18091, new_n18092, new_n18093, new_n18094, new_n18095, new_n18096, new_n18097, new_n18098, new_n18099, new_n18100, new_n18101, new_n18102, new_n18103, new_n18104, new_n18105, new_n18106, new_n18107, new_n18108, new_n18109, new_n18110, new_n18111, new_n18112, new_n18113, new_n18114, new_n18115, new_n18116, new_n18117, new_n18118, new_n18119, new_n18120, new_n18121, new_n18122, new_n18123, new_n18124, new_n18125, new_n18126, new_n18127, new_n18128, new_n18129, new_n18130, new_n18131, new_n18132, new_n18133, new_n18134, new_n18135, new_n18136, new_n18137, new_n18138, new_n18139, new_n18140, new_n18141, new_n18142, new_n18143, new_n18144, new_n18145, new_n18146, new_n18147, new_n18148, new_n18149, new_n18150, new_n18151, new_n18152, new_n18153, new_n18154, new_n18155, new_n18156, new_n18157, new_n18158, new_n18159, new_n18160, new_n18161, new_n18162, new_n18163, new_n18164, new_n18165, new_n18166, new_n18167, new_n18168, new_n18169, new_n18170, new_n18171, new_n18172, new_n18173, new_n18174, new_n18175, new_n18176, new_n18177, new_n18178, new_n18179, new_n18180, new_n18181, new_n18182, new_n18183, new_n18184, new_n18185, new_n18186, new_n18187, new_n18188, new_n18189, new_n18190, new_n18191, new_n18192, new_n18193, new_n18194, new_n18195, new_n18196, new_n18197, new_n18198, new_n18199, new_n18200, new_n18201, new_n18202, new_n18203, new_n18204, new_n18205, new_n18206, new_n18207, new_n18208, new_n18209, new_n18210, new_n18211, new_n18212, new_n18213, new_n18214, new_n18215, new_n18216, new_n18217, new_n18218, new_n18219, new_n18220, new_n18221, new_n18222, new_n18223, new_n18224, new_n18225, new_n18226, new_n18227, new_n18228, new_n18229, new_n18230, new_n18231, new_n18232, new_n18233, new_n18234, new_n18235, new_n18236, new_n18237, new_n18238, new_n18239, new_n18240, new_n18241, new_n18242, new_n18243, new_n18244, new_n18245, new_n18246, new_n18247, new_n18248, new_n18249, new_n18250, new_n18251, new_n18252, new_n18253, new_n18254, new_n18255, new_n18256, new_n18257, new_n18258, new_n18259, new_n18260, new_n18261, new_n18262, new_n18263, new_n18264, new_n18265, new_n18266, new_n18267, new_n18268, new_n18269, new_n18270, new_n18271, new_n18272, new_n18273, new_n18274, new_n18275, new_n18276, new_n18277, new_n18278, new_n18279, new_n18280, new_n18281, new_n18282, new_n18283, new_n18284, new_n18285, new_n18286, new_n18287, new_n18288, new_n18289, new_n18290, new_n18291, new_n18292, new_n18293, new_n18294, new_n18295, new_n18296, new_n18297, new_n18298, new_n18299, new_n18300, new_n18301, new_n18302, new_n18303, new_n18304, new_n18305, new_n18306, new_n18307, new_n18308, new_n18309, new_n18310, new_n18311, new_n18312, new_n18313, new_n18314, new_n18315, new_n18316, new_n18317, new_n18318, new_n18319, new_n18320, new_n18321, new_n18322, new_n18323, new_n18324, new_n18325, new_n18326, new_n18327, new_n18328, new_n18329, new_n18330, new_n18331, new_n18332, new_n18333, new_n18334, new_n18335, new_n18336, new_n18337, new_n18338, new_n18339, new_n18340, new_n18341, new_n18342, new_n18343, new_n18344, new_n18345, new_n18346, new_n18347, new_n18348, new_n18349, new_n18350, new_n18351, new_n18352, new_n18353, new_n18354, new_n18355, new_n18356, new_n18357, new_n18358, new_n18359, new_n18360, new_n18361, new_n18362, new_n18363, new_n18364, new_n18365, new_n18366, new_n18367, new_n18368, new_n18369, new_n18370, new_n18371, new_n18372, new_n18373, new_n18374, new_n18375, new_n18376, new_n18377, new_n18378, new_n18379, new_n18380, new_n18381, new_n18382, new_n18383, new_n18384, new_n18385, new_n18386, new_n18387, new_n18388, new_n18389, new_n18390, new_n18391, new_n18392, new_n18393, new_n18394, new_n18395, new_n18396, new_n18397, new_n18398, new_n18399, new_n18400, new_n18401, new_n18402, new_n18403, new_n18404, new_n18405, new_n18406, new_n18407, new_n18408, new_n18409, new_n18410, new_n18411, new_n18412, new_n18413, new_n18414, new_n18415, new_n18416, new_n18417, new_n18418, new_n18419, new_n18420, new_n18421, new_n18422, new_n18423, new_n18424, new_n18425, new_n18426, new_n18427, new_n18428, new_n18429, new_n18430, new_n18431, new_n18432, new_n18433, new_n18434, new_n18435, new_n18436, new_n18437, new_n18438, new_n18439, new_n18440, new_n18441, new_n18442, new_n18443, new_n18444, new_n18445, new_n18446, new_n18447, new_n18448, new_n18449, new_n18450, new_n18451, new_n18452, new_n18453, new_n18454, new_n18455, new_n18456, new_n18457, new_n18458, new_n18459, new_n18460, new_n18461, new_n18462, new_n18463, new_n18464, new_n18465, new_n18466, new_n18467, new_n18468, new_n18469, new_n18470, new_n18471, new_n18472, new_n18473, new_n18474, new_n18475, new_n18476, new_n18477, new_n18478, new_n18479, new_n18480, new_n18481, new_n18482, new_n18483, new_n18484, new_n18485, new_n18486, new_n18487, new_n18488, new_n18489, new_n18490, new_n18491, new_n18492, new_n18493, new_n18494, new_n18495, new_n18496, new_n18497, new_n18498, new_n18499, new_n18500, new_n18501, new_n18502, new_n18503, new_n18504, new_n18505, new_n18506, new_n18507, new_n18508, new_n18509, new_n18510, new_n18511, new_n18512, new_n18513, new_n18514, new_n18515, new_n18516, new_n18517, new_n18518, new_n18519, new_n18520, new_n18521, new_n18522, new_n18523, new_n18524, new_n18525, new_n18526, new_n18527, new_n18528, new_n18529, new_n18530, new_n18531, new_n18532, new_n18533, new_n18534, new_n18535, new_n18536, new_n18537, new_n18538, new_n18539, new_n18540, new_n18541, new_n18542, new_n18543, new_n18544, new_n18545, new_n18546, new_n18547, new_n18548, new_n18549, new_n18550, new_n18551, new_n18552, new_n18553, new_n18554, new_n18555, new_n18556, new_n18557, new_n18558, new_n18559, new_n18560, new_n18561, new_n18562, new_n18563, new_n18564, new_n18565, new_n18566, new_n18567, new_n18568, new_n18569, new_n18570, new_n18571, new_n18572, new_n18573, new_n18574, new_n18575, new_n18576, new_n18577, new_n18578, new_n18579, new_n18580, new_n18581, new_n18582, new_n18583, new_n18584, new_n18585, new_n18586, new_n18587, new_n18588, new_n18589, new_n18590, new_n18591, new_n18592, new_n18593, new_n18594, new_n18595, new_n18596, new_n18597, new_n18598, new_n18599, new_n18600, new_n18601, new_n18602, new_n18603, new_n18604, new_n18605, new_n18606, new_n18607, new_n18608, new_n18609, new_n18610, new_n18611, new_n18612, new_n18613, new_n18614, new_n18615, new_n18616, new_n18617, new_n18618, new_n18619, new_n18620, new_n18621, new_n18622, new_n18623, new_n18624, new_n18625, new_n18626, new_n18627, new_n18628, new_n18629, new_n18630, new_n18631, new_n18632, new_n18633, new_n18634, new_n18635, new_n18636, new_n18637, new_n18638, new_n18639, new_n18640, new_n18641, new_n18642, new_n18643, new_n18644, new_n18645, new_n18646, new_n18647, new_n18648, new_n18649, new_n18650, new_n18651, new_n18652, new_n18653, new_n18654, new_n18655, new_n18656, new_n18657, new_n18658, new_n18659, new_n18660, new_n18661, new_n18662, new_n18663, new_n18664, new_n18665, new_n18666, new_n18667, new_n18668, new_n18669, new_n18670, new_n18671, new_n18672, new_n18673, new_n18674, new_n18675, new_n18676, new_n18677, new_n18678, new_n18679, new_n18680, new_n18681, new_n18682, new_n18683, new_n18684, new_n18685, new_n18686, new_n18687, new_n18688, new_n18689, new_n18690, new_n18691, new_n18692, new_n18693, new_n18694, new_n18695, new_n18696, new_n18697, new_n18698, new_n18699, new_n18700, new_n18701, new_n18702, new_n18703, new_n18704, new_n18705, new_n18706, new_n18707, new_n18708, new_n18709, new_n18710, new_n18711, new_n18712, new_n18713, new_n18714, new_n18715, new_n18716, new_n18717, new_n18718, new_n18719, new_n18720, new_n18721, new_n18722, new_n18723, new_n18724, new_n18725, new_n18726, new_n18727, new_n18728, new_n18729, new_n18730, new_n18731, new_n18732, new_n18733, new_n18734, new_n18735, new_n18736, new_n18737, new_n18738, new_n18739, new_n18740, new_n18741, new_n18742, new_n18743, new_n18744, new_n18745, new_n18746, new_n18747, new_n18748, new_n18749, new_n18750, new_n18751, new_n18752, new_n18753, new_n18754, new_n18755, new_n18756, new_n18757, new_n18758, new_n18759, new_n18760, new_n18761, new_n18762, new_n18763, new_n18764, new_n18765, new_n18766, new_n18767, new_n18768, new_n18769, new_n18770, new_n18771, new_n18772, new_n18773, new_n18774, new_n18775, new_n18776, new_n18777, new_n18778, new_n18779, new_n18780, new_n18781, new_n18782, new_n18783, new_n18784, new_n18785, new_n18786, new_n18787, new_n18788, new_n18789, new_n18790, new_n18791, new_n18792, new_n18793, new_n18794, new_n18795, new_n18796, new_n18797, new_n18798, new_n18799, new_n18800, new_n18801, new_n18802, new_n18803, new_n18804, new_n18805, new_n18806, new_n18807, new_n18808, new_n18809, new_n18810, new_n18811, new_n18812, new_n18813, new_n18814, new_n18815, new_n18816, new_n18817, new_n18818, new_n18819, new_n18820, new_n18821, new_n18822, new_n18823, new_n18824, new_n18825, new_n18826, new_n18827, new_n18828, new_n18829, new_n18830, new_n18831, new_n18832, new_n18833, new_n18834, new_n18835, new_n18836, new_n18837, new_n18838, new_n18839, new_n18840, new_n18841, new_n18842, new_n18843, new_n18844, new_n18845, new_n18846, new_n18847, new_n18848, new_n18849, new_n18850, new_n18851, new_n18852, new_n18853, new_n18854, new_n18855, new_n18856, new_n18857, new_n18858, new_n18859, new_n18860, new_n18861, new_n18862, new_n18863, new_n18864, new_n18865, new_n18866, new_n18867, new_n18868, new_n18869, new_n18870, new_n18871, new_n18872, new_n18873, new_n18874, new_n18875, new_n18876, new_n18877, new_n18878, new_n18879, new_n18880, new_n18881, new_n18882, new_n18883, new_n18884, new_n18885, new_n18886, new_n18887, new_n18888, new_n18889, new_n18890, new_n18891, new_n18892, new_n18893, new_n18894, new_n18895, new_n18896, new_n18897, new_n18898, new_n18899, new_n18900, new_n18901, new_n18902, new_n18903, new_n18904, new_n18905, new_n18906, new_n18907, new_n18908, new_n18909, new_n18910, new_n18911, new_n18912, new_n18913, new_n18914, new_n18915, new_n18916, new_n18917, new_n18918, new_n18919, new_n18920, new_n18921, new_n18922, new_n18923, new_n18924, new_n18925, new_n18926, new_n18927, new_n18928, new_n18929, new_n18930, new_n18931, new_n18932, new_n18933, new_n18934, new_n18935, new_n18936, new_n18937, new_n18938, new_n18939, new_n18940, new_n18941, new_n18942, new_n18943, new_n18944, new_n18945, new_n18946, new_n18947, new_n18948, new_n18949, new_n18950, new_n18951, new_n18952, new_n18953, new_n18954, new_n18955, new_n18956, new_n18957, new_n18958, new_n18959, new_n18960, new_n18961, new_n18962, new_n18963, new_n18964, new_n18965, new_n18966, new_n18967, new_n18968, new_n18969, new_n18970, new_n18971, new_n18972, new_n18973, new_n18974, new_n18975, new_n18976, new_n18977, new_n18978, new_n18979, new_n18980, new_n18981, new_n18982, new_n18983, new_n18984, new_n18985, new_n18986, new_n18987, new_n18988, new_n18989, new_n18990, new_n18991, new_n18992, new_n18993, new_n18994, new_n18995, new_n18996, new_n18997, new_n18998, new_n18999, new_n19000, new_n19001, new_n19002, new_n19003, new_n19004, new_n19005, new_n19006, new_n19007, new_n19008, new_n19009, new_n19010, new_n19011, new_n19012, new_n19013, new_n19014, new_n19015, new_n19016, new_n19017, new_n19018, new_n19019, new_n19020, new_n19021, new_n19022, new_n19023, new_n19024, new_n19025, new_n19026, new_n19027, new_n19028, new_n19029, new_n19030, new_n19031, new_n19032, new_n19033, new_n19034, new_n19035, new_n19036, new_n19037, new_n19038, new_n19039, new_n19040, new_n19041, new_n19042, new_n19043, new_n19044, new_n19045, new_n19046, new_n19047, new_n19048, new_n19049, new_n19050, new_n19051, new_n19052, new_n19053, new_n19054, new_n19055, new_n19056, new_n19057, new_n19058, new_n19059, new_n19060, new_n19061, new_n19062, new_n19063, new_n19064, new_n19065, new_n19066, new_n19067, new_n19068, new_n19069, new_n19070, new_n19071, new_n19072, new_n19073, new_n19074, new_n19075, new_n19076, new_n19077, new_n19078, new_n19079, new_n19080, new_n19081, new_n19082, new_n19083, new_n19084, new_n19085, new_n19086, new_n19087, new_n19088, new_n19089, new_n19090, new_n19091, new_n19092, new_n19093, new_n19094, new_n19095, new_n19096, new_n19097, new_n19098, new_n19099, new_n19100, new_n19101, new_n19102, new_n19103, new_n19104, new_n19105, new_n19106, new_n19107, new_n19108, new_n19109, new_n19110, new_n19111, new_n19112, new_n19113, new_n19114, new_n19115, new_n19116, new_n19117, new_n19118, new_n19119, new_n19120, new_n19121, new_n19122, new_n19123, new_n19124, new_n19125, new_n19126, new_n19127, new_n19128, new_n19129, new_n19130, new_n19131, new_n19132, new_n19133, new_n19134, new_n19135, new_n19136, new_n19137, new_n19138, new_n19139, new_n19140, new_n19141, new_n19142, new_n19143, new_n19144, new_n19145, new_n19146, new_n19147, new_n19148, new_n19149, new_n19150, new_n19151, new_n19152, new_n19153, new_n19154, new_n19155, new_n19156, new_n19157, new_n19158, new_n19159, new_n19160, new_n19161, new_n19162, new_n19163, new_n19164, new_n19165, new_n19166, new_n19167, new_n19168, new_n19169, new_n19170, new_n19171, new_n19172, new_n19173, new_n19174, new_n19175, new_n19176, new_n19177, new_n19178, new_n19179, new_n19180, new_n19181, new_n19182, new_n19183, new_n19184, new_n19185, new_n19186, new_n19187, new_n19188, new_n19189, new_n19190, new_n19191, new_n19192, new_n19193, new_n19194, new_n19195, new_n19196, new_n19197, new_n19198, new_n19199, new_n19200, new_n19201, new_n19202, new_n19203, new_n19204, new_n19205, new_n19206, new_n19207, new_n19208, new_n19209, new_n19210, new_n19211, new_n19212, new_n19213, new_n19214, new_n19215, new_n19216, new_n19217, new_n19218, new_n19219, new_n19220, new_n19221, new_n19222, new_n19223, new_n19224, new_n19225, new_n19226, new_n19227, new_n19228, new_n19229, new_n19230, new_n19231, new_n19232, new_n19233, new_n19234, new_n19235, new_n19236, new_n19237, new_n19238, new_n19239, new_n19240, new_n19241, new_n19242, new_n19243, new_n19244, new_n19245, new_n19246, new_n19247, new_n19248, new_n19249, new_n19250, new_n19251, new_n19252, new_n19253, new_n19254, new_n19255, new_n19256, new_n19257, new_n19258, new_n19259, new_n19260, new_n19261, new_n19262, new_n19263, new_n19264, new_n19265, new_n19266, new_n19267, new_n19268, new_n19269, new_n19270, new_n19271, new_n19272, new_n19273, new_n19274, new_n19275, new_n19276, new_n19277, new_n19278, new_n19279, new_n19280, new_n19281, new_n19282, new_n19283, new_n19284, new_n19285, new_n19286, new_n19287, new_n19288, new_n19289, new_n19290, new_n19291, new_n19292, new_n19293, new_n19294, new_n19295, new_n19296, new_n19297, new_n19298, new_n19299, new_n19300, new_n19301, new_n19302, new_n19303, new_n19304, new_n19305, new_n19306, new_n19307, new_n19308, new_n19309, new_n19310, new_n19311, new_n19312, new_n19313, new_n19314, new_n19315, new_n19316, new_n19317, new_n19318, new_n19319, new_n19320, new_n19321, new_n19322, new_n19323, new_n19324, new_n19325, new_n19326, new_n19327, new_n19328, new_n19329, new_n19330, new_n19331, new_n19332, new_n19333, new_n19334, new_n19335, new_n19336, new_n19337, new_n19338, new_n19339, new_n19340, new_n19341, new_n19342, new_n19343, new_n19344, new_n19345, new_n19346, new_n19347, new_n19348, new_n19349, new_n19350, new_n19351, new_n19352, new_n19353, new_n19354, new_n19355, new_n19356, new_n19357, new_n19358, new_n19359, new_n19360, new_n19361, new_n19362, new_n19363, new_n19364, new_n19365, new_n19366, new_n19367, new_n19368, new_n19369, new_n19370, new_n19371, new_n19372, new_n19373, new_n19374, new_n19375, new_n19376, new_n19377, new_n19378, new_n19379, new_n19380, new_n19381, new_n19382, new_n19383, new_n19384, new_n19385, new_n19386, new_n19387, new_n19388, new_n19389, new_n19390, new_n19391, new_n19392, new_n19393, new_n19394, new_n19395, new_n19396, new_n19397, new_n19398, new_n19399, new_n19400, new_n19401, new_n19402, new_n19403, new_n19404, new_n19405, new_n19406, new_n19407, new_n19408, new_n19409, new_n19410, new_n19411, new_n19412, new_n19413, new_n19414, new_n19415, new_n19416, new_n19417, new_n19418, new_n19419, new_n19420, new_n19421, new_n19422, new_n19423, new_n19424, new_n19425, new_n19426, new_n19427, new_n19428, new_n19429, new_n19430, new_n19431, new_n19432, new_n19433, new_n19434, new_n19435, new_n19436, new_n19437, new_n19438, new_n19439, new_n19440, new_n19441, new_n19442, new_n19443, new_n19444, new_n19445, new_n19446, new_n19447, new_n19448, new_n19449, new_n19450, new_n19451, new_n19452, new_n19453, new_n19454, new_n19455, new_n19456, new_n19457, new_n19458, new_n19459, new_n19460, new_n19461, new_n19462, new_n19463, new_n19464, new_n19465, new_n19466, new_n19467, new_n19468, new_n19469, new_n19470, new_n19471, new_n19472, new_n19473, new_n19474, new_n19475, new_n19476, new_n19477, new_n19478, new_n19479, new_n19480, new_n19481, new_n19482, new_n19483, new_n19484, new_n19485, new_n19486, new_n19487, new_n19488, new_n19489, new_n19490, new_n19491, new_n19492, new_n19493, new_n19494, new_n19495, new_n19496, new_n19497, new_n19498, new_n19499, new_n19500, new_n19501, new_n19502, new_n19503, new_n19504, new_n19505, new_n19506, new_n19507, new_n19508, new_n19509, new_n19510, new_n19511, new_n19512, new_n19513, new_n19514, new_n19515, new_n19516, new_n19517, new_n19518, new_n19519, new_n19520, new_n19521, new_n19522, new_n19523, new_n19524, new_n19525, new_n19526, new_n19527, new_n19528, new_n19529, new_n19530, new_n19531, new_n19532, new_n19533, new_n19534, new_n19535, new_n19536, new_n19537, new_n19538, new_n19539, new_n19540, new_n19541, new_n19542, new_n19543, new_n19544, new_n19545, new_n19546, new_n19547, new_n19548, new_n19549, new_n19550, new_n19551, new_n19552, new_n19553, new_n19554, new_n19555, new_n19556, new_n19557, new_n19558, new_n19559, new_n19560, new_n19561, new_n19562, new_n19563, new_n19564, new_n19565, new_n19566, new_n19567, new_n19568, new_n19569, new_n19570, new_n19571, new_n19572, new_n19573, new_n19574, new_n19575, new_n19576, new_n19577, new_n19578, new_n19579, new_n19580, new_n19581, new_n19582, new_n19583, new_n19584, new_n19585, new_n19586, new_n19587, new_n19588, new_n19589, new_n19590, new_n19591, new_n19592, new_n19593, new_n19594, new_n19595, new_n19596, new_n19597, new_n19598, new_n19599, new_n19600, new_n19601, new_n19602, new_n19603, new_n19604, new_n19605, new_n19606, new_n19607, new_n19608, new_n19609, new_n19610, new_n19611, new_n19612, new_n19613, new_n19614, new_n19615, new_n19616, new_n19617, new_n19618, new_n19619, new_n19620, new_n19621, new_n19622, new_n19623, new_n19624, new_n19625, new_n19626, new_n19627, new_n19628, new_n19629, new_n19630, new_n19631, new_n19632, new_n19633, new_n19634, new_n19635, new_n19636, new_n19637, new_n19638, new_n19639, new_n19640, new_n19641, new_n19642, new_n19643, new_n19644, new_n19645, new_n19646, new_n19647, new_n19648, new_n19649, new_n19650, new_n19651, new_n19652, new_n19653, new_n19654, new_n19655, new_n19656, new_n19657, new_n19658, new_n19659, new_n19660, new_n19661, new_n19662, new_n19663, new_n19664, new_n19665, new_n19666, new_n19667, new_n19668, new_n19669, new_n19670, new_n19671, new_n19672, new_n19673, new_n19674, new_n19675, new_n19676, new_n19677, new_n19678, new_n19679, new_n19680, new_n19681, new_n19682, new_n19683, new_n19684, new_n19685, new_n19686, new_n19687, new_n19688, new_n19689, new_n19690, new_n19691, new_n19692, new_n19693, new_n19694, new_n19695, new_n19696, new_n19697, new_n19698, new_n19699, new_n19700, new_n19701, new_n19702, new_n19703, new_n19704, new_n19705, new_n19706, new_n19707, new_n19708, new_n19709, new_n19710, new_n19711, new_n19712, new_n19713, new_n19714, new_n19715, new_n19716, new_n19717, new_n19718, new_n19719, new_n19720, new_n19721, new_n19722, new_n19723, new_n19724, new_n19725, new_n19726, new_n19727, new_n19728, new_n19729, new_n19730, new_n19731, new_n19732, new_n19733, new_n19734, new_n19735, new_n19736, new_n19737, new_n19738, new_n19739, new_n19740, new_n19741, new_n19742, new_n19743, new_n19744, new_n19745, new_n19746, new_n19747, new_n19748, new_n19749, new_n19750, new_n19751, new_n19752, new_n19753, new_n19754, new_n19755, new_n19756, new_n19757, new_n19758, new_n19759, new_n19760, new_n19761, new_n19762, new_n19763, new_n19764, new_n19765, new_n19766, new_n19767, new_n19768, new_n19769, new_n19770, new_n19771, new_n19772, new_n19773, new_n19774, new_n19775, new_n19776, new_n19777, new_n19778, new_n19779, new_n19780, new_n19781, new_n19782, new_n19783, new_n19784, new_n19785, new_n19786, new_n19787, new_n19788, new_n19789, new_n19790, new_n19791, new_n19792, new_n19793, new_n19794, new_n19795, new_n19796, new_n19797, new_n19798, new_n19799, new_n19800, new_n19801, new_n19802, new_n19803, new_n19804, new_n19805, new_n19806, new_n19807, new_n19808, new_n19809, new_n19810, new_n19811, new_n19812, new_n19813, new_n19814, new_n19815, new_n19816, new_n19817, new_n19818, new_n19819, new_n19820, new_n19821, new_n19822, new_n19823, new_n19824, new_n19825, new_n19826, new_n19827, new_n19828, new_n19829, new_n19830, new_n19831, new_n19832, new_n19833, new_n19834, new_n19835, new_n19836, new_n19837, new_n19838, new_n19839, new_n19840, new_n19841, new_n19842, new_n19843, new_n19844, new_n19845, new_n19846, new_n19847, new_n19848, new_n19849, new_n19850, new_n19851, new_n19852, new_n19853, new_n19854, new_n19855, new_n19856, new_n19857, new_n19858, new_n19859, new_n19860, new_n19861, new_n19862, new_n19863, new_n19864, new_n19865, new_n19866, new_n19867, new_n19868, new_n19869, new_n19870, new_n19871, new_n19872, new_n19873, new_n19874, new_n19875, new_n19876, new_n19877, new_n19878, new_n19879, new_n19880, new_n19881, new_n19882, new_n19883, new_n19884, new_n19885, new_n19886, new_n19887, new_n19888, new_n19889, new_n19890, new_n19891, new_n19892, new_n19893, new_n19894, new_n19895, new_n19896, new_n19897, new_n19898, new_n19899, new_n19900, new_n19901, new_n19902, new_n19903, new_n19904, new_n19905, new_n19906, new_n19907, new_n19908, new_n19909, new_n19910, new_n19911, new_n19912, new_n19913, new_n19914, new_n19915, new_n19916, new_n19917, new_n19918, new_n19919, new_n19920, new_n19921, new_n19922, new_n19923, new_n19924, new_n19925, new_n19926, new_n19927, new_n19928, new_n19929, new_n19930, new_n19931, new_n19932, new_n19933, new_n19934, new_n19935, new_n19936, new_n19937, new_n19938, new_n19939, new_n19940, new_n19941, new_n19942, new_n19943, new_n19944, new_n19945, new_n19946, new_n19947, new_n19948, new_n19949, new_n19950, new_n19951, new_n19952, new_n19953, new_n19954, new_n19955, new_n19956, new_n19957, new_n19958, new_n19959, new_n19960, new_n19961, new_n19962, new_n19963, new_n19964, new_n19965, new_n19966, new_n19967, new_n19968, new_n19969, new_n19970, new_n19971, new_n19972, new_n19973, new_n19974, new_n19975, new_n19976, new_n19977, new_n19978, new_n19979, new_n19980, new_n19981, new_n19982, new_n19983, new_n19984, new_n19985, new_n19986, new_n19987, new_n19988, new_n19989, new_n19990, new_n19991, new_n19992, new_n19993, new_n19994, new_n19995, new_n19996, new_n19997, new_n19998, new_n19999, new_n20000, new_n20001, new_n20002, new_n20003, new_n20004, new_n20005, new_n20006, new_n20007, new_n20008, new_n20009, new_n20010, new_n20011, new_n20012, new_n20013, new_n20014, new_n20015, new_n20016, new_n20017, new_n20018, new_n20019, new_n20020, new_n20021, new_n20022, new_n20023, new_n20024, new_n20025, new_n20026, new_n20027, new_n20028, new_n20029, new_n20030, new_n20031, new_n20032, new_n20033, new_n20034, new_n20035, new_n20036, new_n20037, new_n20038, new_n20039, new_n20040, new_n20041, new_n20042, new_n20043, new_n20044, new_n20045, new_n20046, new_n20047, new_n20048, new_n20049, new_n20050, new_n20051, new_n20052, new_n20053, new_n20054, new_n20055, new_n20056, new_n20057, new_n20058, new_n20059, new_n20060, new_n20061, new_n20062, new_n20063, new_n20064, new_n20065, new_n20066, new_n20067, new_n20068, new_n20069, new_n20070, new_n20071, new_n20072, new_n20073, new_n20074, new_n20075, new_n20076, new_n20077, new_n20078, new_n20079, new_n20080, new_n20081, new_n20082, new_n20083, new_n20084, new_n20085, new_n20086, new_n20087, new_n20088, new_n20089, new_n20090, new_n20091, new_n20092, new_n20093, new_n20094, new_n20095, new_n20096, new_n20097, new_n20098, new_n20099, new_n20100, new_n20101, new_n20102, new_n20103, new_n20104, new_n20105, new_n20106, new_n20107, new_n20108, new_n20109, new_n20110, new_n20111, new_n20112, new_n20113, new_n20114, new_n20115, new_n20116, new_n20117, new_n20118, new_n20119, new_n20120, new_n20121, new_n20122, new_n20123, new_n20124, new_n20125, new_n20126, new_n20127, new_n20128, new_n20129, new_n20130, new_n20131, new_n20132, new_n20133, new_n20134, new_n20135, new_n20136, new_n20137, new_n20138, new_n20139, new_n20140, new_n20141, new_n20142, new_n20143, new_n20144, new_n20145, new_n20146, new_n20147, new_n20148, new_n20149, new_n20150, new_n20151, new_n20152, new_n20153, new_n20154, new_n20155, new_n20156, new_n20157, new_n20158, new_n20159, new_n20160, new_n20161, new_n20162, new_n20163, new_n20164, new_n20165, new_n20166, new_n20167, new_n20168, new_n20169, new_n20170, new_n20171, new_n20172, new_n20173, new_n20174, new_n20175, new_n20176, new_n20177, new_n20178, new_n20179, new_n20180, new_n20181, new_n20182, new_n20183, new_n20184, new_n20185, new_n20186, new_n20187, new_n20188, new_n20189, new_n20190, new_n20191, new_n20192, new_n20193, new_n20194, new_n20195, new_n20196, new_n20197, new_n20198, new_n20199, new_n20200, new_n20201, new_n20202, new_n20203, new_n20204, new_n20205, new_n20206, new_n20207, new_n20208, new_n20209, new_n20210, new_n20211, new_n20212, new_n20213, new_n20214, new_n20215, new_n20216, new_n20217, new_n20218, new_n20219, new_n20220, new_n20221, new_n20222, new_n20223, new_n20224, new_n20225, new_n20226, new_n20227, new_n20228, new_n20229, new_n20230, new_n20231, new_n20232, new_n20233, new_n20234, new_n20235, new_n20236, new_n20237, new_n20238, new_n20239, new_n20240, new_n20241, new_n20242, new_n20243, new_n20244, new_n20245, new_n20246, new_n20247, new_n20248, new_n20249, new_n20250, new_n20251, new_n20252, new_n20253, new_n20254, new_n20255, new_n20256, new_n20257, new_n20258, new_n20259, new_n20260, new_n20261, new_n20262, new_n20263, new_n20264, new_n20265, new_n20266, new_n20267, new_n20268, new_n20269, new_n20270, new_n20271, new_n20272, new_n20273, new_n20274, new_n20275, new_n20276, new_n20277, new_n20278, new_n20279, new_n20280, new_n20281, new_n20282, new_n20283, new_n20284, new_n20285, new_n20286, new_n20287, new_n20288, new_n20289, new_n20290, new_n20291, new_n20292, new_n20293, new_n20294, new_n20295, new_n20296, new_n20297, new_n20298, new_n20299, new_n20300, new_n20301, new_n20302, new_n20303, new_n20304, new_n20305, new_n20306, new_n20307, new_n20308, new_n20309, new_n20310, new_n20311, new_n20312, new_n20313, new_n20314, new_n20315, new_n20316, new_n20317, new_n20318, new_n20319, new_n20320, new_n20321, new_n20322, new_n20323, new_n20324, new_n20325, new_n20326, new_n20327, new_n20328, new_n20329, new_n20330, new_n20331, new_n20332, new_n20333, new_n20334, new_n20335, new_n20336, new_n20337, new_n20338, new_n20339, new_n20340, new_n20341, new_n20342, new_n20343, new_n20344, new_n20345, new_n20346, new_n20347, new_n20348, new_n20349, new_n20350, new_n20351, new_n20352, new_n20353, new_n20354, new_n20355, new_n20356, new_n20357, new_n20358, new_n20359, new_n20360, new_n20361, new_n20362, new_n20363, new_n20364, new_n20365, new_n20366, new_n20367, new_n20368, new_n20369, new_n20370, new_n20371, new_n20372, new_n20373, new_n20374, new_n20375, new_n20376, new_n20377, new_n20378, new_n20379, new_n20380, new_n20381, new_n20382, new_n20383, new_n20384, new_n20385, new_n20386, new_n20387, new_n20388, new_n20389, new_n20390, new_n20391, new_n20392, new_n20393, new_n20394, new_n20395, new_n20396, new_n20397, new_n20398, new_n20399, new_n20400, new_n20401, new_n20402, new_n20403, new_n20404, new_n20405, new_n20406, new_n20407, new_n20408, new_n20409, new_n20410, new_n20411, new_n20412, new_n20413, new_n20414, new_n20415, new_n20416, new_n20417, new_n20418, new_n20419, new_n20420, new_n20421, new_n20422, new_n20423, new_n20424, new_n20425, new_n20426, new_n20427, new_n20428, new_n20429, new_n20430, new_n20431, new_n20432, new_n20433, new_n20434, new_n20435, new_n20436, new_n20437, new_n20438, new_n20439, new_n20440, new_n20441, new_n20442, new_n20443, new_n20444, new_n20445, new_n20446, new_n20447, new_n20448, new_n20449, new_n20450, new_n20451, new_n20452, new_n20453, new_n20454, new_n20455, new_n20456, new_n20457, new_n20458, new_n20459, new_n20460, new_n20461, new_n20462, new_n20463, new_n20464, new_n20465, new_n20466, new_n20467, new_n20468, new_n20469, new_n20470, new_n20471, new_n20472, new_n20473, new_n20474, new_n20475, new_n20476, new_n20477, new_n20478, new_n20479, new_n20480, new_n20481, new_n20482, new_n20483, new_n20484, new_n20485, new_n20486, new_n20487, new_n20488, new_n20489, new_n20490, new_n20491, new_n20492, new_n20493, new_n20494, new_n20495, new_n20496, new_n20497, new_n20498, new_n20499, new_n20500, new_n20501, new_n20502, new_n20503, new_n20504, new_n20505, new_n20506, new_n20507, new_n20508, new_n20509, new_n20510, new_n20511, new_n20512, new_n20513, new_n20514, new_n20515, new_n20516, new_n20517, new_n20518, new_n20519, new_n20520, new_n20521, new_n20522, new_n20523, new_n20524, new_n20525, new_n20526, new_n20527, new_n20528, new_n20529, new_n20530, new_n20531, new_n20532, new_n20533, new_n20534, new_n20535, new_n20536, new_n20537, new_n20538, new_n20539, new_n20540, new_n20541, new_n20542, new_n20543, new_n20544, new_n20545, new_n20546, new_n20547, new_n20548, new_n20549, new_n20550, new_n20551, new_n20552, new_n20553, new_n20554, new_n20555, new_n20556, new_n20557, new_n20558, new_n20559, new_n20560, new_n20561, new_n20562, new_n20563, new_n20564, new_n20565, new_n20566, new_n20567, new_n20568, new_n20569, new_n20570, new_n20571, new_n20572, new_n20573, new_n20574, new_n20575, new_n20576, new_n20577, new_n20578, new_n20579, new_n20580, new_n20581, new_n20582, new_n20583, new_n20584, new_n20585, new_n20586, new_n20587, new_n20588, new_n20589, new_n20590, new_n20591, new_n20592, new_n20593, new_n20594, new_n20595, new_n20596, new_n20597, new_n20598, new_n20599, new_n20600, new_n20601, new_n20602, new_n20603, new_n20604, new_n20605, new_n20606, new_n20607, new_n20608, new_n20609, new_n20610, new_n20611, new_n20612, new_n20613, new_n20614, new_n20615, new_n20616, new_n20617, new_n20618, new_n20619, new_n20620, new_n20621, new_n20622, new_n20623, new_n20624, new_n20625, new_n20626, new_n20627, new_n20628, new_n20629, new_n20630, new_n20631, new_n20632, new_n20633, new_n20634, new_n20635, new_n20636, new_n20637, new_n20638, new_n20639, new_n20640, new_n20641, new_n20642, new_n20643, new_n20644, new_n20645, new_n20646, new_n20647, new_n20648, new_n20649, new_n20650, new_n20651, new_n20652, new_n20653, new_n20654, new_n20655, new_n20656, new_n20657, new_n20658, new_n20659, new_n20660, new_n20661, new_n20662, new_n20663, new_n20664, new_n20665, new_n20666, new_n20667, new_n20668, new_n20669, new_n20670, new_n20671, new_n20672, new_n20673, new_n20674, new_n20675, new_n20676, new_n20677, new_n20678, new_n20679, new_n20680, new_n20681, new_n20682, new_n20683, new_n20684, new_n20685, new_n20686, new_n20687, new_n20688, new_n20689, new_n20690, new_n20691, new_n20692, new_n20693, new_n20694, new_n20695, new_n20696, new_n20697, new_n20698, new_n20699, new_n20700, new_n20701, new_n20702, new_n20703, new_n20704, new_n20705, new_n20706, new_n20707, new_n20708, new_n20709, new_n20710, new_n20711, new_n20712, new_n20713, new_n20714, new_n20715, new_n20716, new_n20717, new_n20718, new_n20719, new_n20720, new_n20721, new_n20722, new_n20723, new_n20724, new_n20725, new_n20726, new_n20727, new_n20728, new_n20729, new_n20730, new_n20731, new_n20732, new_n20733, new_n20734, new_n20735, new_n20736, new_n20737, new_n20738, new_n20739, new_n20740, new_n20741, new_n20742, new_n20743, new_n20744, new_n20745, new_n20746, new_n20747, new_n20748, new_n20749, new_n20750, new_n20751, new_n20752, new_n20753, new_n20754, new_n20755, new_n20756, new_n20757, new_n20758, new_n20759, new_n20760, new_n20761, new_n20762, new_n20763, new_n20764, new_n20765, new_n20766, new_n20767, new_n20768, new_n20769, new_n20770, new_n20771, new_n20772, new_n20773, new_n20774, new_n20775, new_n20776, new_n20777, new_n20778, new_n20779, new_n20780, new_n20781, new_n20782, new_n20783, new_n20784, new_n20785, new_n20786, new_n20787, new_n20788, new_n20789, new_n20790, new_n20791, new_n20792, new_n20793, new_n20794, new_n20795, new_n20796, new_n20797, new_n20798, new_n20799, new_n20800, new_n20801, new_n20802, new_n20803, new_n20804, new_n20805, new_n20806, new_n20807, new_n20808, new_n20809, new_n20810, new_n20811, new_n20812, new_n20813, new_n20814, new_n20815, new_n20816, new_n20817, new_n20818, new_n20819, new_n20820, new_n20821, new_n20822, new_n20823, new_n20824, new_n20825, new_n20826, new_n20827, new_n20828, new_n20829, new_n20830, new_n20831, new_n20832, new_n20833, new_n20834, new_n20835, new_n20836, new_n20837, new_n20838, new_n20839, new_n20840, new_n20841, new_n20842, new_n20843, new_n20844, new_n20845, new_n20846, new_n20847, new_n20848, new_n20849, new_n20850, new_n20851, new_n20852, new_n20853, new_n20854, new_n20855, new_n20856, new_n20857, new_n20858, new_n20859, new_n20860, new_n20861, new_n20862, new_n20863, new_n20864, new_n20865, new_n20866, new_n20867, new_n20868, new_n20869, new_n20870, new_n20871, new_n20872, new_n20873, new_n20874, new_n20875, new_n20876, new_n20877, new_n20878, new_n20879, new_n20880, new_n20881, new_n20882, new_n20883, new_n20884, new_n20885, new_n20886, new_n20887, new_n20888, new_n20889, new_n20890, new_n20891, new_n20892, new_n20893, new_n20894, new_n20895, new_n20896, new_n20897, new_n20898, new_n20899, new_n20900, new_n20901, new_n20902, new_n20903, new_n20904, new_n20905, new_n20906, new_n20907, new_n20908, new_n20909, new_n20910, new_n20911, new_n20912, new_n20913, new_n20914, new_n20915, new_n20916, new_n20917, new_n20918, new_n20919, new_n20920, new_n20921, new_n20922, new_n20923, new_n20924, new_n20925, new_n20926, new_n20927, new_n20928, new_n20929, new_n20930, new_n20931, new_n20932, new_n20933, new_n20934, new_n20935, new_n20936, new_n20937, new_n20938, new_n20939, new_n20940, new_n20941, new_n20942, new_n20943, new_n20944, new_n20945, new_n20946, new_n20947, new_n20948, new_n20949, new_n20950, new_n20951, new_n20952, new_n20953, new_n20954, new_n20955, new_n20956, new_n20957, new_n20958, new_n20959, new_n20960, new_n20961, new_n20962, new_n20963, new_n20964, new_n20965, new_n20966, new_n20967, new_n20968, new_n20969, new_n20970, new_n20971, new_n20972, new_n20973, new_n20974, new_n20975, new_n20976, new_n20977, new_n20978, new_n20979, new_n20980, new_n20981, new_n20982, new_n20983, new_n20984, new_n20985, new_n20986, new_n20987, new_n20988, new_n20989, new_n20990, new_n20991, new_n20992, new_n20993, new_n20994, new_n20995, new_n20996, new_n20997, new_n20998, new_n20999, new_n21000, new_n21001, new_n21002, new_n21003, new_n21004, new_n21005, new_n21006, new_n21007, new_n21008, new_n21009, new_n21010, new_n21011, new_n21012, new_n21013, new_n21014, new_n21015, new_n21016, new_n21017, new_n21018, new_n21019, new_n21020, new_n21021, new_n21022, new_n21023, new_n21024, new_n21025, new_n21026, new_n21027, new_n21028, new_n21029, new_n21030, new_n21031, new_n21032, new_n21033, new_n21034, new_n21035, new_n21036, new_n21037, new_n21038, new_n21039, new_n21040, new_n21041, new_n21042, new_n21043, new_n21044, new_n21045, new_n21046, new_n21047, new_n21048, new_n21049, new_n21050, new_n21051, new_n21052, new_n21053, new_n21054, new_n21055, new_n21056, new_n21057, new_n21058, new_n21059, new_n21060, new_n21061, new_n21062, new_n21063, new_n21064, new_n21065, new_n21066, new_n21067, new_n21068, new_n21069, new_n21070, new_n21071, new_n21072, new_n21073, new_n21074, new_n21075, new_n21076, new_n21077, new_n21078, new_n21079, new_n21080, new_n21081, new_n21082, new_n21083, new_n21084, new_n21085, new_n21086, new_n21087, new_n21088, new_n21089, new_n21090, new_n21091, new_n21092, new_n21093, new_n21094, new_n21095, new_n21096, new_n21097, new_n21098, new_n21099, new_n21100, new_n21101, new_n21102, new_n21103, new_n21104, new_n21105, new_n21106, new_n21107, new_n21108, new_n21109, new_n21110, new_n21111, new_n21112, new_n21113, new_n21114, new_n21115, new_n21116, new_n21117, new_n21118, new_n21119, new_n21120, new_n21121, new_n21122, new_n21123, new_n21124, new_n21125, new_n21126, new_n21127, new_n21128, new_n21129, new_n21130, new_n21131, new_n21132, new_n21133, new_n21134, new_n21135, new_n21136, new_n21137, new_n21138, new_n21139, new_n21140, new_n21141, new_n21142, new_n21143, new_n21144, new_n21145, new_n21146, new_n21147, new_n21148, new_n21149, new_n21150, new_n21151, new_n21152, new_n21153, new_n21154, new_n21155, new_n21156, new_n21157, new_n21158, new_n21159, new_n21160, new_n21161, new_n21162, new_n21163, new_n21164, new_n21165, new_n21166, new_n21167, new_n21168, new_n21169, new_n21170, new_n21171, new_n21172, new_n21173, new_n21174, new_n21175, new_n21176, new_n21177, new_n21178, new_n21179, new_n21180, new_n21181, new_n21182, new_n21183, new_n21184, new_n21185, new_n21186, new_n21187, new_n21188, new_n21189, new_n21190, new_n21191, new_n21192, new_n21193, new_n21194, new_n21195, new_n21196, new_n21197, new_n21198, new_n21199, new_n21200, new_n21201, new_n21202, new_n21203, new_n21204, new_n21205, new_n21206, new_n21207, new_n21208, new_n21209, new_n21210, new_n21211, new_n21212, new_n21213, new_n21214, new_n21215, new_n21216, new_n21217, new_n21218, new_n21219, new_n21220, new_n21221, new_n21222, new_n21223, new_n21224, new_n21225, new_n21226, new_n21227, new_n21228, new_n21229, new_n21230, new_n21231, new_n21232, new_n21233, new_n21234, new_n21235, new_n21236, new_n21237, new_n21238, new_n21239, new_n21240, new_n21241, new_n21242, new_n21243, new_n21244, new_n21245, new_n21246, new_n21247, new_n21248, new_n21249, new_n21250, new_n21251, new_n21252, new_n21253, new_n21254, new_n21255, new_n21256, new_n21257, new_n21258, new_n21259, new_n21260, new_n21261, new_n21262, new_n21263, new_n21264, new_n21265, new_n21266, new_n21267, new_n21268, new_n21269, new_n21270, new_n21271, new_n21272, new_n21273, new_n21274, new_n21275, new_n21276, new_n21277, new_n21278, new_n21279, new_n21280, new_n21281, new_n21282, new_n21283, new_n21284, new_n21285, new_n21286, new_n21287, new_n21288, new_n21289, new_n21290, new_n21291, new_n21292, new_n21293, new_n21294, new_n21295, new_n21296, new_n21297, new_n21298, new_n21299, new_n21300, new_n21301, new_n21302, new_n21303, new_n21304, new_n21305, new_n21306, new_n21307, new_n21308, new_n21309, new_n21310, new_n21311, new_n21312, new_n21313, new_n21314, new_n21315, new_n21316, new_n21317, new_n21318, new_n21319, new_n21320, new_n21321, new_n21322, new_n21323, new_n21324, new_n21325, new_n21326, new_n21327, new_n21328, new_n21329, new_n21330, new_n21331, new_n21332, new_n21333, new_n21334, new_n21335, new_n21336, new_n21337, new_n21338, new_n21339, new_n21340, new_n21341, new_n21342, new_n21343, new_n21344, new_n21345, new_n21346, new_n21347, new_n21348, new_n21349, new_n21350, new_n21351, new_n21352, new_n21353, new_n21354, new_n21355, new_n21356, new_n21357, new_n21358, new_n21359, new_n21360, new_n21361, new_n21362, new_n21363, new_n21364, new_n21365, new_n21366, new_n21367, new_n21368, new_n21369, new_n21370, new_n21371, new_n21372, new_n21373, new_n21374, new_n21375, new_n21376, new_n21377, new_n21378, new_n21379, new_n21380, new_n21381, new_n21382, new_n21383, new_n21384, new_n21385, new_n21386, new_n21387, new_n21388, new_n21389, new_n21390, new_n21391, new_n21392, new_n21393, new_n21394, new_n21395, new_n21396, new_n21397, new_n21398, new_n21399, new_n21400, new_n21401, new_n21402, new_n21403, new_n21404, new_n21405, new_n21406, new_n21407, new_n21408, new_n21409, new_n21410, new_n21411, new_n21412, new_n21413, new_n21414, new_n21415, new_n21416, new_n21417, new_n21418, new_n21419, new_n21420, new_n21421, new_n21422, new_n21423, new_n21424, new_n21425, new_n21426, new_n21427, new_n21428, new_n21429, new_n21430, new_n21431, new_n21432, new_n21433, new_n21434, new_n21435, new_n21436, new_n21437, new_n21438, new_n21439, new_n21440, new_n21441, new_n21442, new_n21443, new_n21444, new_n21445, new_n21446, new_n21447, new_n21448, new_n21449, new_n21450, new_n21451, new_n21452, new_n21453, new_n21454, new_n21455, new_n21456, new_n21457, new_n21458, new_n21459, new_n21460, new_n21461, new_n21462, new_n21463, new_n21464, new_n21465, new_n21466, new_n21467, new_n21468, new_n21469, new_n21470, new_n21471, new_n21472, new_n21473, new_n21474, new_n21475, new_n21476, new_n21477, new_n21478, new_n21479, new_n21480, new_n21481, new_n21482, new_n21483, new_n21484, new_n21485, new_n21486, new_n21487, new_n21488, new_n21489, new_n21490, new_n21491, new_n21492, new_n21493, new_n21494, new_n21495, new_n21496, new_n21497, new_n21498, new_n21499, new_n21500, new_n21501, new_n21502, new_n21503, new_n21504, new_n21505, new_n21506, new_n21507, new_n21508, new_n21509, new_n21510, new_n21511, new_n21512, new_n21513, new_n21514, new_n21515, new_n21516, new_n21517, new_n21518, new_n21519, new_n21520, new_n21521, new_n21522, new_n21523, new_n21524, new_n21525, new_n21526, new_n21527, new_n21528, new_n21529, new_n21530, new_n21531, new_n21532, new_n21533, new_n21534, new_n21535, new_n21536, new_n21537, new_n21538, new_n21539, new_n21540, new_n21541, new_n21542, new_n21543, new_n21544, new_n21545, new_n21546, new_n21547, new_n21548, new_n21549, new_n21550, new_n21551, new_n21552, new_n21553, new_n21554, new_n21555, new_n21556, new_n21557, new_n21558, new_n21559, new_n21560, new_n21561, new_n21562, new_n21563, new_n21564, new_n21565, new_n21566, new_n21567, new_n21568, new_n21569, new_n21570, new_n21571, new_n21572, new_n21573, new_n21574, new_n21575, new_n21576, new_n21577, new_n21578, new_n21579, new_n21580, new_n21581, new_n21582, new_n21583, new_n21584, new_n21585, new_n21586, new_n21587, new_n21588, new_n21589, new_n21590, new_n21591, new_n21592, new_n21593, new_n21594, new_n21595, new_n21596, new_n21597, new_n21598, new_n21599, new_n21600, new_n21601, new_n21602, new_n21603, new_n21604, new_n21605, new_n21606, new_n21607, new_n21608, new_n21609, new_n21610, new_n21611, new_n21612, new_n21613, new_n21614, new_n21615, new_n21616, new_n21617, new_n21618, new_n21619, new_n21620, new_n21621, new_n21622, new_n21623, new_n21624, new_n21625, new_n21626, new_n21627, new_n21628, new_n21629, new_n21630, new_n21631, new_n21632, new_n21633, new_n21634, new_n21635, new_n21636, new_n21637, new_n21638, new_n21639, new_n21640, new_n21641, new_n21642, new_n21643, new_n21644, new_n21645, new_n21646, new_n21647, new_n21648, new_n21649, new_n21650, new_n21651, new_n21652, new_n21653, new_n21654, new_n21655, new_n21656, new_n21657, new_n21658, new_n21659, new_n21660, new_n21661, new_n21662, new_n21663, new_n21664, new_n21665, new_n21666, new_n21667, new_n21668, new_n21669, new_n21670, new_n21671, new_n21672, new_n21673, new_n21674, new_n21675, new_n21676, new_n21677, new_n21678, new_n21679, new_n21680, new_n21681, new_n21682, new_n21683, new_n21684, new_n21685, new_n21686, new_n21687, new_n21688, new_n21689, new_n21690, new_n21691, new_n21692, new_n21693, new_n21694, new_n21695, new_n21696, new_n21697, new_n21698, new_n21699, new_n21700, new_n21701, new_n21702, new_n21703, new_n21704, new_n21705, new_n21706, new_n21707, new_n21708, new_n21709, new_n21710, new_n21711, new_n21712, new_n21713, new_n21714, new_n21715, new_n21716, new_n21717, new_n21718, new_n21719, new_n21720, new_n21721, new_n21722, new_n21723, new_n21724, new_n21725, new_n21726, new_n21727, new_n21728, new_n21729, new_n21730, new_n21731, new_n21732, new_n21733, new_n21734, new_n21735, new_n21736, new_n21737, new_n21738, new_n21739, new_n21740, new_n21741, new_n21742, new_n21743, new_n21744, new_n21745, new_n21746, new_n21747, new_n21748, new_n21749, new_n21750, new_n21751, new_n21752, new_n21753, new_n21754, new_n21755, new_n21756, new_n21757, new_n21758, new_n21759, new_n21760, new_n21761, new_n21762, new_n21763, new_n21764, new_n21765, new_n21766, new_n21767, new_n21768, new_n21769, new_n21770, new_n21771, new_n21772, new_n21773, new_n21774, new_n21775, new_n21776, new_n21777, new_n21778, new_n21779, new_n21780, new_n21781, new_n21782, new_n21783, new_n21784, new_n21785, new_n21786, new_n21787, new_n21788, new_n21789, new_n21790, new_n21791, new_n21792, new_n21793, new_n21794, new_n21795, new_n21796, new_n21797, new_n21798, new_n21799, new_n21800, new_n21801, new_n21802, new_n21803, new_n21804, new_n21805, new_n21806, new_n21807, new_n21808, new_n21809, new_n21810, new_n21811, new_n21812, new_n21813, new_n21814, new_n21815, new_n21816, new_n21817, new_n21818, new_n21819, new_n21820, new_n21821, new_n21822, new_n21823, new_n21824, new_n21825, new_n21826, new_n21827, new_n21828, new_n21829, new_n21830, new_n21831, new_n21832, new_n21833, new_n21834, new_n21835, new_n21836, new_n21837, new_n21838, new_n21839, new_n21840, new_n21841, new_n21842, new_n21843, new_n21844, new_n21845, new_n21846, new_n21847, new_n21848, new_n21849, new_n21850, new_n21851, new_n21852, new_n21853, new_n21854, new_n21855, new_n21856, new_n21857, new_n21858, new_n21859, new_n21860, new_n21861, new_n21862, new_n21863, new_n21864, new_n21865, new_n21866, new_n21867, new_n21868, new_n21869, new_n21870, new_n21871, new_n21872, new_n21873, new_n21874, new_n21875, new_n21876, new_n21877, new_n21878, new_n21879, new_n21880, new_n21881, new_n21882, new_n21883, new_n21884, new_n21885, new_n21886, new_n21887, new_n21888, new_n21889, new_n21890, new_n21891, new_n21892, new_n21893, new_n21894, new_n21895, new_n21896, new_n21897, new_n21898, new_n21899, new_n21900, new_n21901, new_n21902, new_n21903, new_n21904, new_n21905, new_n21906, new_n21907, new_n21908, new_n21909, new_n21910, new_n21911, new_n21912, new_n21913, new_n21914, new_n21915, new_n21916, new_n21917, new_n21918, new_n21919, new_n21920, new_n21921, new_n21922, new_n21923, new_n21924, new_n21925, new_n21926, new_n21927, new_n21928, new_n21929, new_n21930, new_n21931, new_n21932, new_n21933, new_n21934, new_n21935, new_n21936, new_n21937, new_n21938, new_n21939, new_n21940, new_n21941, new_n21942, new_n21943, new_n21944, new_n21945, new_n21946, new_n21947, new_n21948, new_n21949, new_n21950, new_n21951, new_n21952, new_n21953, new_n21954, new_n21955, new_n21956, new_n21957, new_n21958, new_n21959, new_n21960, new_n21961, new_n21962, new_n21963, new_n21964, new_n21965, new_n21966, new_n21967, new_n21968, new_n21969, new_n21970, new_n21971, new_n21972, new_n21973, new_n21974, new_n21975, new_n21976, new_n21977, new_n21978, new_n21979, new_n21980, new_n21981, new_n21982, new_n21983, new_n21984, new_n21985, new_n21986, new_n21987, new_n21988, new_n21989, new_n21990, new_n21991, new_n21992, new_n21993, new_n21994, new_n21995, new_n21996, new_n21997, new_n21998, new_n21999, new_n22000, new_n22001, new_n22002, new_n22003, new_n22004, new_n22005, new_n22006, new_n22007, new_n22008, new_n22009, new_n22010, new_n22011, new_n22012, new_n22013, new_n22014, new_n22015, new_n22016, new_n22017, new_n22018, new_n22019, new_n22020, new_n22021, new_n22022, new_n22023, new_n22024, new_n22025, new_n22026, new_n22027, new_n22028, new_n22029, new_n22030, new_n22031, new_n22032, new_n22033, new_n22034, new_n22035, new_n22036, new_n22037, new_n22038, new_n22039, new_n22040, new_n22041, new_n22042, new_n22043, new_n22044, new_n22045, new_n22046, new_n22047, new_n22048, new_n22049, new_n22050, new_n22051, new_n22052, new_n22053, new_n22054, new_n22055, new_n22056, new_n22057, new_n22058, new_n22059, new_n22060, new_n22061, new_n22062, new_n22063, new_n22064, new_n22065, new_n22066, new_n22067, new_n22068, new_n22069, new_n22070, new_n22071, new_n22072, new_n22073, new_n22074, new_n22075, new_n22076, new_n22077, new_n22078, new_n22079, new_n22080, new_n22081, new_n22082, new_n22083, new_n22084, new_n22085, new_n22086, new_n22087, new_n22088, new_n22089, new_n22090, new_n22091, new_n22092, new_n22093, new_n22094, new_n22095, new_n22096, new_n22097, new_n22098, new_n22099, new_n22100, new_n22101, new_n22102, new_n22103, new_n22104, new_n22105, new_n22106, new_n22107, new_n22108, new_n22109, new_n22110, new_n22111, new_n22112, new_n22113, new_n22114, new_n22115, new_n22116, new_n22117, new_n22118, new_n22119, new_n22120, new_n22121, new_n22122, new_n22123, new_n22124, new_n22125, new_n22126, new_n22127, new_n22128, new_n22129, new_n22130, new_n22131, new_n22132, new_n22133, new_n22134, new_n22135, new_n22136, new_n22137, new_n22138, new_n22139, new_n22140, new_n22141, new_n22142, new_n22143, new_n22144, new_n22145, new_n22146, new_n22147, new_n22148, new_n22149, new_n22150, new_n22151, new_n22152, new_n22153, new_n22154, new_n22155, new_n22156, new_n22157, new_n22158, new_n22159, new_n22160, new_n22161, new_n22162, new_n22163, new_n22164, new_n22165, new_n22166, new_n22167, new_n22168, new_n22169, new_n22170, new_n22171, new_n22172, new_n22173, new_n22174, new_n22175, new_n22176, new_n22177, new_n22178, new_n22179, new_n22180, new_n22181, new_n22182, new_n22183, new_n22184, new_n22185, new_n22186, new_n22187, new_n22188, new_n22189, new_n22190, new_n22191, new_n22192, new_n22193, new_n22194, new_n22195, new_n22196, new_n22197, new_n22198, new_n22199, new_n22200, new_n22201, new_n22202, new_n22203, new_n22204, new_n22205, new_n22206, new_n22207, new_n22208, new_n22209, new_n22210, new_n22211, new_n22212, new_n22213, new_n22214, new_n22215, new_n22216, new_n22217, new_n22218, new_n22219, new_n22220, new_n22221, new_n22222, new_n22223, new_n22224, new_n22225, new_n22226, new_n22227, new_n22228, new_n22229, new_n22230, new_n22231, new_n22232, new_n22233, new_n22234, new_n22235, new_n22236, new_n22237, new_n22238, new_n22239, new_n22240, new_n22241, new_n22242, new_n22243, new_n22244, new_n22245, new_n22246, new_n22247, new_n22248, new_n22249, new_n22250, new_n22251, new_n22252, new_n22253, new_n22254, new_n22255, new_n22256, new_n22257, new_n22258, new_n22259, new_n22260, new_n22261, new_n22262, new_n22263, new_n22264, new_n22265, new_n22266, new_n22267, new_n22268, new_n22269, new_n22270, new_n22271, new_n22272, new_n22273, new_n22274, new_n22275, new_n22276, new_n22277, new_n22278, new_n22279, new_n22280, new_n22281, new_n22282, new_n22283, new_n22284, new_n22285, new_n22286, new_n22287, new_n22288, new_n22289, new_n22290, new_n22291, new_n22292, new_n22293, new_n22294, new_n22295, new_n22296, new_n22297, new_n22298, new_n22299, new_n22300, new_n22301, new_n22302, new_n22303, new_n22304, new_n22305, new_n22306, new_n22307, new_n22308, new_n22309, new_n22310, new_n22311, new_n22312, new_n22313, new_n22314, new_n22315, new_n22316, new_n22317, new_n22318, new_n22319, new_n22320, new_n22321, new_n22322, new_n22323, new_n22324, new_n22325, new_n22326, new_n22327, new_n22328, new_n22329, new_n22330, new_n22331, new_n22332, new_n22333, new_n22334, new_n22335, new_n22336, new_n22337, new_n22338, new_n22339, new_n22340, new_n22341, new_n22342, new_n22343, new_n22344, new_n22345, new_n22346, new_n22347, new_n22348, new_n22349, new_n22350, new_n22351, new_n22352, new_n22353, new_n22354, new_n22355, new_n22356, new_n22357, new_n22358, new_n22359, new_n22360, new_n22361, new_n22362, new_n22363, new_n22364, new_n22365, new_n22366, new_n22367, new_n22368, new_n22369, new_n22370, new_n22371, new_n22372, new_n22373, new_n22374, new_n22375, new_n22376, new_n22377, new_n22378, new_n22379, new_n22380, new_n22381, new_n22382, new_n22383, new_n22384, new_n22385, new_n22386, new_n22387, new_n22388, new_n22389, new_n22390, new_n22391, new_n22392, new_n22393, new_n22394, new_n22395, new_n22396, new_n22397, new_n22398, new_n22399, new_n22400, new_n22401, new_n22402, new_n22403, new_n22404, new_n22405, new_n22406, new_n22407, new_n22408, new_n22409, new_n22410, new_n22411, new_n22412, new_n22413, new_n22414, new_n22415, new_n22416, new_n22417, new_n22418, new_n22419, new_n22420, new_n22421, new_n22422, new_n22423, new_n22424, new_n22425, new_n22426, new_n22427, new_n22428, new_n22429, new_n22430, new_n22431, new_n22432, new_n22433, new_n22434, new_n22435, new_n22436, new_n22437, new_n22438, new_n22439, new_n22440, new_n22441, new_n22442, new_n22443, new_n22444, new_n22445, new_n22446, new_n22447, new_n22448, new_n22449, new_n22450, new_n22451, new_n22452, new_n22453, new_n22454, new_n22455, new_n22456, new_n22457, new_n22458, new_n22459, new_n22460, new_n22461, new_n22462, new_n22463, new_n22464, new_n22465, new_n22466, new_n22467, new_n22468, new_n22469, new_n22470, new_n22471, new_n22472, new_n22473, new_n22474, new_n22475, new_n22476, new_n22477, new_n22478, new_n22479, new_n22480, new_n22481, new_n22482, new_n22483, new_n22484, new_n22485, new_n22486, new_n22487, new_n22488, new_n22489, new_n22490, new_n22491, new_n22492, new_n22493, new_n22494, new_n22495, new_n22496, new_n22497, new_n22498, new_n22499, new_n22500, new_n22501, new_n22502, new_n22503, new_n22504, new_n22505, new_n22506, new_n22507, new_n22508, new_n22509, new_n22510, new_n22511, new_n22512, new_n22513, new_n22514, new_n22515, new_n22516, new_n22517, new_n22518, new_n22519, new_n22520, new_n22521, new_n22522, new_n22523, new_n22524, new_n22525, new_n22526, new_n22527, new_n22528, new_n22529, new_n22530, new_n22531, new_n22532, new_n22533, new_n22534, new_n22535, new_n22536, new_n22537, new_n22538, new_n22539, new_n22540, new_n22541, new_n22542, new_n22543, new_n22544, new_n22545, new_n22546, new_n22547, new_n22548, new_n22549, new_n22550, new_n22551, new_n22552, new_n22553, new_n22554, new_n22555, new_n22556, new_n22557, new_n22558, new_n22559, new_n22560, new_n22561, new_n22562, new_n22563, new_n22564, new_n22565, new_n22566, new_n22567, new_n22568, new_n22569, new_n22570, new_n22571, new_n22572, new_n22573, new_n22574, new_n22575, new_n22576, new_n22577, new_n22578, new_n22579, new_n22580, new_n22581, new_n22582, new_n22583, new_n22584, new_n22585, new_n22586, new_n22587, new_n22588, new_n22589, new_n22590, new_n22591, new_n22592, new_n22593, new_n22594, new_n22595, new_n22596, new_n22597, new_n22598, new_n22599, new_n22600, new_n22601, new_n22602, new_n22603, new_n22604, new_n22605, new_n22606, new_n22607, new_n22608, new_n22609, new_n22610, new_n22611, new_n22612, new_n22613, new_n22614, new_n22615, new_n22616, new_n22617, new_n22618, new_n22619, new_n22620, new_n22621, new_n22622, new_n22623, new_n22624, new_n22625, new_n22626, new_n22627, new_n22628, new_n22629, new_n22630, new_n22631, new_n22632, new_n22633, new_n22634, new_n22635, new_n22636, new_n22637, new_n22638, new_n22639, new_n22640, new_n22641, new_n22642, new_n22643, new_n22644, new_n22645, new_n22646, new_n22647, new_n22648, new_n22649, new_n22650, new_n22651, new_n22652, new_n22653, new_n22654, new_n22655, new_n22656, new_n22657, new_n22658, new_n22659, new_n22660, new_n22661, new_n22662, new_n22663, new_n22664, new_n22665, new_n22666, new_n22667, new_n22668, new_n22669, new_n22670, new_n22671, new_n22672, new_n22673, new_n22674, new_n22675, new_n22676, new_n22677, new_n22678, new_n22679, new_n22680, new_n22681, new_n22682, new_n22683, new_n22684, new_n22685, new_n22686, new_n22687, new_n22688, new_n22689, new_n22690, new_n22691, new_n22692, new_n22693, new_n22694, new_n22695, new_n22696, new_n22697, new_n22698, new_n22699, new_n22700, new_n22701, new_n22702, new_n22703, new_n22704, new_n22705, new_n22706, new_n22707, new_n22708, new_n22709, new_n22710, new_n22711, new_n22712, new_n22713, new_n22714, new_n22715, new_n22716, new_n22717, new_n22718, new_n22719, new_n22720, new_n22721, new_n22722, new_n22723, new_n22724, new_n22725, new_n22726, new_n22727, new_n22728, new_n22729, new_n22730, new_n22731, new_n22732, new_n22733, new_n22734, new_n22735, new_n22736, new_n22737, new_n22738, new_n22739, new_n22740, new_n22741, new_n22742, new_n22743, new_n22744, new_n22745, new_n22746, new_n22747, new_n22748, new_n22749, new_n22750, new_n22751, new_n22752, new_n22753, new_n22754, new_n22755, new_n22756, new_n22757, new_n22758, new_n22759, new_n22760, new_n22761, new_n22762, new_n22763, new_n22764, new_n22765, new_n22766, new_n22767, new_n22768, new_n22769, new_n22770, new_n22771, new_n22772, new_n22773, new_n22774, new_n22775, new_n22776, new_n22777, new_n22778, new_n22779, new_n22780, new_n22781, new_n22782, new_n22783, new_n22784, new_n22785, new_n22786, new_n22787, new_n22788, new_n22789, new_n22790, new_n22791, new_n22792, new_n22793, new_n22794, new_n22795, new_n22796, new_n22797, new_n22798, new_n22799, new_n22800, new_n22801, new_n22802, new_n22803, new_n22804, new_n22805, new_n22806, new_n22807, new_n22808, new_n22809, new_n22810, new_n22811, new_n22812, new_n22813, new_n22814, new_n22815, new_n22816, new_n22817, new_n22818, new_n22819, new_n22820, new_n22821, new_n22822, new_n22823, new_n22824, new_n22825, new_n22826, new_n22827, new_n22828, new_n22829, new_n22830, new_n22831, new_n22832, new_n22833, new_n22834, new_n22835, new_n22836, new_n22837, new_n22838, new_n22839, new_n22840, new_n22841, new_n22842, new_n22843, new_n22844, new_n22845, new_n22846, new_n22847, new_n22848, new_n22849, new_n22850, new_n22851, new_n22852, new_n22853, new_n22854, new_n22855, new_n22856, new_n22857, new_n22858, new_n22859, new_n22860, new_n22861, new_n22862, new_n22863, new_n22864, new_n22865, new_n22866, new_n22867, new_n22868, new_n22869, new_n22870, new_n22871, new_n22872, new_n22873, new_n22874, new_n22875, new_n22876, new_n22877, new_n22878, new_n22879, new_n22880, new_n22881, new_n22882, new_n22883, new_n22884, new_n22885, new_n22886, new_n22887, new_n22888, new_n22889, new_n22890, new_n22891, new_n22892, new_n22893, new_n22894, new_n22895, new_n22896, new_n22897, new_n22898, new_n22899, new_n22900, new_n22901, new_n22902, new_n22903, new_n22904, new_n22905, new_n22906, new_n22907, new_n22908, new_n22909, new_n22910, new_n22911, new_n22912, new_n22913, new_n22914, new_n22915, new_n22916, new_n22917, new_n22918, new_n22919, new_n22920, new_n22921, new_n22922, new_n22923, new_n22924, new_n22925, new_n22926, new_n22927, new_n22928, new_n22929, new_n22930, new_n22931, new_n22932, new_n22933, new_n22934, new_n22935, new_n22936, new_n22937, new_n22938, new_n22939, new_n22940, new_n22941, new_n22942, new_n22943, new_n22944, new_n22945, new_n22946, new_n22947, new_n22948, new_n22949, new_n22950, new_n22951, new_n22952, new_n22953, new_n22954, new_n22955, new_n22956, new_n22957, new_n22958, new_n22959, new_n22960, new_n22961, new_n22962, new_n22963, new_n22964, new_n22965, new_n22966, new_n22967, new_n22968, new_n22969, new_n22970, new_n22971, new_n22972, new_n22973, new_n22974, new_n22975, new_n22976, new_n22977, new_n22978, new_n22979, new_n22980, new_n22981, new_n22982, new_n22983, new_n22984, new_n22985, new_n22986, new_n22987, new_n22988, new_n22989, new_n22990, new_n22991, new_n22992, new_n22993, new_n22994, new_n22995, new_n22996, new_n22997, new_n22998, new_n22999, new_n23000, new_n23001, new_n23002, new_n23003, new_n23004, new_n23005, new_n23006, new_n23007, new_n23008, new_n23009, new_n23010, new_n23011, new_n23012, new_n23013, new_n23014, new_n23015, new_n23016, new_n23017, new_n23018, new_n23019, new_n23020, new_n23021, new_n23022, new_n23023, new_n23024, new_n23025, new_n23026, new_n23027, new_n23028, new_n23029, new_n23030, new_n23031, new_n23032, new_n23033, new_n23034, new_n23035, new_n23036, new_n23037, new_n23038, new_n23039, new_n23040, new_n23041, new_n23042, new_n23043, new_n23044, new_n23045, new_n23046, new_n23047, new_n23048, new_n23049, new_n23050, new_n23051, new_n23052, new_n23053, new_n23054, new_n23055, new_n23056, new_n23057, new_n23058, new_n23059, new_n23060, new_n23061, new_n23062, new_n23063, new_n23064, new_n23065, new_n23066, new_n23067, new_n23068, new_n23069, new_n23070, new_n23071, new_n23072, new_n23073, new_n23074, new_n23075, new_n23076, new_n23077, new_n23078, new_n23079, new_n23080, new_n23081, new_n23082, new_n23083, new_n23084, new_n23085, new_n23086, new_n23087, new_n23088, new_n23089, new_n23090, new_n23091, new_n23092, new_n23093, new_n23094, new_n23095, new_n23096, new_n23097, new_n23098, new_n23099, new_n23100, new_n23101, new_n23102, new_n23103, new_n23104, new_n23105, new_n23106, new_n23107, new_n23108, new_n23109, new_n23110, new_n23111, new_n23112, new_n23113, new_n23114, new_n23115, new_n23116, new_n23117, new_n23118, new_n23119, new_n23120, new_n23121, new_n23122, new_n23123, new_n23124, new_n23125, new_n23126, new_n23127, new_n23128, new_n23129, new_n23130, new_n23131, new_n23132, new_n23133, new_n23134, new_n23135, new_n23136, new_n23137, new_n23138, new_n23139, new_n23140, new_n23141, new_n23142, new_n23143, new_n23144, new_n23145, new_n23146, new_n23147, new_n23148, new_n23149, new_n23150, new_n23151, new_n23152, new_n23153, new_n23154, new_n23155, new_n23156, new_n23157, new_n23158, new_n23159, new_n23160, new_n23161, new_n23162, new_n23163, new_n23164, new_n23165, new_n23166, new_n23167, new_n23168, new_n23169, new_n23170, new_n23171, new_n23172, new_n23173, new_n23174, new_n23175, new_n23176, new_n23177, new_n23178, new_n23179, new_n23180, new_n23181, new_n23182, new_n23183, new_n23184, new_n23185, new_n23186, new_n23187, new_n23188, new_n23189, new_n23190, new_n23191, new_n23192, new_n23193, new_n23194, new_n23195, new_n23196, new_n23197, new_n23198, new_n23199, new_n23200, new_n23201, new_n23202, new_n23203, new_n23204, new_n23205, new_n23206, new_n23207, new_n23208, new_n23209, new_n23210, new_n23211, new_n23212, new_n23213, new_n23214, new_n23215, new_n23216, new_n23217, new_n23218, new_n23219, new_n23220, new_n23221, new_n23222, new_n23223, new_n23224, new_n23225, new_n23226, new_n23227, new_n23228, new_n23229, new_n23230, new_n23231, new_n23232, new_n23233, new_n23234, new_n23235, new_n23236, new_n23237, new_n23238, new_n23239, new_n23240, new_n23241, new_n23242, new_n23243, new_n23244, new_n23245, new_n23246, new_n23247, new_n23248, new_n23249, new_n23250, new_n23251, new_n23252, new_n23253, new_n23254, new_n23255, new_n23256, new_n23257, new_n23258, new_n23259, new_n23260, new_n23261, new_n23262, new_n23263, new_n23264, new_n23265, new_n23266, new_n23267, new_n23268, new_n23269, new_n23270, new_n23271, new_n23272, new_n23273, new_n23274, new_n23275, new_n23276, new_n23277, new_n23278, new_n23279, new_n23280, new_n23281, new_n23282, new_n23283, new_n23284, new_n23285, new_n23286, new_n23287, new_n23288, new_n23289, new_n23290, new_n23291, new_n23292, new_n23293, new_n23294, new_n23295, new_n23296, new_n23297, new_n23298, new_n23299, new_n23300, new_n23301, new_n23302, new_n23303, new_n23304, new_n23305, new_n23306, new_n23307, new_n23308, new_n23309, new_n23310, new_n23311, new_n23312, new_n23313, new_n23314, new_n23315, new_n23316, new_n23317, new_n23318, new_n23319, new_n23320, new_n23321, new_n23322, new_n23323, new_n23324, new_n23325, new_n23326, new_n23327, new_n23328, new_n23329, new_n23330, new_n23331, new_n23332, new_n23333, new_n23334, new_n23335, new_n23336, new_n23337, new_n23338, new_n23339, new_n23340, new_n23341, new_n23342, new_n23343, new_n23344, new_n23345, new_n23346, new_n23347, new_n23348, new_n23349, new_n23350, new_n23351, new_n23352, new_n23353, new_n23354, new_n23355, new_n23356, new_n23357, new_n23358, new_n23359, new_n23360, new_n23361, new_n23362, new_n23363, new_n23364, new_n23365, new_n23366, new_n23367, new_n23368, new_n23369, new_n23370, new_n23371, new_n23372, new_n23373, new_n23374, new_n23375, new_n23376, new_n23377, new_n23378, new_n23379, new_n23380, new_n23381, new_n23382, new_n23383, new_n23384, new_n23385, new_n23386, new_n23387, new_n23388, new_n23389, new_n23390, new_n23391, new_n23392, new_n23393, new_n23394, new_n23395, new_n23396, new_n23397, new_n23398, new_n23399, new_n23400, new_n23401, new_n23402, new_n23403, new_n23404, new_n23405, new_n23406, new_n23407, new_n23408, new_n23409, new_n23410, new_n23411, new_n23412, new_n23413, new_n23414, new_n23415, new_n23416, new_n23417, new_n23418, new_n23419, new_n23420, new_n23421, new_n23422, new_n23423, new_n23424, new_n23425, new_n23426, new_n23427, new_n23428, new_n23429, new_n23430, new_n23431, new_n23432, new_n23433, new_n23434, new_n23435, new_n23436, new_n23437, new_n23438, new_n23439, new_n23440, new_n23441, new_n23442, new_n23443, new_n23444, new_n23445, new_n23446, new_n23447, new_n23448, new_n23449, new_n23450, new_n23451, new_n23452, new_n23453, new_n23454, new_n23455, new_n23456, new_n23457, new_n23458, new_n23459, new_n23460, new_n23461, new_n23462, new_n23463, new_n23464, new_n23465, new_n23466, new_n23467, new_n23468, new_n23469, new_n23470, new_n23471, new_n23472, new_n23473, new_n23474, new_n23475, new_n23476, new_n23477, new_n23478, new_n23479, new_n23480, new_n23481, new_n23482, new_n23483, new_n23484, new_n23485, new_n23486, new_n23487, new_n23488, new_n23489, new_n23490, new_n23491, new_n23492, new_n23493, new_n23494, new_n23495, new_n23496, new_n23497, new_n23498, new_n23499, new_n23500, new_n23501, new_n23502, new_n23503, new_n23504, new_n23505, new_n23506, new_n23507, new_n23508, new_n23509, new_n23510, new_n23511, new_n23512, new_n23513, new_n23514, new_n23515, new_n23516, new_n23517, new_n23518, new_n23519, new_n23520, new_n23521, new_n23522, new_n23523, new_n23524, new_n23525, new_n23526, new_n23527, new_n23528, new_n23529, new_n23530, new_n23531, new_n23532, new_n23533, new_n23534, new_n23535, new_n23536, new_n23537, new_n23538, new_n23539, new_n23540, new_n23541, new_n23542, new_n23543, new_n23544, new_n23545, new_n23546, new_n23547, new_n23548, new_n23549, new_n23550, new_n23551, new_n23552, new_n23553, new_n23554, new_n23555, new_n23556, new_n23557, new_n23558, new_n23559, new_n23560, new_n23561, new_n23562, new_n23563, new_n23564, new_n23565, new_n23566, new_n23567, new_n23568, new_n23569, new_n23570, new_n23571, new_n23572, new_n23573, new_n23574, new_n23575, new_n23576, new_n23577, new_n23578, new_n23579, new_n23580, new_n23581, new_n23582, new_n23583, new_n23584, new_n23585, new_n23586, new_n23587, new_n23588, new_n23589, new_n23590, new_n23591, new_n23592, new_n23593, new_n23594, new_n23595, new_n23596, new_n23597, new_n23598, new_n23599, new_n23600, new_n23601, new_n23602, new_n23603, new_n23604, new_n23605, new_n23606, new_n23607, new_n23608, new_n23609, new_n23610, new_n23611, new_n23612, new_n23613, new_n23614, new_n23615, new_n23616, new_n23617, new_n23618, new_n23619, new_n23620, new_n23621, new_n23622, new_n23623, new_n23624, new_n23625, new_n23626, new_n23627, new_n23628, new_n23629, new_n23630, new_n23631, new_n23632, new_n23633, new_n23634, new_n23635, new_n23636, new_n23637, new_n23638, new_n23639, new_n23640, new_n23641, new_n23642, new_n23643, new_n23644, new_n23645, new_n23646, new_n23647, new_n23648, new_n23649, new_n23650, new_n23651, new_n23652, new_n23653, new_n23654, new_n23655, new_n23656, new_n23657, new_n23658, new_n23659, new_n23660, new_n23661, new_n23662, new_n23663, new_n23664, new_n23665, new_n23666, new_n23667, new_n23668, new_n23669, new_n23670, new_n23671, new_n23672, new_n23673, new_n23674, new_n23675, new_n23676, new_n23677, new_n23678, new_n23679, new_n23680, new_n23681, new_n23682, new_n23683, new_n23684, new_n23685, new_n23686, new_n23687, new_n23688, new_n23689, new_n23690, new_n23691, new_n23692, new_n23693, new_n23694, new_n23695, new_n23696, new_n23697, new_n23698, new_n23699, new_n23700, new_n23701, new_n23702, new_n23703, new_n23704, new_n23705, new_n23706, new_n23707, new_n23708, new_n23709, new_n23710, new_n23711, new_n23712, new_n23713, new_n23714, new_n23715, new_n23716, new_n23717, new_n23718, new_n23719, new_n23720, new_n23721, new_n23722, new_n23723, new_n23724, new_n23725, new_n23726, new_n23727, new_n23728, new_n23729, new_n23730, new_n23731, new_n23732, new_n23733, new_n23734, new_n23735, new_n23736, new_n23737, new_n23738, new_n23739, new_n23740, new_n23741, new_n23742, new_n23743, new_n23744, new_n23745, new_n23746, new_n23747, new_n23748, new_n23749, new_n23750, new_n23751, new_n23752, new_n23753, new_n23754, new_n23755, new_n23756, new_n23757, new_n23758, new_n23759, new_n23760, new_n23761, new_n23762, new_n23763, new_n23764, new_n23765, new_n23766, new_n23767, new_n23768, new_n23769, new_n23770, new_n23771, new_n23772, new_n23773, new_n23774, new_n23775, new_n23776, new_n23777, new_n23778, new_n23779, new_n23780, new_n23781, new_n23782, new_n23783, new_n23784, new_n23785, new_n23786, new_n23787, new_n23788, new_n23789, new_n23790, new_n23791, new_n23792, new_n23793, new_n23794, new_n23795, new_n23796, new_n23797, new_n23798, new_n23799, new_n23800, new_n23801, new_n23802, new_n23803, new_n23804, new_n23805, new_n23806, new_n23807, new_n23808, new_n23809, new_n23810, new_n23811, new_n23812, new_n23813, new_n23814, new_n23815, new_n23816, new_n23817, new_n23818, new_n23819, new_n23820, new_n23821, new_n23822, new_n23823, new_n23824, new_n23825, new_n23826, new_n23827, new_n23828, new_n23829, new_n23830, new_n23831, new_n23832, new_n23833, new_n23834, new_n23835, new_n23836, new_n23837, new_n23838, new_n23839, new_n23840, new_n23841, new_n23842, new_n23843, new_n23844, new_n23845, new_n23846, new_n23847, new_n23848, new_n23849, new_n23850, new_n23851, new_n23852, new_n23853, new_n23854, new_n23855, new_n23856, new_n23857, new_n23858, new_n23859, new_n23860, new_n23861, new_n23862, new_n23863, new_n23864, new_n23865, new_n23866, new_n23867, new_n23868, new_n23869, new_n23870, new_n23871, new_n23872, new_n23873, new_n23874, new_n23875, new_n23876, new_n23877, new_n23878, new_n23879, new_n23880, new_n23881, new_n23882, new_n23883, new_n23884, new_n23885, new_n23886, new_n23887, new_n23888, new_n23889, new_n23890, new_n23891, new_n23892, new_n23893, new_n23894, new_n23895, new_n23896, new_n23897, new_n23898, new_n23899, new_n23900, new_n23901, new_n23902, new_n23903, new_n23904, new_n23905, new_n23906, new_n23907, new_n23908, new_n23909, new_n23910, new_n23911, new_n23912, new_n23913, new_n23914, new_n23915, new_n23916, new_n23917, new_n23918, new_n23919, new_n23920, new_n23921, new_n23922, new_n23923, new_n23924, new_n23925, new_n23926, new_n23927, new_n23928, new_n23929, new_n23930, new_n23931, new_n23932, new_n23933, new_n23934, new_n23935, new_n23936, new_n23937, new_n23938, new_n23939, new_n23940, new_n23941, new_n23942, new_n23943, new_n23944, new_n23945, new_n23946, new_n23947, new_n23948, new_n23949, new_n23950, new_n23951, new_n23952, new_n23953, new_n23954, new_n23955, new_n23956, new_n23957, new_n23958, new_n23959, new_n23960, new_n23961, new_n23962, new_n23963, new_n23964, new_n23965, new_n23966, new_n23967, new_n23968, new_n23969, new_n23970, new_n23971, new_n23972, new_n23973, new_n23974, new_n23975, new_n23976, new_n23977, new_n23978, new_n23979, new_n23980, new_n23981, new_n23982, new_n23983, new_n23984, new_n23985, new_n23986, new_n23987, new_n23988, new_n23989, new_n23990, new_n23991, new_n23992, new_n23993, new_n23994, new_n23995, new_n23996, new_n23997, new_n23998, new_n23999, new_n24000, new_n24001, new_n24002, new_n24003, new_n24004, new_n24005, new_n24006, new_n24007, new_n24008, new_n24009, new_n24010, new_n24011, new_n24012, new_n24013, new_n24014, new_n24015, new_n24016, new_n24017, new_n24018, new_n24019, new_n24020, new_n24021, new_n24022, new_n24023, new_n24024, new_n24025, new_n24026, new_n24027, new_n24028, new_n24029, new_n24030, new_n24031, new_n24032, new_n24033, new_n24034, new_n24035, new_n24036, new_n24037, new_n24038, new_n24039, new_n24040, new_n24041, new_n24042, new_n24043, new_n24044, new_n24045, new_n24046, new_n24047, new_n24048, new_n24049, new_n24050, new_n24051, new_n24052, new_n24053, new_n24054, new_n24055, new_n24056, new_n24057, new_n24058, new_n24059, new_n24060, new_n24061, new_n24062, new_n24063, new_n24064, new_n24065, new_n24066, new_n24067, new_n24068, new_n24069, new_n24070, new_n24071, new_n24072, new_n24073, new_n24074, new_n24075, new_n24076, new_n24077, new_n24078, new_n24079, new_n24080, new_n24081, new_n24082, new_n24083, new_n24084, new_n24085, new_n24086, new_n24087, new_n24088, new_n24089, new_n24090, new_n24091, new_n24092, new_n24093, new_n24094, new_n24095, new_n24096, new_n24097, new_n24098, new_n24099, new_n24100, new_n24101, new_n24102, new_n24103, new_n24104, new_n24105, new_n24106, new_n24107, new_n24108, new_n24109, new_n24110, new_n24111, new_n24112, new_n24113, new_n24114, new_n24115, new_n24116, new_n24117, new_n24118, new_n24119, new_n24120, new_n24121, new_n24122, new_n24123, new_n24124, new_n24125, new_n24126, new_n24127, new_n24128, new_n24129, new_n24130, new_n24131, new_n24132, new_n24133, new_n24134, new_n24135, new_n24136, new_n24137, new_n24138, new_n24139, new_n24140, new_n24141, new_n24142, new_n24143, new_n24144, new_n24145, new_n24146, new_n24147, new_n24148, new_n24149, new_n24150, new_n24151, new_n24152, new_n24153, new_n24154, new_n24155, new_n24156, new_n24157, new_n24158, new_n24159, new_n24160, new_n24161, new_n24162, new_n24163, new_n24164, new_n24165, new_n24166, new_n24167, new_n24168, new_n24169, new_n24170, new_n24171, new_n24172, new_n24173, new_n24174, new_n24175, new_n24176, new_n24177, new_n24178, new_n24179, new_n24180, new_n24181, new_n24182, new_n24183, new_n24184, new_n24185, new_n24186, new_n24187, new_n24188, new_n24189, new_n24190, new_n24191, new_n24192, new_n24193, new_n24194, new_n24195, new_n24196, new_n24197, new_n24198, new_n24199, new_n24200, new_n24201, new_n24202, new_n24203, new_n24204, new_n24205, new_n24206, new_n24207, new_n24208, new_n24209, new_n24210, new_n24211, new_n24212, new_n24213, new_n24214, new_n24215, new_n24216, new_n24217, new_n24218, new_n24219, new_n24220, new_n24221, new_n24222, new_n24223, new_n24224, new_n24225, new_n24226, new_n24227, new_n24228, new_n24229, new_n24230, new_n24231, new_n24232, new_n24233, new_n24234, new_n24235, new_n24236, new_n24237, new_n24238, new_n24239, new_n24240, new_n24241, new_n24242, new_n24243, new_n24244, new_n24245, new_n24246, new_n24247, new_n24248, new_n24249, new_n24250, new_n24251, new_n24252, new_n24253, new_n24254, new_n24255, new_n24256, new_n24257, new_n24258, new_n24259, new_n24260, new_n24261, new_n24262, new_n24263, new_n24264, new_n24265, new_n24266, new_n24267, new_n24268, new_n24269, new_n24270, new_n24271, new_n24272, new_n24273, new_n24274, new_n24275, new_n24276, new_n24277, new_n24278, new_n24279, new_n24280, new_n24281, new_n24282, new_n24283, new_n24284, new_n24285, new_n24286, new_n24287, new_n24288, new_n24289, new_n24290, new_n24291, new_n24292, new_n24293, new_n24294, new_n24295, new_n24296, new_n24297, new_n24298, new_n24299, new_n24300, new_n24301, new_n24302, new_n24303, new_n24304, new_n24305, new_n24306, new_n24307, new_n24308, new_n24309, new_n24310, new_n24311, new_n24312, new_n24313, new_n24314, new_n24315, new_n24316, new_n24317, new_n24318, new_n24319, new_n24320, new_n24321, new_n24322, new_n24323, new_n24324, new_n24325, new_n24326, new_n24327, new_n24328, new_n24329, new_n24330, new_n24331, new_n24332, new_n24333, new_n24334, new_n24335, new_n24336, new_n24337, new_n24338, new_n24339, new_n24340, new_n24341, new_n24342, new_n24343, new_n24344, new_n24345, new_n24346, new_n24347, new_n24348, new_n24349, new_n24350, new_n24351, new_n24352, new_n24353, new_n24354, new_n24355, new_n24356, new_n24357, new_n24358, new_n24359, new_n24360, new_n24361, new_n24362, new_n24363, new_n24364, new_n24365, new_n24366, new_n24367, new_n24368, new_n24369, new_n24370, new_n24371, new_n24372, new_n24373, new_n24374, new_n24375, new_n24376, new_n24377, new_n24378, new_n24379, new_n24380, new_n24381, new_n24382, new_n24383, new_n24384, new_n24385, new_n24386, new_n24387, new_n24388, new_n24389, new_n24390, new_n24391, new_n24392, new_n24393, new_n24394, new_n24395, new_n24396, new_n24397, new_n24398, new_n24399, new_n24400, new_n24401, new_n24402, new_n24403, new_n24404, new_n24405, new_n24406, new_n24407, new_n24408, new_n24409, new_n24410, new_n24411, new_n24412, new_n24413, new_n24414, new_n24415, new_n24416, new_n24417, new_n24418, new_n24419, new_n24420, new_n24421, new_n24422, new_n24423, new_n24424, new_n24425, new_n24426, new_n24427, new_n24428, new_n24429, new_n24430, new_n24431, new_n24432, new_n24433, new_n24434, new_n24435, new_n24436, new_n24437, new_n24438, new_n24439, new_n24440, new_n24441, new_n24442, new_n24443, new_n24444, new_n24445, new_n24446, new_n24447, new_n24448, new_n24449, new_n24450, new_n24451, new_n24452, new_n24453, new_n24454, new_n24455, new_n24456, new_n24457, new_n24458, new_n24459, new_n24460, new_n24461, new_n24462, new_n24463, new_n24464, new_n24465, new_n24466, new_n24467, new_n24468, new_n24469, new_n24470, new_n24471, new_n24472, new_n24473, new_n24474, new_n24475, new_n24476, new_n24477, new_n24478, new_n24479, new_n24480, new_n24481, new_n24482, new_n24483, new_n24484, new_n24485, new_n24486, new_n24487, new_n24488, new_n24489, new_n24490, new_n24491, new_n24492, new_n24493, new_n24494, new_n24495, new_n24496, new_n24497, new_n24498, new_n24499, new_n24500, new_n24501, new_n24502, new_n24503, new_n24504, new_n24505, new_n24506, new_n24507, new_n24508, new_n24509, new_n24510, new_n24511, new_n24512, new_n24513, new_n24514, new_n24515, new_n24516, new_n24517, new_n24518, new_n24519, new_n24520, new_n24521, new_n24522, new_n24523, new_n24524, new_n24525, new_n24526, new_n24527, new_n24528, new_n24529, new_n24530, new_n24531, new_n24532, new_n24533, new_n24534, new_n24535, new_n24536, new_n24537, new_n24538, new_n24539, new_n24540, new_n24541, new_n24542, new_n24543, new_n24544, new_n24545, new_n24546, new_n24547, new_n24548, new_n24549, new_n24550, new_n24551, new_n24552, new_n24553, new_n24554, new_n24555, new_n24556, new_n24557, new_n24558, new_n24559, new_n24560, new_n24561, new_n24562, new_n24563, new_n24564, new_n24565, new_n24566, new_n24567, new_n24568, new_n24569, new_n24570, new_n24571, new_n24572, new_n24573, new_n24574, new_n24575, new_n24576, new_n24577, new_n24578, new_n24579, new_n24580, new_n24581, new_n24582, new_n24583, new_n24584, new_n24585, new_n24586, new_n24587, new_n24588, new_n24589, new_n24590, new_n24591, new_n24592, new_n24593, new_n24594, new_n24595, new_n24596, new_n24597, new_n24598, new_n24599, new_n24600, new_n24601, new_n24602, new_n24603, new_n24604, new_n24605, new_n24606, new_n24607, new_n24608, new_n24609, new_n24610, new_n24611, new_n24612, new_n24613, new_n24614, new_n24615, new_n24616, new_n24617, new_n24618, new_n24619, new_n24620, new_n24621, new_n24622, new_n24623, new_n24624, new_n24625, new_n24626, new_n24627, new_n24628, new_n24629, new_n24630, new_n24631, new_n24632, new_n24633, new_n24634, new_n24635, new_n24636, new_n24637, new_n24638, new_n24639, new_n24640, new_n24641, new_n24642, new_n24643, new_n24644, new_n24645, new_n24646, new_n24647, new_n24648, new_n24649, new_n24650, new_n24651, new_n24652, new_n24653, new_n24654, new_n24655, new_n24656, new_n24657, new_n24658, new_n24659, new_n24660, new_n24661, new_n24662, new_n24663, new_n24664, new_n24665, new_n24666, new_n24667, new_n24668, new_n24669, new_n24670, new_n24671, new_n24672, new_n24673, new_n24674, new_n24675, new_n24676, new_n24677, new_n24678, new_n24679, new_n24680, new_n24681, new_n24682, new_n24683, new_n24684, new_n24685, new_n24686, new_n24687, new_n24688, new_n24689, new_n24690, new_n24691, new_n24692, new_n24693, new_n24694, new_n24695, new_n24696, new_n24697, new_n24698, new_n24699, new_n24700, new_n24701, new_n24702, new_n24703, new_n24704, new_n24705, new_n24706, new_n24707, new_n24708, new_n24709, new_n24710, new_n24711, new_n24712, new_n24713, new_n24714, new_n24715, new_n24716, new_n24717, new_n24718, new_n24719, new_n24720, new_n24721, new_n24722, new_n24723, new_n24724, new_n24725, new_n24726, new_n24727, new_n24728, new_n24729, new_n24730, new_n24731, new_n24732, new_n24733, new_n24734, new_n24735, new_n24736, new_n24737, new_n24738, new_n24739, new_n24740, new_n24741, new_n24742, new_n24743, new_n24744, new_n24745, new_n24746, new_n24747, new_n24748, new_n24749, new_n24750, new_n24751, new_n24752, new_n24753, new_n24754, new_n24755, new_n24756, new_n24757, new_n24758, new_n24759, new_n24760, new_n24761, new_n24762, new_n24763, new_n24764, new_n24765, new_n24766, new_n24767, new_n24768, new_n24769, new_n24770, new_n24771, new_n24772, new_n24773, new_n24774, new_n24775, new_n24776, new_n24777, new_n24778, new_n24779, new_n24780, new_n24781, new_n24782, new_n24783, new_n24784, new_n24785, new_n24786, new_n24787, new_n24788, new_n24789, new_n24790, new_n24791, new_n24792, new_n24793, new_n24794, new_n24795, new_n24796, new_n24797, new_n24798, new_n24799, new_n24800, new_n24801, new_n24802, new_n24803, new_n24804, new_n24805, new_n24806, new_n24807, new_n24808, new_n24809, new_n24810, new_n24811, new_n24812, new_n24813, new_n24814, new_n24815, new_n24816, new_n24817, new_n24818, new_n24819, new_n24820, new_n24821, new_n24822, new_n24823, new_n24824, new_n24825, new_n24826, new_n24827, new_n24828, new_n24829, new_n24830, new_n24831, new_n24832, new_n24833, new_n24834, new_n24835, new_n24836, new_n24837, new_n24838, new_n24839, new_n24840, new_n24841, new_n24842, new_n24843, new_n24844, new_n24845, new_n24846, new_n24847, new_n24848, new_n24849, new_n24850, new_n24851, new_n24852, new_n24853, new_n24854, new_n24855, new_n24856, new_n24857, new_n24858, new_n24859, new_n24860, new_n24861, new_n24862, new_n24863, new_n24864, new_n24865, new_n24866, new_n24867, new_n24868, new_n24869, new_n24870, new_n24871, new_n24872, new_n24873, new_n24874, new_n24875, new_n24876, new_n24877, new_n24878, new_n24879, new_n24880, new_n24881, new_n24882, new_n24883, new_n24884, new_n24885, new_n24886, new_n24887, new_n24888, new_n24889, new_n24890, new_n24891, new_n24892, new_n24893, new_n24894, new_n24895, new_n24896, new_n24897, new_n24898, new_n24899, new_n24900, new_n24901, new_n24902, new_n24903, new_n24904, new_n24905, new_n24906, new_n24907, new_n24908, new_n24909, new_n24910, new_n24911, new_n24912, new_n24913, new_n24914, new_n24915, new_n24916, new_n24917, new_n24918, new_n24919, new_n24920, new_n24921, new_n24922, new_n24923, new_n24924, new_n24925, new_n24926, new_n24927, new_n24928, new_n24929, new_n24930, new_n24931, new_n24932, new_n24933, new_n24934, new_n24935, new_n24936, new_n24937, new_n24938, new_n24939, new_n24940, new_n24941, new_n24942, new_n24943, new_n24944, new_n24945, new_n24946, new_n24947, new_n24948, new_n24949, new_n24950, new_n24951, new_n24952, new_n24953, new_n24954, new_n24955, new_n24956, new_n24957, new_n24958, new_n24959, new_n24960, new_n24961, new_n24962, new_n24963, new_n24964, new_n24965, new_n24966, new_n24967, new_n24968, new_n24969, new_n24970, new_n24971, new_n24972, new_n24973, new_n24974, new_n24975, new_n24976, new_n24977, new_n24978, new_n24979, new_n24980, new_n24981, new_n24982, new_n24983, new_n24984, new_n24985, new_n24986, new_n24987, new_n24988, new_n24989, new_n24990, new_n24991, new_n24992, new_n24993, new_n24994, new_n24995, new_n24996, new_n24997, new_n24998, new_n24999, new_n25000, new_n25001, new_n25002, new_n25003, new_n25004, new_n25005, new_n25006, new_n25007, new_n25008, new_n25009, new_n25010, new_n25011, new_n25012, new_n25013, new_n25014, new_n25015, new_n25016, new_n25017, new_n25018, new_n25019, new_n25020, new_n25021, new_n25022, new_n25023, new_n25024, new_n25025, new_n25026, new_n25027, new_n25028, new_n25029, new_n25030, new_n25031, new_n25032, new_n25033, new_n25034, new_n25035, new_n25036, new_n25037, new_n25038, new_n25039, new_n25040, new_n25041, new_n25042, new_n25043, new_n25044, new_n25045, new_n25046, new_n25047, new_n25048, new_n25049, new_n25050, new_n25051, new_n25052, new_n25053, new_n25054, new_n25055, new_n25056, new_n25057, new_n25058, new_n25059, new_n25060, new_n25061, new_n25062, new_n25063, new_n25064, new_n25065, new_n25066, new_n25067, new_n25068, new_n25069, new_n25070, new_n25071, new_n25072, new_n25073, new_n25074, new_n25075, new_n25076, new_n25077, new_n25078, new_n25079, new_n25080, new_n25081, new_n25082, new_n25083, new_n25084, new_n25085, new_n25086, new_n25087, new_n25088, new_n25089, new_n25090, new_n25091, new_n25092, new_n25093, new_n25094, new_n25095, new_n25096, new_n25097, new_n25098, new_n25099, new_n25100, new_n25101, new_n25102, new_n25103, new_n25104, new_n25105, new_n25106, new_n25107, new_n25108, new_n25109, new_n25110, new_n25111, new_n25112, new_n25113, new_n25114, new_n25115, new_n25116, new_n25117, new_n25118, new_n25119, new_n25120, new_n25121, new_n25122, new_n25123, new_n25124, new_n25125, new_n25126, new_n25127, new_n25128, new_n25129, new_n25130, new_n25131, new_n25132, new_n25133, new_n25134, new_n25135, new_n25136, new_n25137, new_n25138, new_n25139, new_n25140, new_n25141, new_n25142, new_n25143, new_n25144, new_n25145, new_n25146, new_n25147, new_n25148, new_n25149, new_n25150, new_n25151, new_n25152, new_n25153, new_n25154, new_n25155, new_n25156, new_n25157, new_n25158, new_n25159, new_n25160, new_n25161, new_n25162, new_n25163, new_n25164, new_n25165, new_n25166, new_n25167, new_n25168, new_n25169, new_n25170, new_n25171, new_n25172, new_n25173, new_n25174, new_n25175, new_n25176, new_n25177, new_n25178, new_n25179, new_n25180, new_n25181, new_n25182, new_n25183, new_n25184, new_n25185, new_n25186, new_n25187, new_n25188, new_n25189, new_n25190, new_n25191, new_n25192, new_n25193, new_n25194, new_n25195, new_n25196, new_n25197, new_n25198, new_n25199, new_n25200, new_n25201, new_n25202, new_n25203, new_n25204, new_n25205, new_n25206, new_n25207, new_n25208, new_n25209, new_n25210, new_n25211, new_n25212, new_n25213, new_n25214, new_n25215, new_n25216, new_n25217, new_n25218, new_n25219, new_n25220, new_n25221, new_n25222, new_n25223, new_n25224, new_n25225, new_n25226, new_n25227, new_n25228, new_n25229, new_n25230, new_n25231, new_n25232, new_n25233, new_n25234, new_n25235, new_n25236, new_n25237, new_n25238, new_n25239, new_n25240, new_n25241, new_n25242, new_n25243, new_n25244, new_n25245, new_n25246, new_n25247, new_n25248, new_n25249, new_n25250, new_n25251, new_n25252, new_n25253, new_n25254, new_n25255, new_n25256, new_n25257, new_n25258, new_n25259, new_n25260, new_n25261, new_n25262, new_n25263, new_n25264, new_n25265, new_n25266, new_n25267, new_n25268, new_n25269, new_n25270, new_n25271, new_n25272, new_n25273, new_n25274, new_n25275, new_n25276, new_n25277, new_n25278, new_n25279, new_n25280, new_n25281, new_n25282, new_n25283, new_n25284, new_n25285, new_n25286, new_n25287, new_n25288, new_n25289, new_n25290, new_n25291, new_n25292, new_n25293, new_n25294, new_n25295, new_n25296, new_n25297, new_n25298, new_n25299, new_n25300, new_n25301, new_n25302, new_n25303, new_n25304, new_n25305, new_n25306, new_n25307, new_n25308, new_n25309, new_n25310, new_n25311, new_n25312, new_n25313, new_n25314, new_n25315, new_n25316, new_n25317, new_n25318, new_n25319, new_n25320, new_n25321, new_n25322, new_n25323, new_n25324, new_n25325, new_n25326, new_n25327, new_n25328, new_n25329, new_n25330, new_n25331, new_n25332, new_n25333, new_n25334, new_n25335, new_n25336, new_n25337, new_n25338, new_n25339, new_n25340, new_n25341, new_n25342, new_n25343, new_n25344, new_n25345, new_n25346, new_n25347, new_n25348, new_n25349, new_n25350, new_n25351, new_n25352, new_n25353, new_n25354, new_n25355, new_n25356, new_n25357, new_n25358, new_n25359, new_n25360, new_n25361, new_n25362, new_n25363, new_n25364, new_n25365, new_n25366, new_n25367, new_n25368, new_n25369, new_n25370, new_n25371, new_n25372, new_n25373, new_n25374, new_n25375, new_n25376, new_n25377, new_n25378, new_n25379, new_n25380, new_n25381, new_n25382, new_n25383, new_n25384, new_n25385, new_n25386, new_n25387, new_n25388, new_n25389, new_n25390, new_n25391, new_n25392, new_n25393, new_n25394, new_n25395, new_n25396, new_n25397, new_n25398, new_n25399, new_n25400, new_n25401, new_n25402, new_n25403, new_n25404, new_n25405, new_n25406, new_n25407, new_n25408, new_n25409, new_n25410, new_n25411, new_n25412, new_n25413, new_n25414, new_n25415, new_n25416, new_n25417, new_n25418, new_n25419, new_n25420, new_n25421, new_n25422, new_n25423, new_n25424, new_n25425, new_n25426, new_n25427, new_n25428, new_n25429, new_n25430, new_n25431, new_n25432, new_n25433, new_n25434, new_n25435, new_n25436, new_n25437, new_n25438, new_n25439, new_n25440, new_n25441, new_n25442, new_n25443, new_n25444, new_n25445, new_n25446, new_n25447, new_n25448, new_n25449, new_n25450, new_n25451, new_n25452, new_n25453, new_n25454, new_n25455, new_n25456, new_n25457, new_n25458, new_n25459, new_n25460, new_n25461, new_n25462, new_n25463, new_n25464, new_n25465, new_n25466, new_n25467, new_n25468, new_n25469, new_n25470, new_n25471, new_n25472, new_n25473, new_n25474, new_n25475, new_n25476, new_n25477, new_n25478, new_n25479, new_n25480, new_n25481, new_n25482, new_n25483, new_n25484, new_n25485, new_n25486, new_n25487, new_n25488, new_n25489, new_n25490, new_n25491, new_n25492, new_n25493, new_n25494, new_n25495, new_n25496, new_n25497, new_n25498, new_n25499, new_n25500, new_n25501, new_n25502, new_n25503, new_n25504, new_n25505, new_n25506, new_n25507, new_n25508, new_n25509, new_n25510, new_n25511, new_n25512, new_n25513, new_n25514, new_n25515, new_n25516, new_n25517, new_n25518, new_n25519, new_n25520, new_n25521, new_n25522, new_n25523, new_n25524, new_n25525, new_n25526, new_n25527, new_n25528, new_n25529, new_n25530, new_n25531, new_n25532, new_n25533, new_n25534, new_n25535, new_n25536, new_n25537, new_n25538, new_n25539, new_n25540, new_n25541, new_n25542, new_n25543, new_n25544, new_n25545, new_n25546, new_n25547, new_n25548, new_n25549, new_n25550, new_n25551, new_n25552, new_n25553, new_n25554, new_n25555, new_n25556, new_n25557, new_n25558, new_n25559, new_n25560, new_n25561, new_n25562, new_n25563, new_n25564, new_n25565, new_n25566, new_n25567, new_n25568, new_n25569, new_n25570, new_n25571, new_n25572, new_n25573, new_n25574, new_n25575, new_n25576, new_n25577, new_n25578, new_n25579, new_n25580, new_n25581, new_n25582, new_n25583, new_n25584, new_n25585, new_n25586, new_n25587, new_n25588, new_n25589, new_n25590, new_n25591, new_n25592, new_n25593, new_n25594, new_n25595, new_n25596, new_n25597, new_n25598, new_n25599, new_n25600, new_n25601, new_n25602, new_n25603, new_n25604, new_n25605, new_n25606, new_n25607, new_n25608, new_n25609, new_n25610, new_n25611, new_n25612, new_n25613, new_n25614, new_n25615, new_n25616, new_n25617, new_n25618, new_n25619, new_n25620, new_n25621, new_n25622, new_n25623, new_n25624, new_n25625, new_n25626, new_n25627, new_n25628, new_n25629, new_n25630, new_n25631, new_n25632, new_n25633, new_n25634, new_n25635, new_n25636, new_n25637, new_n25638, new_n25639, new_n25640, new_n25641, new_n25642, new_n25643, new_n25644, new_n25645, new_n25646, new_n25647, new_n25648, new_n25649, new_n25650, new_n25651, new_n25652, new_n25653, new_n25654, new_n25655, new_n25656, new_n25657, new_n25658, new_n25659, new_n25660, new_n25661, new_n25662, new_n25663, new_n25664, new_n25665, new_n25666, new_n25667, new_n25668, new_n25669, new_n25670, new_n25671, new_n25672, new_n25673, new_n25674, new_n25675, new_n25676, new_n25677, new_n25678, new_n25679, new_n25680, new_n25681, new_n25682, new_n25683, new_n25684, new_n25685, new_n25686, new_n25687, new_n25688, new_n25689, new_n25690, new_n25691, new_n25692, new_n25693, new_n25694, new_n25695, new_n25696, new_n25697, new_n25698, new_n25699, new_n25700, new_n25701, new_n25702, new_n25703, new_n25704, new_n25705, new_n25706, new_n25707, new_n25708, new_n25709, new_n25710, new_n25711, new_n25712, new_n25713, new_n25714, new_n25715, new_n25716, new_n25717, new_n25718, new_n25719, new_n25720, new_n25721, new_n25722, new_n25723, new_n25724, new_n25725, new_n25726, new_n25727, new_n25728, new_n25729, new_n25730, new_n25731, new_n25732, new_n25733, new_n25734, new_n25735, new_n25736, new_n25737, new_n25738, new_n25739, new_n25740, new_n25741, new_n25742, new_n25743, new_n25744, new_n25745, new_n25746, new_n25747, new_n25748, new_n25749, new_n25750, new_n25751, new_n25752, new_n25753, new_n25754, new_n25755, new_n25756, new_n25757, new_n25758, new_n25759, new_n25760, new_n25761, new_n25762, new_n25763, new_n25764, new_n25765, new_n25766, new_n25767, new_n25768, new_n25769, new_n25770, new_n25771, new_n25772, new_n25773, new_n25774, new_n25775, new_n25776, new_n25777, new_n25778, new_n25779, new_n25780, new_n25781, new_n25782, new_n25783, new_n25784, new_n25785, new_n25786, new_n25787, new_n25788, new_n25789, new_n25790, new_n25791, new_n25792, new_n25793, new_n25794, new_n25795, new_n25796, new_n25797, new_n25798, new_n25799, new_n25800, new_n25801, new_n25802, new_n25803, new_n25804, new_n25805, new_n25806, new_n25807, new_n25808, new_n25809, new_n25810, new_n25811, new_n25812, new_n25813, new_n25814, new_n25815, new_n25816, new_n25817, new_n25818, new_n25819, new_n25820, new_n25821, new_n25822, new_n25823, new_n25824, new_n25825, new_n25826, new_n25827, new_n25828, new_n25829, new_n25830, new_n25831, new_n25832, new_n25833, new_n25834, new_n25835, new_n25836, new_n25837, new_n25838, new_n25839, new_n25840, new_n25841, new_n25842, new_n25843, new_n25844, new_n25845, new_n25846, new_n25847, new_n25848, new_n25849, new_n25850, new_n25851, new_n25852, new_n25853, new_n25854, new_n25855, new_n25856, new_n25857, new_n25858, new_n25859, new_n25860, new_n25861, new_n25862, new_n25863, new_n25864, new_n25865, new_n25866, new_n25867, new_n25868, new_n25869, new_n25870, new_n25871, new_n25872, new_n25873, new_n25874, new_n25875, new_n25876, new_n25877, new_n25878, new_n25879, new_n25880, new_n25881, new_n25882, new_n25883, new_n25884, new_n25885, new_n25886, new_n25887, new_n25888, new_n25889, new_n25890, new_n25891, new_n25892, new_n25893, new_n25894, new_n25895, new_n25896, new_n25897, new_n25898, new_n25899, new_n25900, new_n25901, new_n25902, new_n25903, new_n25904, new_n25905, new_n25906, new_n25907, new_n25908, new_n25909, new_n25910, new_n25911, new_n25912, new_n25913, new_n25914, new_n25915, new_n25916, new_n25917, new_n25918, new_n25919, new_n25920, new_n25921, new_n25922, new_n25923, new_n25924, new_n25925, new_n25926, new_n25927, new_n25928, new_n25929, new_n25930, new_n25931, new_n25932, new_n25933, new_n25934, new_n25935, new_n25936, new_n25937, new_n25938, new_n25939, new_n25940, new_n25941, new_n25942, new_n25943, new_n25944, new_n25945, new_n25946, new_n25947, new_n25948, new_n25949, new_n25950, new_n25951, new_n25952, new_n25953, new_n25954, new_n25955, new_n25956, new_n25957, new_n25958, new_n25959, new_n25960, new_n25961, new_n25962, new_n25963, new_n25964, new_n25965, new_n25966, new_n25967, new_n25968, new_n25969, new_n25970, new_n25971, new_n25972, new_n25973, new_n25974, new_n25975, new_n25976, new_n25977, new_n25978, new_n25979, new_n25980, new_n25981, new_n25982, new_n25983, new_n25984, new_n25985, new_n25986, new_n25987, new_n25988, new_n25989, new_n25990, new_n25991, new_n25992, new_n25993, new_n25994, new_n25995, new_n25996, new_n25997, new_n25998, new_n25999, new_n26000, new_n26001, new_n26002, new_n26003, new_n26004, new_n26005, new_n26006, new_n26007, new_n26008, new_n26009, new_n26010, new_n26011, new_n26012, new_n26013, new_n26014, new_n26015, new_n26016, new_n26017, new_n26018, new_n26019, new_n26020, new_n26021, new_n26022, new_n26023, new_n26024, new_n26025, new_n26026, new_n26027, new_n26028, new_n26029, new_n26030, new_n26031, new_n26032, new_n26033, new_n26034, new_n26035, new_n26036, new_n26037, new_n26038, new_n26039, new_n26040, new_n26041, new_n26042, new_n26043, new_n26044, new_n26045, new_n26046, new_n26047, new_n26048, new_n26049, new_n26050, new_n26051, new_n26052, new_n26053, new_n26054, new_n26055, new_n26056, new_n26057, new_n26058, new_n26059, new_n26060, new_n26061, new_n26062, new_n26063, new_n26064, new_n26065, new_n26066, new_n26067, new_n26068, new_n26069, new_n26070, new_n26071, new_n26072, new_n26073, new_n26074, new_n26075, new_n26076, new_n26077, new_n26078, new_n26079, new_n26080, new_n26081, new_n26082, new_n26083, new_n26084, new_n26085, new_n26086, new_n26087, new_n26088, new_n26089, new_n26090, new_n26091, new_n26092, new_n26093, new_n26094, new_n26095, new_n26096, new_n26097, new_n26098, new_n26099, new_n26100, new_n26101, new_n26102, new_n26103, new_n26104, new_n26105, new_n26106, new_n26107, new_n26108, new_n26109, new_n26110, new_n26111, new_n26112, new_n26113, new_n26114, new_n26115, new_n26116, new_n26117, new_n26118, new_n26119, new_n26120, new_n26121, new_n26122, new_n26123, new_n26124, new_n26125, new_n26126, new_n26127, new_n26128, new_n26129, new_n26130, new_n26131, new_n26132, new_n26133, new_n26134, new_n26135, new_n26136, new_n26137, new_n26138, new_n26139, new_n26140, new_n26141, new_n26142, new_n26143, new_n26144, new_n26145, new_n26146, new_n26147, new_n26148, new_n26149, new_n26150, new_n26151, new_n26152, new_n26153, new_n26154, new_n26155, new_n26156, new_n26157, new_n26158, new_n26159, new_n26160, new_n26161, new_n26162, new_n26163, new_n26164, new_n26165, new_n26166, new_n26167, new_n26168, new_n26169, new_n26170, new_n26171, new_n26172, new_n26173, new_n26174, new_n26175, new_n26176, new_n26177, new_n26178, new_n26179, new_n26180, new_n26181, new_n26182, new_n26183, new_n26184, new_n26185, new_n26186, new_n26187, new_n26188, new_n26189, new_n26190, new_n26191, new_n26192, new_n26193, new_n26194, new_n26195, new_n26196, new_n26197, new_n26198, new_n26199, new_n26200, new_n26201, new_n26202, new_n26203, new_n26204, new_n26205, new_n26206, new_n26207, new_n26208, new_n26209, new_n26210, new_n26211, new_n26212, new_n26213, new_n26214, new_n26215, new_n26216, new_n26217, new_n26218, new_n26219, new_n26220, new_n26221, new_n26222, new_n26223, new_n26224, new_n26225, new_n26226, new_n26227, new_n26228, new_n26229, new_n26230, new_n26231, new_n26232, new_n26233, new_n26234, new_n26235, new_n26236, new_n26237, new_n26238, new_n26239, new_n26240, new_n26241, new_n26242, new_n26243, new_n26244, new_n26245, new_n26246, new_n26247, new_n26248, new_n26249, new_n26250, new_n26251, new_n26252, new_n26253, new_n26254, new_n26255, new_n26256, new_n26257, new_n26258, new_n26259, new_n26260, new_n26261, new_n26262, new_n26263, new_n26264, new_n26265, new_n26266, new_n26267, new_n26268, new_n26269, new_n26270, new_n26271, new_n26272, new_n26273, new_n26274, new_n26275, new_n26276, new_n26277, new_n26278, new_n26279, new_n26280, new_n26281, new_n26282, new_n26283, new_n26284, new_n26285, new_n26286, new_n26287, new_n26288, new_n26289, new_n26290, new_n26291, new_n26292, new_n26293, new_n26294, new_n26295, new_n26296, new_n26297, new_n26298, new_n26299, new_n26300, new_n26301, new_n26302, new_n26303, new_n26304, new_n26305, new_n26306, new_n26307, new_n26308, new_n26309, new_n26310, new_n26311, new_n26312, new_n26313, new_n26314, new_n26315, new_n26316, new_n26317, new_n26318, new_n26319, new_n26320, new_n26321, new_n26322, new_n26323, new_n26324, new_n26325, new_n26326, new_n26327, new_n26328, new_n26329, new_n26330, new_n26331, new_n26332, new_n26333, new_n26334, new_n26335, new_n26336, new_n26337, new_n26338, new_n26339, new_n26340, new_n26341, new_n26342, new_n26343, new_n26344, new_n26345, new_n26346, new_n26347, new_n26348, new_n26349, new_n26350, new_n26351, new_n26352, new_n26353, new_n26354, new_n26355, new_n26356, new_n26357, new_n26358, new_n26359, new_n26360, new_n26361, new_n26362, new_n26363, new_n26364, new_n26365, new_n26366, new_n26367, new_n26368, new_n26369, new_n26370, new_n26371, new_n26372, new_n26373, new_n26374, new_n26375, new_n26376, new_n26377, new_n26378, new_n26379, new_n26380, new_n26381, new_n26382, new_n26383, new_n26384, new_n26385, new_n26386, new_n26387, new_n26388, new_n26389, new_n26390, new_n26391, new_n26392, new_n26393, new_n26394, new_n26395, new_n26396, new_n26397, new_n26398, new_n26399, new_n26400, new_n26401, new_n26402, new_n26403, new_n26404, new_n26405, new_n26406, new_n26407, new_n26408, new_n26409, new_n26410, new_n26411, new_n26412, new_n26413, new_n26414, new_n26415, new_n26416, new_n26417, new_n26418, new_n26419, new_n26420, new_n26421, new_n26422, new_n26423, new_n26424, new_n26425, new_n26426, new_n26427, new_n26428, new_n26429, new_n26430, new_n26431, new_n26432, new_n26433, new_n26434, new_n26435, new_n26436, new_n26437, new_n26438, new_n26439, new_n26440, new_n26441, new_n26442, new_n26443, new_n26444, new_n26445, new_n26446, new_n26447, new_n26448, new_n26449, new_n26450, new_n26451, new_n26452, new_n26453, new_n26454, new_n26455, new_n26456, new_n26457, new_n26458, new_n26459, new_n26460, new_n26461, new_n26462, new_n26463, new_n26464, new_n26465, new_n26466, new_n26467, new_n26468, new_n26469, new_n26470, new_n26471, new_n26472, new_n26473, new_n26474, new_n26475, new_n26476, new_n26477, new_n26478, new_n26479, new_n26480, new_n26481, new_n26482, new_n26483, new_n26484, new_n26485, new_n26486, new_n26487, new_n26488, new_n26489, new_n26490, new_n26491, new_n26492, new_n26493, new_n26494, new_n26495, new_n26496, new_n26497, new_n26498, new_n26499, new_n26500, new_n26501, new_n26502, new_n26503, new_n26504, new_n26505, new_n26506, new_n26507, new_n26508, new_n26509, new_n26510, new_n26511, new_n26512, new_n26513, new_n26514, new_n26515, new_n26516, new_n26517, new_n26518, new_n26519, new_n26520, new_n26521, new_n26522, new_n26523, new_n26524, new_n26525, new_n26526, new_n26527, new_n26528, new_n26529, new_n26530, new_n26531, new_n26532, new_n26533, new_n26534, new_n26535, new_n26536, new_n26537, new_n26538, new_n26539, new_n26540, new_n26541, new_n26542, new_n26543, new_n26544, new_n26545, new_n26546, new_n26547, new_n26548, new_n26549, new_n26550, new_n26551, new_n26552, new_n26553, new_n26554, new_n26555, new_n26556, new_n26557, new_n26558, new_n26559, new_n26560, new_n26561, new_n26562, new_n26563, new_n26564, new_n26565, new_n26566, new_n26567, new_n26568, new_n26569, new_n26570, new_n26571, new_n26572, new_n26573, new_n26574, new_n26575, new_n26576, new_n26577, new_n26578, new_n26579, new_n26580, new_n26581, new_n26582, new_n26583, new_n26584, new_n26585, new_n26586, new_n26587, new_n26588, new_n26589, new_n26590, new_n26591, new_n26592, new_n26593, new_n26594, new_n26595, new_n26596, new_n26597, new_n26598, new_n26599, new_n26600, new_n26601, new_n26602, new_n26603, new_n26604, new_n26605, new_n26606, new_n26607, new_n26608, new_n26609, new_n26610, new_n26611, new_n26612, new_n26613, new_n26614, new_n26615, new_n26616, new_n26617, new_n26618, new_n26619, new_n26620, new_n26621, new_n26622, new_n26623, new_n26624, new_n26625, new_n26626, new_n26627, new_n26628, new_n26629, new_n26630, new_n26631, new_n26632, new_n26633, new_n26634, new_n26635, new_n26636, new_n26637, new_n26638, new_n26639, new_n26640, new_n26641, new_n26642, new_n26643, new_n26644, new_n26645, new_n26646, new_n26647, new_n26648, new_n26649, new_n26650, new_n26651, new_n26652, new_n26653, new_n26654, new_n26655, new_n26656, new_n26657, new_n26658, new_n26659, new_n26660, new_n26661, new_n26662, new_n26663, new_n26664, new_n26665, new_n26666, new_n26667, new_n26668, new_n26669, new_n26670, new_n26671, new_n26672, new_n26673, new_n26674, new_n26675, new_n26676, new_n26677, new_n26678, new_n26679, new_n26680, new_n26681, new_n26682, new_n26683, new_n26684, new_n26685, new_n26686, new_n26687, new_n26688, new_n26689, new_n26690, new_n26691, new_n26692, new_n26693, new_n26694, new_n26695, new_n26696, new_n26697, new_n26698, new_n26699, new_n26700, new_n26701, new_n26702, new_n26703, new_n26704, new_n26705, new_n26706, new_n26707, new_n26708, new_n26709, new_n26710, new_n26711, new_n26712, new_n26713, new_n26714, new_n26715, new_n26716, new_n26717, new_n26718, new_n26719, new_n26720, new_n26721, new_n26722, new_n26723, new_n26724, new_n26725, new_n26726, new_n26727, new_n26728, new_n26729, new_n26730, new_n26731, new_n26732, new_n26733, new_n26734, new_n26735, new_n26736, new_n26737, new_n26738, new_n26739, new_n26740, new_n26741, new_n26742, new_n26743, new_n26744, new_n26745, new_n26746, new_n26747, new_n26748, new_n26749, new_n26750, new_n26751, new_n26752, new_n26753, new_n26754, new_n26755, new_n26756, new_n26757, new_n26758, new_n26759, new_n26760, new_n26761, new_n26762, new_n26763, new_n26764, new_n26765, new_n26766, new_n26767, new_n26768, new_n26769, new_n26770, new_n26771, new_n26772, new_n26773, new_n26774, new_n26775, new_n26776, new_n26777, new_n26778, new_n26779, new_n26780, new_n26781, new_n26782, new_n26783, new_n26784, new_n26785, new_n26786, new_n26787, new_n26788, new_n26789, new_n26790, new_n26791, new_n26792, new_n26793, new_n26794, new_n26795, new_n26796, new_n26797, new_n26798, new_n26799, new_n26800, new_n26801, new_n26802, new_n26803, new_n26804, new_n26805, new_n26806, new_n26807, new_n26808, new_n26809, new_n26810, new_n26811, new_n26812, new_n26813, new_n26814, new_n26815, new_n26816, new_n26817, new_n26818, new_n26819, new_n26820, new_n26821, new_n26822, new_n26823, new_n26824, new_n26825, new_n26826, new_n26827, new_n26828, new_n26829, new_n26830, new_n26831, new_n26832, new_n26833, new_n26834, new_n26835, new_n26836, new_n26837, new_n26838, new_n26839, new_n26840, new_n26841, new_n26842, new_n26843, new_n26844, new_n26845, new_n26846, new_n26847, new_n26848, new_n26849, new_n26850, new_n26851, new_n26852, new_n26853, new_n26854, new_n26855, new_n26856, new_n26857, new_n26858, new_n26859, new_n26860, new_n26861, new_n26862, new_n26863, new_n26864, new_n26865, new_n26866, new_n26867, new_n26868, new_n26869, new_n26870, new_n26871, new_n26872, new_n26873, new_n26874, new_n26875, new_n26876, new_n26877, new_n26878, new_n26879, new_n26880, new_n26881, new_n26882, new_n26883, new_n26884, new_n26885, new_n26886, new_n26887, new_n26888, new_n26889, new_n26890, new_n26891, new_n26892, new_n26893, new_n26894, new_n26895, new_n26896, new_n26897, new_n26898, new_n26899, new_n26900, new_n26901, new_n26902, new_n26903, new_n26904, new_n26905, new_n26906, new_n26907, new_n26908, new_n26909, new_n26910, new_n26911, new_n26912, new_n26913, new_n26914, new_n26915, new_n26916, new_n26917, new_n26918, new_n26919, new_n26920, new_n26921, new_n26922, new_n26923, new_n26924, new_n26925, new_n26926, new_n26927, new_n26928, new_n26929, new_n26930, new_n26931, new_n26932, new_n26933, new_n26934, new_n26935, new_n26936, new_n26937, new_n26938, new_n26939, new_n26940, new_n26941, new_n26942, new_n26943, new_n26944, new_n26945, new_n26946, new_n26947, new_n26948, new_n26949, new_n26950, new_n26951, new_n26952, new_n26953, new_n26954, new_n26955, new_n26956, new_n26957, new_n26958, new_n26959, new_n26960, new_n26961, new_n26962, new_n26963, new_n26964, new_n26965, new_n26966, new_n26967, new_n26968, new_n26969, new_n26970, new_n26971, new_n26972, new_n26973, new_n26974, new_n26975, new_n26976, new_n26977, new_n26978, new_n26979, new_n26980, new_n26981, new_n26982, new_n26983, new_n26984, new_n26985, new_n26986, new_n26987, new_n26988, new_n26989, new_n26990, new_n26991, new_n26992, new_n26993, new_n26994, new_n26995, new_n26996, new_n26997, new_n26998, new_n26999, li0000, li0001, li0002, li0003, li0004, li0005, li0006, li0007, li0008, li0009, li0010, li0011, li0012, li0013, li0014, li0015, li0016, li0017, li0018, li0019, li0020, li0021, li0022, li0023, li0024, li0025, li0026, li0027, li0028, li0029, li0030, li0031, li0032, li0033, li0034, li0035, li0036, li0037, li0038, li0039, li0040, li0041, li0042, li0043, li0044, li0045, li0046, li0047, li0048, li0049, li0050, li0051, li0052, li0053, li0054, li0055, li0056, li0057, li0058, li0059, li0060, li0061, li0062, li0063, li0064, li0065, li0066, li0067, li0068, li0069, li0070, li0071, li0072, li0073, li0074, li0075, li0076, li0077, li0078, li0079, li0080, li0081, li0082, li0083, li0084, li0085, li0086, li0087, li0088, li0089, li0090, li0091, li0092, li0093, li0094, li0095, li0096, li0097, li0098, li0099, li0100, li0101, li0102, li0103, li0104, li0105, li0106, li0107, li0108, li0109, li0110, li0111, li0112, li0113, li0114, li0115, li0116, li0117, li0118, li0119, li0120, li0121, li0122, li0123, li0124, li0125, li0126, li0127, li0128, li0129, li0130, li0131, li0132, li0133, li0134, li0135, li0136, li0137, li0138, li0139, li0140, li0141, li0142, li0143, li0144, li0145, li0146, li0147, li0148, li0149, li0150, li0151, li0152, li0153, li0154, li0155, li0156, li0157, li0158, li0159, li0160, li0161, li0162, li0163, li0164, li0165, li0166, li0167, li0168, li0169, li0170, li0171, li0172, li0173, li0174, li0175, li0176, li0177, li0178, li0179, li0180, li0181, li0182, li0183, li0184, li0185, li0186, li0187, li0188, li0189, li0190, li0191, li0192, li0193, li0194, li0195, li0196, li0197, li0198, li0199, li0200, li0201, li0202, li0203, li0204, li0205, li0206, li0207, li0208, li0209, li0210, li0211, li0212, li0213, li0214, li0215, li0216, li0217, li0218, li0219, li0220, li0221, li0222, li0223, li0224, li0225, li0226, li0227, li0228, li0229, li0230, li0231, li0232, li0233, li0234, li0235, li0236, li0237, li0238, li0239, li0240, li0241, li0242, li0243, li0244, li0245, li0246, li0247, li0248, li0249, li0250, li0251, li0252, li0253, li0254, li0255, li0256, li0257, li0258, li0259, li0260, li0261, li0262, li0263, li0264, li0265, li0266, li0267, li0268, li0269, li0270, li0271, li0272, li0273, li0274, li0275, li0276, li0277, li0278, li0279, li0280, li0281, li0282, li0283, li0284, li0285, li0286, li0287, li0288, li0289, li0290, li0291, li0292, li0293, li0294, li0295, li0296, li0297, li0298, li0299, li0300, li0301, li0302, li0303, li0304, li0305, li0306, li0307, li0308, li0309, li0310, li0311, li0312, li0313, li0314, li0315, li0316, li0317, li0318, li0319, li0320, li0321, li0322, li0323, li0324, li0325, li0326, li0327, li0328, li0329, li0330, li0331, li0332, li0333, li0334, li0335, li0336, li0337, li0338, li0339, li0340, li0341, li0342, li0343, li0344, li0345, li0346, li0347, li0348, li0349, li0350, li0351, li0352, li0353, li0354, li0355, li0356, li0357, li0358, li0359, li0360, li0361, li0362, li0363, li0364, li0365, li0366, li0367, li0368, li0369, li0370, li0371, li0372, li0373, li0374, li0375, li0376, li0377, li0378, li0379, li0380, li0381, li0382, li0383, li0384, li0385, li0386, li0387, li0388, li0389, li0390, li0391, li0392, li0393, li0394, li0395, li0396, li0397, li0398, li0399, li0400, li0401, li0402, li0403, li0404, li0405, li0406, li0407, li0408, li0409, li0410, li0411, li0412, li0413, li0414, li0415, li0416, li0417, li0418, li0419, li0420, li0421, li0422, li0423, li0424, li0425, li0426, li0427, li0428, li0429, li0430, li0431, li0432, li0433, li0434, li0435, li0436, li0437, li0438, li0439, li0440, li0441, li0442, li0443, li0444, li0445, li0446, li0447, li0448, li0449, li0450, li0451, li0452, li0453, li0454, li0455, li0456, li0457, li0458, li0459, li0460, li0461, li0462, li0463, li0464, li0465, li0466, li0467, li0468, li0469, li0470, li0471, li0472, li0473, li0474, li0475, li0476, li0477, li0478, li0479, li0480, li0481, li0482, li0483, li0484, li0485, li0486, li0487, li0488, li0489, li0490, li0491, li0492, li0493, li0494, li0495, li0496, li0497, li0498, li0499, li0500, li0501, li0502, li0503, li0504, li0505, li0506, li0507, li0508, li0509, li0510, li0511, li0512, li0513, li0514, li0515, li0516, li0517, li0518, li0519, li0520, li0521, li0522, li0523, li0524, li0525, li0526, li0527, li0528, li0529, li0530, li0531, li0532, li0533, li0534, li0535, li0536, li0537, li0538, li0539, li0540, li0541, li0542, li0543, li0544, li0545, li0546, li0547, li0548, li0549, li0550, li0551, li0552, li0553, li0554, li0555, li0556, li0557, li0558, li0559, li0560, li0561, li0562, li0563, li0564, li0565, li0566, li0567, li0568, li0569, li0570, li0571, li0572, li0573, li0574, li0575, li0576, li0577, li0578, li0579, li0580, li0581, li0582, li0583, li0584, li0585, li0586, li0587, li0588, li0589, li0590, li0591, li0592, li0593, li0594, li0595, li0596, li0597, li0598, li0599, li0600, li0601, li0602, li0603, li0604, li0605, li0606, li0607, li0608, li0609, li0610, li0611, li0612, li0613, li0614, li0615, li0616, li0617, li0618, li0619, li0620, li0621, li0622, li0623, li0624, li0625, li0626, li0627, li0628, li0629, li0630, li0631, li0632, li0633, li0634, li0635, li0636, li0637, li0638, li0639, li0640, li0641, li0642, li0643, li0644, li0645, li0646, li0647, li0648, li0649, li0650, li0651, li0652, li0653, li0654, li0655, li0656, li0657, li0658, li0659, li0660, li0661, li0662, li0663, li0664, li0665, li0666, li0667, li0668, li0669, li0670, li0671, li0672, li0673, li0674, li0675, li0676, li0677, li0678, li0679, li0680, li0681, li0682, li0683, li0684, li0685, li0686, li0687, li0688, li0689, li0690, li0691, li0692, li0693, li0694, li0695, li0696, li0697, li0698, li0699, li0700, li0701, li0702, li0703, li0704, li0705, li0706, li0707, li0708, li0709, li0710, li0711, li0712, li0713, li0714, li0715, li0716, li0717, li0718, li0719, li0720, li0721, li0722, li0723, li0724, li0725, li0726, li0727, li0728, li0729, li0730, li0731, li0732, li0733, li0734, li0735, li0736, li0737, li0738, li0739, li0740, li0741, li0742, li0743, li0744, li0745, li0746, li0747, li0748, li0749, li0750, li0751, li0752, li0753, li0754, li0755, li0756, li0757, li0758, li0759, li0760, li0761, li0762, li0763, li0764, li0765, li0766, li0767, li0768, li0769, li0770, li0771, li0772, li0773, li0774, li0775, li0776, li0777, li0778, li0779, li0780, li0781, li0782, li0783, li0784, li0785, li0786, li0787, li0788, li0789, li0790, li0791, li0792, li0793, li0794, li0795, li0796, li0797, li0798, li0799, li0800, li0801, li0802, li0803, li0804, li0805, li0806, li0807, li0808, li0809, li0810, li0811, li0812, li0813, li0814, li0815, li0816, li0817, li0818, li0819, li0820, li0821, li0822, li0823, li0824, li0825, li0826, li0827, li0828, li0829, li0830, li0831, li0832, li0833, li0834, li0835, li0836, li0837, li0838, li0839, li0840, li0841, li0842, li0843, li0844, li0845, li0846, li0847, li0848, li0849, li0850, li0851, li0852, li0853, li0854, li0855, li0856, li0857, li0858, li0859, li0860, li0861, li0862, li0863, li0864, li0865, li0866, li0867, li0868, li0869, li0870, li0871, li0872, li0873, li0874, li0875, li0876, li0877, li0878, li0879, li0880, li0881, li0882, li0883, li0884, li0885, li0886, li0887, li0888, li0889, li0890, li0891, li0892, li0893, li0894, li0895, li0896, li0897, li0898, li0899, li0900, li0901, li0902, li0903, li0904, li0905, li0906, li0907, li0908, li0909, li0910, li0911, li0912, li0913, li0914, li0915, li0916, li0917, li0918, li0919, li0920, li0921, li0922, li0923, li0924, li0925, li0926, li0927, li0928, li0929, li0930, li0931, li0932, li0933, li0934, li0935, li0936, li0937, li0938, li0939, li0940, li0941, li0942, li0943, li0944, li0945, li0946, li0947, li0948, li0949, li0950, li0951, li0952, li0953, li0954, li0955, li0956, li0957, li0958, li0959, li0960, li0961, li0962, li0963, li0964, li0965, li0966, li0967, li0968, li0969, li0970, li0971, li0972, li0973, li0974, li0975, li0976, li0977, li0978, li0979, li0980, li0981, li0982, li0983, li0984, li0985, li0986, li0987, li0988, li0989, li0990, li0991, li0992, li0993, li0994, li0995, li0996, li0997, li0998, li0999, li1000, li1001, li1002, li1003, li1004, li1005, li1006, li1007, li1008, li1009, li1010, li1011, li1012, li1013, li1014, li1015, li1016, li1017, li1018, li1019, li1020, li1021, li1022, li1023, li1024, li1025, li1026, li1027, li1028, li1029, li1030, li1031, li1032, li1033, li1034, li1035, li1036, li1037, li1038, li1039, li1040, li1041, li1042, li1043, li1044, li1045, li1046, li1047, li1048, li1049, li1050, li1051, li1052, li1053, li1054, li1055, li1056, li1057, li1058, li1059, li1060, li1061, li1062, li1063, li1064, li1065, li1066, li1067, li1068, li1069, li1070, li1071, li1072, li1073, li1074, li1075, li1076, li1077, li1078, li1079, li1080, li1081, li1082, li1083, li1084, li1085, li1086, li1087, li1088, li1089, li1090, li1091, li1092, li1093, li1094, li1095, li1096, li1097, li1098, li1099, li1100, li1101, li1102, li1103, li1104, li1105, li1106, li1107, li1108, li1109, li1110, li1111, li1112, li1113, li1114, li1115, li1116, li1117, li1118, li1119, li1120, li1121, li1122, li1123, li1124, li1125, li1126, li1127, li1128, li1129, li1130, li1131, li1132, li1133, li1134, li1135, li1136, li1137, li1138, li1139, li1140, li1141, li1142, li1143, li1144, li1145, li1146, li1147, li1148, li1149, li1150, li1151, li1152, li1153, li1154, li1155, li1156, li1157, li1158, li1159, li1160, li1161, li1162, li1163, li1164, li1165, li1166, li1167, li1168, li1169, li1170, li1171, li1172, li1173, li1174, li1175, li1176, li1177, li1178, li1179, li1180, li1181, li1182, li1183, li1184, li1185, li1186, li1187, li1188, li1189, li1190, li1191, li1192, li1193, li1194, li1195, li1196, li1197, li1198, li1199, li1200, li1201, li1202, li1203, li1204, li1205, li1206, li1207, li1208, li1209, li1210, li1211, li1212, li1213, li1214, li1215, li1216, li1217, li1218, li1219, li1220, li1221, li1222, li1223, li1224, li1225, li1226, li1227, li1228, li1229, li1230, li1231, li1232, li1233, li1234, li1235, li1236, li1237, li1238, li1239, li1240, li1241, li1242, li1243, li1244, li1245, li1246, li1247, li1248, li1249, li1250, li1251, li1252, li1253, li1254, li1255, li1256, li1257, li1258, li1259, li1260, li1261, li1262, li1263, li1264, li1265, li1266, li1267, li1268, li1269, li1270, li1271, li1272, li1273, li1274, li1275, li1276, li1277, li1278, li1279, li1280, li1281, li1282, li1283, li1284, li1285, li1286, li1287, li1288, li1289, li1290, li1291, li1292, li1293, li1294, li1295, li1296, li1297, li1298, li1299, li1300, li1301, li1302, li1303, li1304, li1305, li1306, li1307, li1308, li1309, li1310, li1311, li1312, li1313, li1314, li1315, li1316, li1317, li1318, li1319, li1320, li1321, li1322, li1323, li1324, li1325, li1326, li1327, li1328, li1329, li1330, li1331, li1332, li1333, li1334, li1335, li1336, li1337, li1338, li1339, li1340, li1341, li1342, li1343, li1344, li1345, li1346, li1347, li1348, li1349, li1350, li1351, li1352, li1353, li1354, li1355, li1356, li1357, li1358, li1359, li1360, li1361, li1362, li1363, li1364, li1365, li1366, li1367, li1368, li1369, li1370, li1371, li1372, li1373, li1374, li1375, li1376, li1377, li1378, li1379, li1380, li1381, li1382, li1383, li1384, li1385, li1386, li1387, li1388, li1389, li1390, li1391, li1392, li1393, li1394, li1395, li1396, li1397, li1398, li1399, li1400, li1401, li1402, li1403, li1404, li1405, li1406, li1407, li1408, li1409, li1410, li1411, li1412, li1413, li1414, li1415, li1416, li1417, li1418, li1419, li1420, li1421, li1422, li1423, li1424, li1425, li1426, li1427, li1428, li1429, li1430, li1431, li1432, li1433, li1434, li1435, li1436, li1437, li1438, li1439, li1440, li1441, li1442, li1443, li1444, li1445, li1446, li1447, li1448, li1449, li1450, li1451, li1452, li1453, li1454, li1455, li1456, li1457, li1458, li1459, li1460, li1461, li1462, li1463, li1464, li1465, li1466, li1467, li1468, li1469, li1470, li1471, li1472, li1473, li1474, li1475, li1476;
  assign new_n1942 = lo0044 & lo0046 ;
  assign new_n1943 = ~lo0041 & ~lo0042 ;
  assign new_n1944 = ~lo0039 & ~lo0040 ;
  assign new_n1945 = ~lo0037 & ~lo0038 ;
  assign new_n1946 = new_n1944 & new_n1945 ;
  assign new_n1947 = new_n1943 & new_n1946 ;
  assign new_n1948 = lo0031 & lo0032 ;
  assign new_n1949 = lo0029 & lo0030 ;
  assign new_n1950 = new_n1948 & new_n1949 ;
  assign new_n1951 = lo0035 & lo0036 ;
  assign new_n1952 = ~lo0033 & ~lo0034 ;
  assign new_n1953 = new_n1951 & new_n1952 ;
  assign new_n1954 = new_n1950 & new_n1953 ;
  assign new_n1955 = ~lo0021 & ~lo0024 ;
  assign new_n1956 = lo0022 & lo0023 ;
  assign new_n1957 = new_n1955 & new_n1956 ;
  assign new_n1958 = lo0027 & ~lo0028 ;
  assign new_n1959 = lo0025 & ~lo0026 ;
  assign new_n1960 = new_n1958 & new_n1959 ;
  assign new_n1961 = new_n1957 & new_n1960 ;
  assign new_n1962 = new_n1954 & new_n1961 ;
  assign new_n1963 = new_n1947 & new_n1962 ;
  assign new_n1964 = ~lo0019 & lo0020 ;
  assign new_n1965 = new_n1963 & new_n1964 ;
  assign new_n1966 = ~lo0020 & new_n1963 ;
  assign new_n1967 = ~lo0019 & new_n1966 ;
  assign new_n1968 = lo0019 & new_n1966 ;
  assign new_n1969 = lo0018 & ~new_n1968 ;
  assign new_n1970 = ~new_n1967 & new_n1969 ;
  assign new_n1971 = ~new_n1965 & new_n1970 ;
  assign new_n1972 = lo0021 & new_n1971 ;
  assign new_n1973 = new_n1943 & new_n1972 ;
  assign new_n1974 = new_n1942 & new_n1973 ;
  assign new_n1975 = lo0041 & ~lo0042 ;
  assign new_n1976 = new_n1972 & new_n1975 ;
  assign new_n1977 = new_n1942 & new_n1976 ;
  assign new_n1978 = ~lo0021 & new_n1971 ;
  assign new_n1979 = new_n1943 & new_n1978 ;
  assign new_n1980 = new_n1942 & new_n1979 ;
  assign new_n1981 = lo0041 & lo0042 ;
  assign new_n1982 = new_n1978 & new_n1981 ;
  assign new_n1983 = new_n1942 & new_n1982 ;
  assign new_n1984 = ~lo0041 & lo0042 ;
  assign new_n1985 = new_n1972 & new_n1984 ;
  assign new_n1986 = new_n1942 & new_n1985 ;
  assign new_n1987 = new_n1978 & new_n1984 ;
  assign new_n1988 = new_n1942 & new_n1987 ;
  assign new_n1989 = new_n1975 & new_n1978 ;
  assign new_n1990 = new_n1942 & new_n1989 ;
  assign new_n1991 = new_n1972 & new_n1981 ;
  assign new_n1992 = new_n1942 & new_n1991 ;
  assign new_n1993 = lo0043 & lo0044 ;
  assign new_n1994 = new_n1973 & new_n1993 ;
  assign new_n1995 = new_n1979 & new_n1993 ;
  assign new_n1996 = new_n1987 & new_n1993 ;
  assign new_n1997 = new_n1989 & new_n1993 ;
  assign new_n1998 = new_n1985 & new_n1993 ;
  assign new_n1999 = new_n1976 & new_n1993 ;
  assign new_n2000 = new_n1982 & new_n1993 ;
  assign new_n2001 = new_n1991 & new_n1993 ;
  assign new_n2002 = lo0044 & lo1051 ;
  assign new_n2003 = new_n1987 & new_n2002 ;
  assign new_n2004 = new_n1989 & new_n2002 ;
  assign new_n2005 = new_n1976 & new_n2002 ;
  assign new_n2006 = new_n1979 & new_n2002 ;
  assign new_n2007 = new_n1982 & new_n2002 ;
  assign new_n2008 = new_n1985 & new_n2002 ;
  assign new_n2009 = new_n1973 & new_n2002 ;
  assign new_n2010 = new_n1991 & new_n2002 ;
  assign new_n2011 = lo0044 & lo0045 ;
  assign new_n2012 = new_n1987 & new_n2011 ;
  assign new_n2013 = new_n1991 & new_n2011 ;
  assign new_n2014 = new_n1989 & new_n2011 ;
  assign new_n2015 = new_n1973 & new_n2011 ;
  assign new_n2016 = new_n1976 & new_n2011 ;
  assign new_n2017 = new_n1979 & new_n2011 ;
  assign new_n2018 = new_n1982 & new_n2011 ;
  assign new_n2019 = new_n1985 & new_n2011 ;
  assign new_n2020 = ~lo0890 & ~lo0891 ;
  assign new_n2021 = ~lo0936 & ~lo0937 ;
  assign new_n2022 = new_n2020 & new_n2021 ;
  assign new_n2023 = lo1127 & ~new_n2022 ;
  assign new_n2024 = lo1128 & new_n2022 ;
  assign new_n2025 = ~new_n2023 & ~new_n2024 ;
  assign new_n2026 = lo1146 & ~new_n2022 ;
  assign new_n2027 = lo1147 & new_n2022 ;
  assign new_n2028 = ~new_n2026 & ~new_n2027 ;
  assign new_n2029 = lo1148 & ~new_n2022 ;
  assign new_n2030 = lo1149 & new_n2022 ;
  assign new_n2031 = ~new_n2029 & ~new_n2030 ;
  assign new_n2032 = lo1150 & ~new_n2022 ;
  assign new_n2033 = lo1151 & new_n2022 ;
  assign new_n2034 = ~new_n2032 & ~new_n2033 ;
  assign new_n2035 = lo1152 & ~new_n2022 ;
  assign new_n2036 = lo1153 & new_n2022 ;
  assign new_n2037 = ~new_n2035 & ~new_n2036 ;
  assign new_n2038 = lo1154 & ~new_n2022 ;
  assign new_n2039 = lo1155 & new_n2022 ;
  assign new_n2040 = ~new_n2038 & ~new_n2039 ;
  assign new_n2041 = lo1156 & ~new_n2022 ;
  assign new_n2042 = lo1157 & new_n2022 ;
  assign new_n2043 = ~new_n2041 & ~new_n2042 ;
  assign new_n2044 = lo1158 & ~new_n2022 ;
  assign new_n2045 = lo1159 & new_n2022 ;
  assign new_n2046 = ~new_n2044 & ~new_n2045 ;
  assign new_n2047 = lo1160 & ~new_n2022 ;
  assign new_n2048 = lo1161 & new_n2022 ;
  assign new_n2049 = ~new_n2047 & ~new_n2048 ;
  assign new_n2050 = lo1162 & ~new_n2022 ;
  assign new_n2051 = lo1163 & new_n2022 ;
  assign new_n2052 = ~new_n2050 & ~new_n2051 ;
  assign new_n2053 = lo1164 & ~new_n2022 ;
  assign new_n2054 = lo1165 & new_n2022 ;
  assign new_n2055 = ~new_n2053 & ~new_n2054 ;
  assign new_n2056 = lo1166 & ~new_n2022 ;
  assign new_n2057 = lo1167 & new_n2022 ;
  assign new_n2058 = ~new_n2056 & ~new_n2057 ;
  assign new_n2059 = lo1168 & ~new_n2022 ;
  assign new_n2060 = lo1169 & new_n2022 ;
  assign new_n2061 = ~new_n2059 & ~new_n2060 ;
  assign new_n2062 = lo1170 & ~new_n2022 ;
  assign new_n2063 = lo1171 & new_n2022 ;
  assign new_n2064 = ~new_n2062 & ~new_n2063 ;
  assign new_n2065 = lo1172 & ~new_n2022 ;
  assign new_n2066 = lo1173 & new_n2022 ;
  assign new_n2067 = ~new_n2065 & ~new_n2066 ;
  assign new_n2068 = ~lo0939 & ~lo0941 ;
  assign new_n2069 = ~lo0940 & new_n2068 ;
  assign new_n2070 = ~lo0886 & lo0938 ;
  assign new_n2071 = new_n2069 & new_n2070 ;
  assign new_n2072 = lo1124 & ~new_n2022 ;
  assign new_n2073 = lo1125 & new_n2022 ;
  assign new_n2074 = ~new_n2072 & ~new_n2073 ;
  assign new_n2075 = new_n2071 & ~new_n2074 ;
  assign new_n2076 = lo1120 & ~new_n2022 ;
  assign new_n2077 = lo1121 & new_n2022 ;
  assign new_n2078 = ~new_n2076 & ~new_n2077 ;
  assign new_n2079 = new_n2071 & ~new_n2078 ;
  assign new_n2080 = lo1174 & ~new_n2022 ;
  assign new_n2081 = lo1175 & new_n2022 ;
  assign new_n2082 = ~new_n2080 & ~new_n2081 ;
  assign new_n2083 = new_n2071 & ~new_n2082 ;
  assign new_n2084 = lo1176 & ~new_n2022 ;
  assign new_n2085 = lo1177 & new_n2022 ;
  assign new_n2086 = ~new_n2084 & ~new_n2085 ;
  assign new_n2087 = new_n2071 & ~new_n2086 ;
  assign new_n2088 = lo1178 & ~new_n2022 ;
  assign new_n2089 = lo1179 & new_n2022 ;
  assign new_n2090 = ~new_n2088 & ~new_n2089 ;
  assign new_n2091 = new_n2071 & ~new_n2090 ;
  assign new_n2092 = lo1180 & ~new_n2022 ;
  assign new_n2093 = lo1181 & new_n2022 ;
  assign new_n2094 = ~new_n2092 & ~new_n2093 ;
  assign new_n2095 = new_n2071 & ~new_n2094 ;
  assign new_n2096 = lo1182 & ~new_n2022 ;
  assign new_n2097 = lo1183 & new_n2022 ;
  assign new_n2098 = ~new_n2096 & ~new_n2097 ;
  assign new_n2099 = new_n2071 & ~new_n2098 ;
  assign new_n2100 = lo1184 & ~new_n2022 ;
  assign new_n2101 = lo1185 & new_n2022 ;
  assign new_n2102 = ~new_n2100 & ~new_n2101 ;
  assign new_n2103 = new_n2071 & ~new_n2102 ;
  assign new_n2104 = lo1186 & ~new_n2022 ;
  assign new_n2105 = lo1187 & new_n2022 ;
  assign new_n2106 = ~new_n2104 & ~new_n2105 ;
  assign new_n2107 = new_n2071 & ~new_n2106 ;
  assign new_n2108 = lo1188 & ~new_n2022 ;
  assign new_n2109 = lo1189 & new_n2022 ;
  assign new_n2110 = ~new_n2108 & ~new_n2109 ;
  assign new_n2111 = new_n2071 & ~new_n2110 ;
  assign new_n2112 = lo1190 & ~new_n2022 ;
  assign new_n2113 = lo1191 & new_n2022 ;
  assign new_n2114 = ~new_n2112 & ~new_n2113 ;
  assign new_n2115 = new_n2071 & ~new_n2114 ;
  assign new_n2116 = lo1192 & ~new_n2022 ;
  assign new_n2117 = lo1193 & new_n2022 ;
  assign new_n2118 = ~new_n2116 & ~new_n2117 ;
  assign new_n2119 = new_n2071 & ~new_n2118 ;
  assign new_n2120 = lo1194 & ~new_n2022 ;
  assign new_n2121 = lo1195 & new_n2022 ;
  assign new_n2122 = ~new_n2120 & ~new_n2121 ;
  assign new_n2123 = new_n2071 & ~new_n2122 ;
  assign new_n2124 = lo1196 & ~new_n2022 ;
  assign new_n2125 = lo1197 & new_n2022 ;
  assign new_n2126 = ~new_n2124 & ~new_n2125 ;
  assign new_n2127 = new_n2071 & ~new_n2126 ;
  assign new_n2128 = lo1198 & ~new_n2022 ;
  assign new_n2129 = lo1199 & new_n2022 ;
  assign new_n2130 = ~new_n2128 & ~new_n2129 ;
  assign new_n2131 = new_n2071 & ~new_n2130 ;
  assign new_n2132 = lo1200 & ~new_n2022 ;
  assign new_n2133 = lo1201 & new_n2022 ;
  assign new_n2134 = ~new_n2132 & ~new_n2133 ;
  assign new_n2135 = new_n2071 & ~new_n2134 ;
  assign new_n2136 = ~lo0934 & ~lo0935 ;
  assign new_n2137 = ~lo0933 & new_n2136 ;
  assign new_n2138 = new_n2021 & new_n2137 ;
  assign new_n2139 = new_n2071 & ~new_n2138 ;
  assign new_n2140 = lo1126 & ~new_n2139 ;
  assign new_n2141 = lo1122 & new_n2139 ;
  assign new_n2142 = ~new_n2140 & ~new_n2141 ;
  assign new_n2143 = lo1202 & ~new_n2139 ;
  assign new_n2144 = lo1203 & new_n2139 ;
  assign new_n2145 = ~new_n2143 & ~new_n2144 ;
  assign new_n2146 = lo1204 & ~new_n2139 ;
  assign new_n2147 = lo1205 & new_n2139 ;
  assign new_n2148 = ~new_n2146 & ~new_n2147 ;
  assign new_n2149 = lo1206 & ~new_n2139 ;
  assign new_n2150 = lo1207 & new_n2139 ;
  assign new_n2151 = ~new_n2149 & ~new_n2150 ;
  assign new_n2152 = lo1208 & ~new_n2139 ;
  assign new_n2153 = lo1209 & new_n2139 ;
  assign new_n2154 = ~new_n2152 & ~new_n2153 ;
  assign new_n2155 = lo1210 & ~new_n2139 ;
  assign new_n2156 = lo1211 & new_n2139 ;
  assign new_n2157 = ~new_n2155 & ~new_n2156 ;
  assign new_n2158 = lo1212 & ~new_n2139 ;
  assign new_n2159 = lo1213 & new_n2139 ;
  assign new_n2160 = ~new_n2158 & ~new_n2159 ;
  assign new_n2161 = lo1214 & ~new_n2139 ;
  assign new_n2162 = lo1215 & new_n2139 ;
  assign new_n2163 = ~new_n2161 & ~new_n2162 ;
  assign new_n2164 = lo1216 & ~new_n2139 ;
  assign new_n2165 = lo1217 & new_n2139 ;
  assign new_n2166 = ~new_n2164 & ~new_n2165 ;
  assign new_n2167 = lo1218 & ~new_n2139 ;
  assign new_n2168 = lo1219 & new_n2139 ;
  assign new_n2169 = ~new_n2167 & ~new_n2168 ;
  assign new_n2170 = lo1220 & ~new_n2139 ;
  assign new_n2171 = lo1221 & new_n2139 ;
  assign new_n2172 = ~new_n2170 & ~new_n2171 ;
  assign new_n2173 = lo1222 & ~new_n2139 ;
  assign new_n2174 = lo1223 & new_n2139 ;
  assign new_n2175 = ~new_n2173 & ~new_n2174 ;
  assign new_n2176 = lo1224 & ~new_n2139 ;
  assign new_n2177 = lo1225 & new_n2139 ;
  assign new_n2178 = ~new_n2176 & ~new_n2177 ;
  assign new_n2179 = lo1226 & ~new_n2139 ;
  assign new_n2180 = lo1227 & new_n2139 ;
  assign new_n2181 = ~new_n2179 & ~new_n2180 ;
  assign new_n2182 = lo1228 & ~new_n2139 ;
  assign new_n2183 = lo1229 & new_n2139 ;
  assign new_n2184 = ~new_n2182 & ~new_n2183 ;
  assign new_n2185 = new_n2071 & new_n2138 ;
  assign new_n2186 = lo1123 & new_n2185 ;
  assign new_n2187 = lo0018 & new_n1967 ;
  assign new_n2188 = new_n1993 & new_n2187 ;
  assign new_n2189 = lo0000 & ~new_n2188 ;
  assign new_n2190 = lo1269 & new_n2188 ;
  assign new_n2191 = ~new_n2189 & ~new_n2190 ;
  assign new_n2192 = lo0001 & ~new_n2188 ;
  assign new_n2193 = lo1270 & new_n2188 ;
  assign new_n2194 = ~new_n2192 & ~new_n2193 ;
  assign new_n2195 = lo0002 & ~new_n2188 ;
  assign new_n2196 = lo1271 & new_n2188 ;
  assign new_n2197 = ~new_n2195 & ~new_n2196 ;
  assign new_n2198 = new_n2011 & new_n2187 ;
  assign new_n2199 = lo0003 & ~new_n2198 ;
  assign new_n2200 = lo1272 & new_n2198 ;
  assign new_n2201 = ~new_n2199 & ~new_n2200 ;
  assign new_n2202 = lo0004 & ~new_n2198 ;
  assign new_n2203 = lo1273 & new_n2198 ;
  assign new_n2204 = ~new_n2202 & ~new_n2203 ;
  assign new_n2205 = lo0005 & ~new_n2198 ;
  assign new_n2206 = lo1274 & new_n2198 ;
  assign new_n2207 = ~new_n2205 & ~new_n2206 ;
  assign new_n2208 = lo0006 & ~new_n2198 ;
  assign new_n2209 = lo1275 & new_n2198 ;
  assign new_n2210 = ~new_n2208 & ~new_n2209 ;
  assign new_n2211 = lo0007 & ~new_n2198 ;
  assign new_n2212 = lo1276 & new_n2198 ;
  assign new_n2213 = ~new_n2211 & ~new_n2212 ;
  assign new_n2214 = lo0008 & ~new_n2198 ;
  assign new_n2215 = lo1277 & new_n2198 ;
  assign new_n2216 = ~new_n2214 & ~new_n2215 ;
  assign new_n2217 = lo0009 & ~new_n2198 ;
  assign new_n2218 = lo1278 & new_n2198 ;
  assign new_n2219 = ~new_n2217 & ~new_n2218 ;
  assign new_n2220 = lo0010 & ~new_n2198 ;
  assign new_n2221 = lo1279 & new_n2198 ;
  assign new_n2222 = ~new_n2220 & ~new_n2221 ;
  assign new_n2223 = new_n1942 & new_n2187 ;
  assign new_n2224 = lo0011 & ~new_n2223 ;
  assign new_n2225 = lo1280 & new_n2223 ;
  assign new_n2226 = ~new_n2224 & ~new_n2225 ;
  assign new_n2227 = lo0012 & ~new_n2223 ;
  assign new_n2228 = lo1281 & new_n2223 ;
  assign new_n2229 = ~new_n2227 & ~new_n2228 ;
  assign new_n2230 = lo0013 & ~new_n2223 ;
  assign new_n2231 = lo1282 & new_n2223 ;
  assign new_n2232 = ~new_n2230 & ~new_n2231 ;
  assign new_n2233 = lo0014 & ~new_n2223 ;
  assign new_n2234 = lo1283 & new_n2223 ;
  assign new_n2235 = ~new_n2233 & ~new_n2234 ;
  assign new_n2236 = lo0015 & ~new_n2223 ;
  assign new_n2237 = lo1284 & new_n2223 ;
  assign new_n2238 = ~new_n2236 & ~new_n2237 ;
  assign new_n2239 = lo0053 & ~lo0054 ;
  assign new_n2240 = ~lo0053 & lo0054 ;
  assign new_n2241 = ~new_n2239 & ~new_n2240 ;
  assign new_n2242 = lo0051 & ~lo0052 ;
  assign new_n2243 = ~lo0051 & lo0052 ;
  assign new_n2244 = ~new_n2242 & ~new_n2243 ;
  assign new_n2245 = new_n2241 & new_n2244 ;
  assign new_n2246 = lo1285 & new_n2245 ;
  assign new_n2247 = lo0018 & ~lo0022 ;
  assign new_n2248 = lo0115 & lo0116 ;
  assign new_n2249 = ~new_n2247 & ~new_n2248 ;
  assign new_n2250 = ~lo0118 & lo0119 ;
  assign new_n2251 = ~lo0117 & ~new_n2250 ;
  assign new_n2252 = new_n2249 & ~new_n2251 ;
  assign new_n2253 = lo0018 & new_n2252 ;
  assign new_n2254 = lo0117 & new_n2249 ;
  assign new_n2255 = ~lo0117 & ~new_n2249 ;
  assign new_n2256 = lo0118 & ~lo0119 ;
  assign new_n2257 = ~new_n2250 & ~new_n2256 ;
  assign new_n2258 = ~lo0118 & ~new_n2257 ;
  assign new_n2259 = ~new_n2255 & new_n2258 ;
  assign new_n2260 = lo0120 & ~new_n2259 ;
  assign new_n2261 = ~new_n2254 & ~new_n2260 ;
  assign new_n2262 = ~lo1293 & ~lo1294 ;
  assign new_n2263 = ~lo1292 & new_n2262 ;
  assign new_n2264 = ~lo1291 & new_n2263 ;
  assign new_n2265 = ~lo0122 & new_n2264 ;
  assign new_n2266 = lo0121 & ~new_n2265 ;
  assign new_n2267 = ~lo0124 & ~lo0125 ;
  assign new_n2268 = lo0123 & ~new_n2267 ;
  assign new_n2269 = lo0126 & lo0127 ;
  assign new_n2270 = ~lo0126 & lo0128 ;
  assign new_n2271 = ~new_n2269 & ~new_n2270 ;
  assign new_n2272 = new_n2267 & ~new_n2271 ;
  assign new_n2273 = ~new_n2268 & ~new_n2272 ;
  assign new_n2274 = lo0130 & ~new_n2267 ;
  assign new_n2275 = lo0126 & lo0131 ;
  assign new_n2276 = ~lo0126 & lo0132 ;
  assign new_n2277 = ~new_n2275 & ~new_n2276 ;
  assign new_n2278 = new_n2267 & ~new_n2277 ;
  assign new_n2279 = ~new_n2274 & ~new_n2278 ;
  assign new_n2280 = lo0133 & ~new_n2267 ;
  assign new_n2281 = lo0126 & lo0134 ;
  assign new_n2282 = ~lo0126 & lo0135 ;
  assign new_n2283 = ~new_n2281 & ~new_n2282 ;
  assign new_n2284 = new_n2267 & ~new_n2283 ;
  assign new_n2285 = ~new_n2280 & ~new_n2284 ;
  assign new_n2286 = ~new_n2279 & ~new_n2285 ;
  assign new_n2287 = lo0139 & ~new_n2267 ;
  assign new_n2288 = lo0126 & lo0140 ;
  assign new_n2289 = ~lo0126 & lo0141 ;
  assign new_n2290 = ~new_n2288 & ~new_n2289 ;
  assign new_n2291 = new_n2267 & ~new_n2290 ;
  assign new_n2292 = ~new_n2287 & ~new_n2291 ;
  assign new_n2293 = lo0142 & ~new_n2267 ;
  assign new_n2294 = lo0126 & lo0143 ;
  assign new_n2295 = ~lo0126 & lo0144 ;
  assign new_n2296 = ~new_n2294 & ~new_n2295 ;
  assign new_n2297 = new_n2267 & ~new_n2296 ;
  assign new_n2298 = ~new_n2293 & ~new_n2297 ;
  assign new_n2299 = new_n2292 & new_n2298 ;
  assign new_n2300 = lo0145 & ~new_n2267 ;
  assign new_n2301 = lo0126 & lo0146 ;
  assign new_n2302 = ~lo0126 & lo0147 ;
  assign new_n2303 = ~new_n2301 & ~new_n2302 ;
  assign new_n2304 = new_n2267 & ~new_n2303 ;
  assign new_n2305 = ~new_n2300 & ~new_n2304 ;
  assign new_n2306 = lo0136 & ~new_n2267 ;
  assign new_n2307 = lo0126 & lo0137 ;
  assign new_n2308 = ~lo0126 & lo0138 ;
  assign new_n2309 = ~new_n2307 & ~new_n2308 ;
  assign new_n2310 = new_n2267 & ~new_n2309 ;
  assign new_n2311 = ~new_n2306 & ~new_n2310 ;
  assign new_n2312 = lo0148 & ~new_n2267 ;
  assign new_n2313 = lo0126 & lo0149 ;
  assign new_n2314 = ~lo0126 & lo0150 ;
  assign new_n2315 = ~new_n2313 & ~new_n2314 ;
  assign new_n2316 = new_n2267 & ~new_n2315 ;
  assign new_n2317 = ~new_n2312 & ~new_n2316 ;
  assign new_n2318 = new_n2311 & new_n2317 ;
  assign new_n2319 = ~new_n2305 & new_n2318 ;
  assign new_n2320 = new_n2299 & new_n2319 ;
  assign new_n2321 = ~new_n2279 & ~new_n2320 ;
  assign new_n2322 = new_n2285 & ~new_n2321 ;
  assign new_n2323 = ~new_n2286 & ~new_n2322 ;
  assign new_n2324 = lo0151 & ~new_n2267 ;
  assign new_n2325 = lo0126 & lo0152 ;
  assign new_n2326 = ~lo0126 & lo0153 ;
  assign new_n2327 = ~new_n2325 & ~new_n2326 ;
  assign new_n2328 = new_n2267 & ~new_n2327 ;
  assign new_n2329 = ~new_n2324 & ~new_n2328 ;
  assign new_n2330 = lo0160 & ~new_n2267 ;
  assign new_n2331 = lo0126 & lo0161 ;
  assign new_n2332 = ~lo0126 & lo0162 ;
  assign new_n2333 = ~new_n2331 & ~new_n2332 ;
  assign new_n2334 = new_n2267 & ~new_n2333 ;
  assign new_n2335 = ~new_n2330 & ~new_n2334 ;
  assign new_n2336 = new_n2273 & new_n2335 ;
  assign new_n2337 = new_n2329 & new_n2336 ;
  assign new_n2338 = lo0154 & ~new_n2267 ;
  assign new_n2339 = lo0126 & lo0155 ;
  assign new_n2340 = ~lo0126 & lo0156 ;
  assign new_n2341 = ~new_n2339 & ~new_n2340 ;
  assign new_n2342 = new_n2267 & ~new_n2341 ;
  assign new_n2343 = ~new_n2338 & ~new_n2342 ;
  assign new_n2344 = lo0157 & ~new_n2267 ;
  assign new_n2345 = lo0126 & lo0158 ;
  assign new_n2346 = ~lo0126 & lo0159 ;
  assign new_n2347 = ~new_n2345 & ~new_n2346 ;
  assign new_n2348 = new_n2267 & ~new_n2347 ;
  assign new_n2349 = ~new_n2344 & ~new_n2348 ;
  assign new_n2350 = new_n2343 & new_n2349 ;
  assign new_n2351 = lo0169 & ~new_n2267 ;
  assign new_n2352 = lo0126 & lo0170 ;
  assign new_n2353 = ~lo0126 & lo0171 ;
  assign new_n2354 = ~new_n2352 & ~new_n2353 ;
  assign new_n2355 = new_n2267 & ~new_n2354 ;
  assign new_n2356 = ~new_n2351 & ~new_n2355 ;
  assign new_n2357 = lo0172 & ~new_n2267 ;
  assign new_n2358 = lo0126 & lo0173 ;
  assign new_n2359 = ~lo0126 & lo0174 ;
  assign new_n2360 = ~new_n2358 & ~new_n2359 ;
  assign new_n2361 = new_n2267 & ~new_n2360 ;
  assign new_n2362 = ~new_n2357 & ~new_n2361 ;
  assign new_n2363 = new_n2356 & ~new_n2362 ;
  assign new_n2364 = lo0163 & ~new_n2267 ;
  assign new_n2365 = lo0126 & lo0164 ;
  assign new_n2366 = ~lo0126 & lo0165 ;
  assign new_n2367 = ~new_n2365 & ~new_n2366 ;
  assign new_n2368 = new_n2267 & ~new_n2367 ;
  assign new_n2369 = ~new_n2364 & ~new_n2368 ;
  assign new_n2370 = lo0166 & ~new_n2267 ;
  assign new_n2371 = lo0126 & lo0167 ;
  assign new_n2372 = ~lo0126 & lo0168 ;
  assign new_n2373 = ~new_n2371 & ~new_n2372 ;
  assign new_n2374 = new_n2267 & ~new_n2373 ;
  assign new_n2375 = ~new_n2370 & ~new_n2374 ;
  assign new_n2376 = new_n2369 & ~new_n2375 ;
  assign new_n2377 = new_n2363 & new_n2376 ;
  assign new_n2378 = new_n2350 & new_n2377 ;
  assign new_n2379 = new_n2337 & new_n2378 ;
  assign new_n2380 = ~new_n2323 & new_n2379 ;
  assign new_n2381 = new_n2285 & ~new_n2343 ;
  assign new_n2382 = ~new_n2285 & ~new_n2311 ;
  assign new_n2383 = new_n2299 & new_n2382 ;
  assign new_n2384 = new_n2350 & new_n2383 ;
  assign new_n2385 = ~new_n2298 & ~new_n2349 ;
  assign new_n2386 = ~new_n2311 & ~new_n2343 ;
  assign new_n2387 = new_n2385 & new_n2386 ;
  assign new_n2388 = new_n2285 & new_n2349 ;
  assign new_n2389 = ~new_n2387 & ~new_n2388 ;
  assign new_n2390 = ~new_n2292 & ~new_n2389 ;
  assign new_n2391 = ~new_n2384 & ~new_n2390 ;
  assign new_n2392 = ~new_n2317 & ~new_n2391 ;
  assign new_n2393 = ~new_n2381 & ~new_n2392 ;
  assign new_n2394 = ~new_n2273 & ~new_n2393 ;
  assign new_n2395 = ~new_n2380 & ~new_n2394 ;
  assign new_n2396 = lo0129 & new_n2395 ;
  assign new_n2397 = ~new_n2273 & ~new_n2317 ;
  assign new_n2398 = ~new_n2285 & ~new_n2292 ;
  assign new_n2399 = new_n2397 & new_n2398 ;
  assign new_n2400 = new_n2387 & new_n2399 ;
  assign new_n2401 = ~lo0129 & ~new_n2400 ;
  assign new_n2402 = ~new_n2396 & ~new_n2401 ;
  assign new_n2403 = ~lo0176 & ~lo0177 ;
  assign new_n2404 = ~lo0175 & new_n2403 ;
  assign new_n2405 = lo0179 & ~lo0180 ;
  assign new_n2406 = ~lo0175 & ~new_n2405 ;
  assign new_n2407 = ~lo0177 & ~new_n2406 ;
  assign new_n2408 = ~lo0176 & ~new_n2407 ;
  assign new_n2409 = ~lo0179 & ~lo0180 ;
  assign new_n2410 = ~lo0175 & ~lo0177 ;
  assign new_n2411 = new_n2409 & new_n2410 ;
  assign new_n2412 = ~lo0176 & ~new_n2411 ;
  assign new_n2413 = new_n2408 & new_n2412 ;
  assign new_n2414 = ~lo0180 & new_n2404 ;
  assign new_n2415 = ~lo0182 & new_n2414 ;
  assign new_n2416 = ~lo0181 & ~new_n2415 ;
  assign new_n2417 = ~lo0184 & new_n2414 ;
  assign new_n2418 = ~lo0183 & ~new_n2417 ;
  assign new_n2419 = ~lo0186 & new_n2414 ;
  assign new_n2420 = ~lo0185 & ~new_n2419 ;
  assign new_n2421 = lo0185 & new_n2419 ;
  assign new_n2422 = ~lo0188 & new_n2414 ;
  assign new_n2423 = ~lo0187 & ~new_n2422 ;
  assign new_n2424 = ~new_n2421 & new_n2423 ;
  assign new_n2425 = ~new_n2420 & new_n2424 ;
  assign new_n2426 = ~new_n2420 & ~new_n2425 ;
  assign new_n2427 = lo0183 & new_n2417 ;
  assign new_n2428 = ~new_n2418 & ~new_n2427 ;
  assign new_n2429 = ~new_n2426 & new_n2428 ;
  assign new_n2430 = ~new_n2418 & ~new_n2429 ;
  assign new_n2431 = lo0181 & new_n2415 ;
  assign new_n2432 = ~new_n2416 & ~new_n2431 ;
  assign new_n2433 = ~new_n2430 & new_n2432 ;
  assign new_n2434 = ~new_n2416 & ~new_n2433 ;
  assign new_n2435 = new_n2404 & ~new_n2409 ;
  assign new_n2436 = ~new_n2408 & new_n2412 ;
  assign new_n2437 = new_n2435 & new_n2436 ;
  assign new_n2438 = ~new_n2434 & new_n2437 ;
  assign new_n2439 = ~new_n2413 & ~new_n2438 ;
  assign new_n2440 = ~lo0178 & ~new_n2439 ;
  assign new_n2441 = new_n2404 & ~new_n2440 ;
  assign new_n2442 = ~lo0129 & ~new_n2441 ;
  assign new_n2443 = ~new_n2402 & ~new_n2442 ;
  assign new_n2444 = new_n2273 & new_n2443 ;
  assign new_n2445 = new_n2265 & ~new_n2444 ;
  assign new_n2446 = ~new_n2266 & ~new_n2445 ;
  assign new_n2447 = lo0189 & ~new_n2265 ;
  assign new_n2448 = new_n2343 & new_n2443 ;
  assign new_n2449 = new_n2265 & ~new_n2448 ;
  assign new_n2450 = ~new_n2447 & ~new_n2449 ;
  assign new_n2451 = lo0190 & ~new_n2265 ;
  assign new_n2452 = new_n2349 & new_n2443 ;
  assign new_n2453 = new_n2265 & ~new_n2452 ;
  assign new_n2454 = ~new_n2451 & ~new_n2453 ;
  assign new_n2455 = new_n2450 & new_n2454 ;
  assign new_n2456 = ~lo1291 & new_n2262 ;
  assign new_n2457 = lo0194 & ~new_n2265 ;
  assign new_n2458 = new_n2404 & new_n2442 ;
  assign new_n2459 = ~new_n2443 & ~new_n2458 ;
  assign new_n2460 = new_n2409 & new_n2442 ;
  assign new_n2461 = ~new_n2311 & ~new_n2442 ;
  assign new_n2462 = ~new_n2460 & ~new_n2461 ;
  assign new_n2463 = ~new_n2459 & new_n2462 ;
  assign new_n2464 = new_n2265 & ~new_n2463 ;
  assign new_n2465 = ~new_n2457 & ~new_n2464 ;
  assign new_n2466 = ~lo0062 & lo0251 ;
  assign new_n2467 = ~lo0058 & lo0249 ;
  assign new_n2468 = lo0060 & ~lo0250 ;
  assign new_n2469 = ~new_n2467 & ~new_n2468 ;
  assign new_n2470 = ~new_n2466 & new_n2469 ;
  assign new_n2471 = ~lo0064 & lo0252 ;
  assign new_n2472 = lo0057 & lo0247 ;
  assign new_n2473 = ~new_n2471 & new_n2472 ;
  assign new_n2474 = lo0058 & ~lo0249 ;
  assign new_n2475 = lo0064 & ~lo0252 ;
  assign new_n2476 = ~new_n2474 & ~new_n2475 ;
  assign new_n2477 = ~lo0060 & lo0250 ;
  assign new_n2478 = lo0062 & ~lo0251 ;
  assign new_n2479 = ~new_n2477 & ~new_n2478 ;
  assign new_n2480 = new_n2476 & new_n2479 ;
  assign new_n2481 = new_n2473 & new_n2480 ;
  assign new_n2482 = new_n2470 & new_n2481 ;
  assign new_n2483 = ~lo0248 & ~new_n2482 ;
  assign new_n2484 = ~lo0254 & ~lo0255 ;
  assign new_n2485 = ~lo0253 & new_n2484 ;
  assign new_n2486 = ~lo0256 & ~lo0257 ;
  assign new_n2487 = lo0247 & new_n2486 ;
  assign new_n2488 = new_n2485 & new_n2487 ;
  assign new_n2489 = new_n2483 & new_n2488 ;
  assign new_n2490 = ~lo0249 & ~lo0250 ;
  assign new_n2491 = lo0745 & new_n2490 ;
  assign new_n2492 = lo0249 & lo0250 ;
  assign new_n2493 = ~lo0249 & lo0250 ;
  assign new_n2494 = lo0744 & new_n2493 ;
  assign new_n2495 = ~new_n2492 & ~new_n2494 ;
  assign new_n2496 = ~new_n2491 & new_n2495 ;
  assign new_n2497 = ~lo0249 & ~new_n2496 ;
  assign new_n2498 = lo0249 & new_n2496 ;
  assign new_n2499 = ~new_n2497 & ~new_n2498 ;
  assign new_n2500 = lo0743 & ~new_n2499 ;
  assign new_n2501 = ~lo0743 & new_n2497 ;
  assign new_n2502 = lo0249 & lo0746 ;
  assign new_n2503 = ~new_n2496 & new_n2502 ;
  assign new_n2504 = ~new_n2501 & ~new_n2503 ;
  assign new_n2505 = ~new_n2500 & new_n2504 ;
  assign new_n2506 = ~lo0251 & ~lo0252 ;
  assign new_n2507 = lo0742 & new_n2490 ;
  assign new_n2508 = lo0752 & new_n2493 ;
  assign new_n2509 = ~new_n2492 & ~new_n2508 ;
  assign new_n2510 = ~new_n2507 & new_n2509 ;
  assign new_n2511 = ~lo0249 & ~new_n2510 ;
  assign new_n2512 = lo0249 & new_n2510 ;
  assign new_n2513 = ~new_n2511 & ~new_n2512 ;
  assign new_n2514 = lo0751 & ~new_n2513 ;
  assign new_n2515 = ~lo0751 & new_n2511 ;
  assign new_n2516 = lo0249 & lo0753 ;
  assign new_n2517 = ~new_n2510 & new_n2516 ;
  assign new_n2518 = ~new_n2515 & ~new_n2517 ;
  assign new_n2519 = ~new_n2514 & new_n2518 ;
  assign new_n2520 = new_n2506 & ~new_n2519 ;
  assign new_n2521 = lo0251 & lo0252 ;
  assign new_n2522 = ~lo0251 & lo0252 ;
  assign new_n2523 = lo0749 & new_n2490 ;
  assign new_n2524 = ~lo0250 & lo0748 ;
  assign new_n2525 = lo0249 & new_n2524 ;
  assign new_n2526 = ~new_n2492 & ~new_n2525 ;
  assign new_n2527 = ~new_n2523 & new_n2526 ;
  assign new_n2528 = ~lo0250 & ~new_n2527 ;
  assign new_n2529 = lo0250 & new_n2527 ;
  assign new_n2530 = ~new_n2528 & ~new_n2529 ;
  assign new_n2531 = lo0747 & ~new_n2530 ;
  assign new_n2532 = ~lo0747 & new_n2528 ;
  assign new_n2533 = lo0250 & lo0750 ;
  assign new_n2534 = ~new_n2527 & new_n2533 ;
  assign new_n2535 = ~new_n2532 & ~new_n2534 ;
  assign new_n2536 = ~new_n2531 & new_n2535 ;
  assign new_n2537 = new_n2522 & ~new_n2536 ;
  assign new_n2538 = ~new_n2521 & ~new_n2537 ;
  assign new_n2539 = ~new_n2520 & new_n2538 ;
  assign new_n2540 = ~lo0251 & ~new_n2539 ;
  assign new_n2541 = lo0251 & new_n2539 ;
  assign new_n2542 = ~new_n2540 & ~new_n2541 ;
  assign new_n2543 = ~new_n2505 & ~new_n2542 ;
  assign new_n2544 = new_n2505 & new_n2540 ;
  assign new_n2545 = lo0756 & new_n2490 ;
  assign new_n2546 = ~lo0250 & lo0755 ;
  assign new_n2547 = lo0249 & new_n2546 ;
  assign new_n2548 = ~new_n2492 & ~new_n2547 ;
  assign new_n2549 = ~new_n2545 & new_n2548 ;
  assign new_n2550 = ~lo0250 & ~new_n2549 ;
  assign new_n2551 = lo0250 & new_n2549 ;
  assign new_n2552 = ~new_n2550 & ~new_n2551 ;
  assign new_n2553 = lo0754 & ~new_n2552 ;
  assign new_n2554 = ~lo0754 & new_n2550 ;
  assign new_n2555 = lo0250 & lo0757 ;
  assign new_n2556 = ~new_n2549 & new_n2555 ;
  assign new_n2557 = ~new_n2554 & ~new_n2556 ;
  assign new_n2558 = ~new_n2553 & new_n2557 ;
  assign new_n2559 = lo0251 & ~new_n2558 ;
  assign new_n2560 = ~new_n2539 & new_n2559 ;
  assign new_n2561 = ~new_n2544 & ~new_n2560 ;
  assign new_n2562 = ~new_n2543 & new_n2561 ;
  assign new_n2563 = new_n2489 & ~new_n2562 ;
  assign new_n2564 = ~lo0093 & ~lo0095 ;
  assign new_n2565 = ~lo0091 & new_n2564 ;
  assign new_n2566 = ~lo0092 & new_n2565 ;
  assign new_n2567 = lo0092 & ~new_n2564 ;
  assign new_n2568 = ~lo0091 & ~new_n2567 ;
  assign new_n2569 = ~new_n2566 & new_n2568 ;
  assign new_n2570 = lo0099 & new_n2565 ;
  assign new_n2571 = new_n2569 & new_n2570 ;
  assign new_n2572 = ~new_n2565 & ~new_n2569 ;
  assign new_n2573 = lo0555 & ~new_n2565 ;
  assign new_n2574 = new_n2569 & new_n2573 ;
  assign new_n2575 = ~new_n2572 & ~new_n2574 ;
  assign new_n2576 = ~new_n2571 & new_n2575 ;
  assign new_n2577 = new_n2569 & ~new_n2576 ;
  assign new_n2578 = ~new_n2569 & new_n2576 ;
  assign new_n2579 = ~new_n2577 & ~new_n2578 ;
  assign new_n2580 = lo0100 & ~new_n2579 ;
  assign new_n2581 = ~lo0100 & new_n2577 ;
  assign new_n2582 = lo0758 & ~new_n2569 ;
  assign new_n2583 = ~new_n2576 & new_n2582 ;
  assign new_n2584 = ~new_n2581 & ~new_n2583 ;
  assign new_n2585 = ~new_n2580 & new_n2584 ;
  assign new_n2586 = lo0090 & ~new_n2585 ;
  assign new_n2587 = ~new_n2483 & new_n2586 ;
  assign new_n2588 = ~lo0247 & ~lo0248 ;
  assign new_n2589 = new_n2485 & new_n2588 ;
  assign new_n2590 = ~lo0256 & lo0257 ;
  assign new_n2591 = new_n2589 & new_n2590 ;
  assign new_n2592 = ~lo0107 & ~lo0108 ;
  assign new_n2593 = ~lo0102 & lo0222 ;
  assign new_n2594 = ~lo0103 & new_n2593 ;
  assign new_n2595 = ~lo0105 & ~new_n2594 ;
  assign new_n2596 = new_n2592 & ~new_n2595 ;
  assign new_n2597 = ~lo0106 & ~new_n2596 ;
  assign new_n2598 = lo0641 & ~new_n2597 ;
  assign new_n2599 = new_n2591 & new_n2598 ;
  assign new_n2600 = lo0256 & ~lo0257 ;
  assign new_n2601 = new_n2589 & new_n2600 ;
  assign new_n2602 = lo0759 & new_n2601 ;
  assign new_n2603 = new_n2486 & new_n2588 ;
  assign new_n2604 = lo0253 & new_n2484 ;
  assign new_n2605 = new_n2603 & new_n2604 ;
  assign new_n2606 = lo0762 & new_n2605 ;
  assign new_n2607 = ~new_n2602 & ~new_n2606 ;
  assign new_n2608 = ~lo0253 & new_n2603 ;
  assign new_n2609 = ~lo0254 & lo0255 ;
  assign new_n2610 = new_n2608 & new_n2609 ;
  assign new_n2611 = lo1360 & new_n2610 ;
  assign new_n2612 = lo0254 & ~lo0255 ;
  assign new_n2613 = new_n2608 & new_n2612 ;
  assign new_n2614 = lo0761 & new_n2613 ;
  assign new_n2615 = ~new_n2611 & ~new_n2614 ;
  assign new_n2616 = new_n2607 & new_n2615 ;
  assign new_n2617 = ~new_n2599 & new_n2616 ;
  assign new_n2618 = ~new_n2587 & new_n2617 ;
  assign new_n2619 = ~new_n2563 & new_n2618 ;
  assign new_n2620 = lo0298 & ~new_n2619 ;
  assign new_n2621 = ~lo0249 & lo0462 ;
  assign new_n2622 = ~lo0250 & new_n2621 ;
  assign new_n2623 = ~lo0249 & lo0461 ;
  assign new_n2624 = lo0250 & new_n2623 ;
  assign new_n2625 = ~new_n2492 & ~new_n2624 ;
  assign new_n2626 = ~new_n2622 & new_n2625 ;
  assign new_n2627 = ~lo0249 & ~new_n2626 ;
  assign new_n2628 = lo0249 & new_n2626 ;
  assign new_n2629 = ~new_n2627 & ~new_n2628 ;
  assign new_n2630 = lo0460 & ~new_n2629 ;
  assign new_n2631 = ~lo0460 & new_n2627 ;
  assign new_n2632 = lo0249 & lo0463 ;
  assign new_n2633 = ~new_n2626 & new_n2632 ;
  assign new_n2634 = ~new_n2631 & ~new_n2633 ;
  assign new_n2635 = ~new_n2630 & new_n2634 ;
  assign new_n2636 = ~lo0249 & lo0470 ;
  assign new_n2637 = ~lo0250 & new_n2636 ;
  assign new_n2638 = ~lo0249 & lo0469 ;
  assign new_n2639 = lo0250 & new_n2638 ;
  assign new_n2640 = ~new_n2492 & ~new_n2639 ;
  assign new_n2641 = ~new_n2637 & new_n2640 ;
  assign new_n2642 = ~lo0249 & ~new_n2641 ;
  assign new_n2643 = lo0249 & new_n2641 ;
  assign new_n2644 = ~new_n2642 & ~new_n2643 ;
  assign new_n2645 = lo0468 & ~new_n2644 ;
  assign new_n2646 = ~lo0468 & new_n2642 ;
  assign new_n2647 = lo0249 & lo0471 ;
  assign new_n2648 = ~new_n2641 & new_n2647 ;
  assign new_n2649 = ~new_n2646 & ~new_n2648 ;
  assign new_n2650 = ~new_n2645 & new_n2649 ;
  assign new_n2651 = new_n2506 & ~new_n2650 ;
  assign new_n2652 = ~lo0250 & lo0466 ;
  assign new_n2653 = ~lo0249 & new_n2652 ;
  assign new_n2654 = ~lo0250 & lo0465 ;
  assign new_n2655 = lo0249 & new_n2654 ;
  assign new_n2656 = ~new_n2492 & ~new_n2655 ;
  assign new_n2657 = ~new_n2653 & new_n2656 ;
  assign new_n2658 = ~lo0250 & ~new_n2657 ;
  assign new_n2659 = lo0250 & new_n2657 ;
  assign new_n2660 = ~new_n2658 & ~new_n2659 ;
  assign new_n2661 = lo0464 & ~new_n2660 ;
  assign new_n2662 = ~lo0464 & new_n2658 ;
  assign new_n2663 = lo0250 & lo0467 ;
  assign new_n2664 = ~new_n2657 & new_n2663 ;
  assign new_n2665 = ~new_n2662 & ~new_n2664 ;
  assign new_n2666 = ~new_n2661 & new_n2665 ;
  assign new_n2667 = new_n2522 & ~new_n2666 ;
  assign new_n2668 = ~new_n2521 & ~new_n2667 ;
  assign new_n2669 = ~new_n2651 & new_n2668 ;
  assign new_n2670 = ~lo0251 & ~new_n2669 ;
  assign new_n2671 = lo0251 & new_n2669 ;
  assign new_n2672 = ~new_n2670 & ~new_n2671 ;
  assign new_n2673 = ~new_n2635 & ~new_n2672 ;
  assign new_n2674 = new_n2635 & new_n2670 ;
  assign new_n2675 = ~lo0250 & lo0474 ;
  assign new_n2676 = ~lo0249 & new_n2675 ;
  assign new_n2677 = ~lo0250 & lo0473 ;
  assign new_n2678 = lo0249 & new_n2677 ;
  assign new_n2679 = ~new_n2492 & ~new_n2678 ;
  assign new_n2680 = ~new_n2676 & new_n2679 ;
  assign new_n2681 = ~lo0250 & ~new_n2680 ;
  assign new_n2682 = lo0250 & new_n2680 ;
  assign new_n2683 = ~new_n2681 & ~new_n2682 ;
  assign new_n2684 = lo0472 & ~new_n2683 ;
  assign new_n2685 = ~lo0472 & new_n2681 ;
  assign new_n2686 = lo0250 & lo0475 ;
  assign new_n2687 = ~new_n2680 & new_n2686 ;
  assign new_n2688 = ~new_n2685 & ~new_n2687 ;
  assign new_n2689 = ~new_n2684 & new_n2688 ;
  assign new_n2690 = lo0251 & ~new_n2689 ;
  assign new_n2691 = ~new_n2669 & new_n2690 ;
  assign new_n2692 = ~new_n2674 & ~new_n2691 ;
  assign new_n2693 = ~new_n2673 & new_n2692 ;
  assign new_n2694 = new_n2489 & ~new_n2693 ;
  assign new_n2695 = ~lo0092 & lo0097 ;
  assign new_n2696 = ~lo0095 & new_n2695 ;
  assign new_n2697 = lo0092 & lo0095 ;
  assign new_n2698 = lo0092 & lo0096 ;
  assign new_n2699 = ~lo0095 & new_n2698 ;
  assign new_n2700 = ~new_n2697 & ~new_n2699 ;
  assign new_n2701 = ~new_n2696 & new_n2700 ;
  assign new_n2702 = ~lo0095 & ~new_n2701 ;
  assign new_n2703 = lo0095 & new_n2701 ;
  assign new_n2704 = ~new_n2702 & ~new_n2703 ;
  assign new_n2705 = lo0094 & ~new_n2704 ;
  assign new_n2706 = ~lo0094 & new_n2702 ;
  assign new_n2707 = lo0095 & lo0098 ;
  assign new_n2708 = ~new_n2701 & new_n2707 ;
  assign new_n2709 = ~new_n2706 & ~new_n2708 ;
  assign new_n2710 = ~new_n2705 & new_n2709 ;
  assign new_n2711 = ~lo0093 & ~new_n2710 ;
  assign new_n2712 = ~new_n2695 & ~new_n2698 ;
  assign new_n2713 = lo0093 & ~new_n2712 ;
  assign new_n2714 = ~new_n2711 & ~new_n2713 ;
  assign new_n2715 = ~lo0091 & ~new_n2714 ;
  assign new_n2716 = lo0091 & lo0097 ;
  assign new_n2717 = ~new_n2715 & ~new_n2716 ;
  assign new_n2718 = lo0090 & ~new_n2717 ;
  assign new_n2719 = ~new_n2483 & new_n2718 ;
  assign new_n2720 = ~lo0222 & ~lo0228 ;
  assign new_n2721 = lo0104 & ~new_n2720 ;
  assign new_n2722 = lo0229 & new_n2720 ;
  assign new_n2723 = ~new_n2721 & ~new_n2722 ;
  assign new_n2724 = ~lo0106 & new_n2592 ;
  assign new_n2725 = ~lo0105 & new_n2724 ;
  assign new_n2726 = ~lo0103 & new_n2725 ;
  assign new_n2727 = ~lo0102 & new_n2726 ;
  assign new_n2728 = ~new_n2723 & new_n2727 ;
  assign new_n2729 = new_n2591 & new_n2728 ;
  assign new_n2730 = lo0476 & new_n2601 ;
  assign new_n2731 = lo0478 & new_n2605 ;
  assign new_n2732 = ~new_n2730 & ~new_n2731 ;
  assign new_n2733 = lo0477 & new_n2613 ;
  assign new_n2734 = lo1319 & new_n2610 ;
  assign new_n2735 = ~new_n2733 & ~new_n2734 ;
  assign new_n2736 = new_n2732 & new_n2735 ;
  assign new_n2737 = ~new_n2729 & new_n2736 ;
  assign new_n2738 = ~new_n2719 & new_n2737 ;
  assign new_n2739 = ~new_n2694 & new_n2738 ;
  assign new_n2740 = ~lo0298 & ~new_n2739 ;
  assign new_n2741 = ~new_n2620 & ~new_n2740 ;
  assign new_n2742 = lo0853 & ~new_n2741 ;
  assign new_n2743 = lo0605 & new_n2490 ;
  assign new_n2744 = lo0604 & new_n2493 ;
  assign new_n2745 = ~new_n2492 & ~new_n2744 ;
  assign new_n2746 = ~new_n2743 & new_n2745 ;
  assign new_n2747 = ~lo0249 & ~new_n2746 ;
  assign new_n2748 = lo0249 & new_n2746 ;
  assign new_n2749 = ~new_n2747 & ~new_n2748 ;
  assign new_n2750 = lo0603 & ~new_n2749 ;
  assign new_n2751 = ~lo0603 & new_n2747 ;
  assign new_n2752 = lo0249 & lo0606 ;
  assign new_n2753 = ~new_n2746 & new_n2752 ;
  assign new_n2754 = ~new_n2751 & ~new_n2753 ;
  assign new_n2755 = ~new_n2750 & new_n2754 ;
  assign new_n2756 = lo0613 & new_n2490 ;
  assign new_n2757 = lo0612 & new_n2493 ;
  assign new_n2758 = ~new_n2492 & ~new_n2757 ;
  assign new_n2759 = ~new_n2756 & new_n2758 ;
  assign new_n2760 = ~lo0249 & ~new_n2759 ;
  assign new_n2761 = lo0249 & new_n2759 ;
  assign new_n2762 = ~new_n2760 & ~new_n2761 ;
  assign new_n2763 = lo0611 & ~new_n2762 ;
  assign new_n2764 = ~lo0611 & new_n2760 ;
  assign new_n2765 = lo0249 & lo0614 ;
  assign new_n2766 = ~new_n2759 & new_n2765 ;
  assign new_n2767 = ~new_n2764 & ~new_n2766 ;
  assign new_n2768 = ~new_n2763 & new_n2767 ;
  assign new_n2769 = new_n2506 & ~new_n2768 ;
  assign new_n2770 = lo0609 & new_n2490 ;
  assign new_n2771 = ~lo0250 & lo0608 ;
  assign new_n2772 = lo0249 & new_n2771 ;
  assign new_n2773 = ~new_n2492 & ~new_n2772 ;
  assign new_n2774 = ~new_n2770 & new_n2773 ;
  assign new_n2775 = ~lo0250 & ~new_n2774 ;
  assign new_n2776 = lo0250 & new_n2774 ;
  assign new_n2777 = ~new_n2775 & ~new_n2776 ;
  assign new_n2778 = lo0607 & ~new_n2777 ;
  assign new_n2779 = ~lo0607 & new_n2775 ;
  assign new_n2780 = lo0250 & lo0610 ;
  assign new_n2781 = ~new_n2774 & new_n2780 ;
  assign new_n2782 = ~new_n2779 & ~new_n2781 ;
  assign new_n2783 = ~new_n2778 & new_n2782 ;
  assign new_n2784 = new_n2522 & ~new_n2783 ;
  assign new_n2785 = ~new_n2521 & ~new_n2784 ;
  assign new_n2786 = ~new_n2769 & new_n2785 ;
  assign new_n2787 = ~lo0251 & ~new_n2786 ;
  assign new_n2788 = lo0251 & new_n2786 ;
  assign new_n2789 = ~new_n2787 & ~new_n2788 ;
  assign new_n2790 = ~new_n2755 & ~new_n2789 ;
  assign new_n2791 = new_n2755 & new_n2787 ;
  assign new_n2792 = lo0617 & new_n2490 ;
  assign new_n2793 = ~lo0250 & lo0616 ;
  assign new_n2794 = lo0249 & new_n2793 ;
  assign new_n2795 = ~new_n2492 & ~new_n2794 ;
  assign new_n2796 = ~new_n2792 & new_n2795 ;
  assign new_n2797 = ~lo0250 & ~new_n2796 ;
  assign new_n2798 = lo0250 & new_n2796 ;
  assign new_n2799 = ~new_n2797 & ~new_n2798 ;
  assign new_n2800 = lo0615 & ~new_n2799 ;
  assign new_n2801 = ~lo0615 & new_n2797 ;
  assign new_n2802 = lo0250 & lo0618 ;
  assign new_n2803 = ~new_n2796 & new_n2802 ;
  assign new_n2804 = ~new_n2801 & ~new_n2803 ;
  assign new_n2805 = ~new_n2800 & new_n2804 ;
  assign new_n2806 = lo0251 & ~new_n2805 ;
  assign new_n2807 = ~new_n2786 & new_n2806 ;
  assign new_n2808 = ~new_n2791 & ~new_n2807 ;
  assign new_n2809 = ~new_n2790 & new_n2808 ;
  assign new_n2810 = new_n2489 & ~new_n2809 ;
  assign new_n2811 = lo0091 & lo0094 ;
  assign new_n2812 = ~new_n2715 & ~new_n2811 ;
  assign new_n2813 = lo0090 & ~new_n2812 ;
  assign new_n2814 = ~new_n2483 & new_n2813 ;
  assign new_n2815 = lo0619 & new_n2601 ;
  assign new_n2816 = lo0621 & new_n2605 ;
  assign new_n2817 = ~new_n2815 & ~new_n2816 ;
  assign new_n2818 = lo0620 & new_n2613 ;
  assign new_n2819 = lo1344 & new_n2610 ;
  assign new_n2820 = ~new_n2818 & ~new_n2819 ;
  assign new_n2821 = new_n2817 & new_n2820 ;
  assign new_n2822 = ~new_n2729 & new_n2821 ;
  assign new_n2823 = ~new_n2814 & new_n2822 ;
  assign new_n2824 = ~new_n2810 & new_n2823 ;
  assign new_n2825 = lo0297 & ~lo0298 ;
  assign new_n2826 = ~lo0846 & new_n2825 ;
  assign new_n2827 = ~lo0299 & lo0300 ;
  assign new_n2828 = new_n2826 & new_n2827 ;
  assign new_n2829 = ~new_n2824 & new_n2828 ;
  assign new_n2830 = lo0404 & new_n2506 ;
  assign new_n2831 = lo0251 & ~lo0252 ;
  assign new_n2832 = lo0403 & new_n2831 ;
  assign new_n2833 = ~new_n2521 & ~new_n2832 ;
  assign new_n2834 = ~new_n2830 & new_n2833 ;
  assign new_n2835 = ~lo0252 & ~new_n2834 ;
  assign new_n2836 = lo0252 & new_n2834 ;
  assign new_n2837 = ~new_n2835 & ~new_n2836 ;
  assign new_n2838 = lo0402 & ~new_n2837 ;
  assign new_n2839 = ~lo0402 & new_n2835 ;
  assign new_n2840 = lo0252 & lo0405 ;
  assign new_n2841 = ~new_n2834 & new_n2840 ;
  assign new_n2842 = ~new_n2839 & ~new_n2841 ;
  assign new_n2843 = ~new_n2838 & new_n2842 ;
  assign new_n2844 = lo0401 & new_n2506 ;
  assign new_n2845 = lo0411 & new_n2831 ;
  assign new_n2846 = ~new_n2521 & ~new_n2845 ;
  assign new_n2847 = ~new_n2844 & new_n2846 ;
  assign new_n2848 = ~lo0252 & ~new_n2847 ;
  assign new_n2849 = lo0252 & new_n2847 ;
  assign new_n2850 = ~new_n2848 & ~new_n2849 ;
  assign new_n2851 = lo0410 & ~new_n2850 ;
  assign new_n2852 = ~lo0410 & new_n2848 ;
  assign new_n2853 = lo0252 & lo0412 ;
  assign new_n2854 = ~new_n2847 & new_n2853 ;
  assign new_n2855 = ~new_n2852 & ~new_n2854 ;
  assign new_n2856 = ~new_n2851 & new_n2855 ;
  assign new_n2857 = new_n2490 & ~new_n2856 ;
  assign new_n2858 = lo0408 & new_n2506 ;
  assign new_n2859 = lo0407 & new_n2522 ;
  assign new_n2860 = ~new_n2521 & ~new_n2859 ;
  assign new_n2861 = ~new_n2858 & new_n2860 ;
  assign new_n2862 = ~lo0251 & ~new_n2861 ;
  assign new_n2863 = lo0251 & new_n2861 ;
  assign new_n2864 = ~new_n2862 & ~new_n2863 ;
  assign new_n2865 = lo0406 & ~new_n2864 ;
  assign new_n2866 = ~lo0406 & new_n2862 ;
  assign new_n2867 = lo0251 & lo0409 ;
  assign new_n2868 = ~new_n2861 & new_n2867 ;
  assign new_n2869 = ~new_n2866 & ~new_n2868 ;
  assign new_n2870 = ~new_n2865 & new_n2869 ;
  assign new_n2871 = new_n2493 & ~new_n2870 ;
  assign new_n2872 = ~new_n2492 & ~new_n2871 ;
  assign new_n2873 = ~new_n2857 & new_n2872 ;
  assign new_n2874 = ~lo0249 & ~new_n2873 ;
  assign new_n2875 = lo0249 & new_n2873 ;
  assign new_n2876 = ~new_n2874 & ~new_n2875 ;
  assign new_n2877 = ~new_n2843 & ~new_n2876 ;
  assign new_n2878 = new_n2843 & new_n2874 ;
  assign new_n2879 = lo0415 & new_n2506 ;
  assign new_n2880 = lo0414 & new_n2522 ;
  assign new_n2881 = ~new_n2521 & ~new_n2880 ;
  assign new_n2882 = ~new_n2879 & new_n2881 ;
  assign new_n2883 = ~lo0251 & ~new_n2882 ;
  assign new_n2884 = lo0251 & new_n2882 ;
  assign new_n2885 = ~new_n2883 & ~new_n2884 ;
  assign new_n2886 = lo0413 & ~new_n2885 ;
  assign new_n2887 = ~lo0413 & new_n2883 ;
  assign new_n2888 = lo0251 & lo0416 ;
  assign new_n2889 = ~new_n2882 & new_n2888 ;
  assign new_n2890 = ~new_n2887 & ~new_n2889 ;
  assign new_n2891 = ~new_n2886 & new_n2890 ;
  assign new_n2892 = lo0249 & ~new_n2891 ;
  assign new_n2893 = ~new_n2873 & new_n2892 ;
  assign new_n2894 = ~new_n2878 & ~new_n2893 ;
  assign new_n2895 = ~new_n2877 & new_n2894 ;
  assign new_n2896 = new_n2489 & ~new_n2895 ;
  assign new_n2897 = lo0091 & lo0096 ;
  assign new_n2898 = ~new_n2715 & ~new_n2897 ;
  assign new_n2899 = lo0090 & ~new_n2898 ;
  assign new_n2900 = ~new_n2483 & new_n2899 ;
  assign new_n2901 = lo0417 & new_n2601 ;
  assign new_n2902 = lo0538 & new_n2605 ;
  assign new_n2903 = ~new_n2901 & ~new_n2902 ;
  assign new_n2904 = lo0418 & new_n2613 ;
  assign new_n2905 = lo1314 & new_n2610 ;
  assign new_n2906 = ~new_n2904 & ~new_n2905 ;
  assign new_n2907 = new_n2903 & new_n2906 ;
  assign new_n2908 = ~new_n2729 & new_n2907 ;
  assign new_n2909 = ~new_n2900 & new_n2908 ;
  assign new_n2910 = ~new_n2896 & new_n2909 ;
  assign new_n2911 = lo0299 & ~lo0300 ;
  assign new_n2912 = new_n2826 & new_n2911 ;
  assign new_n2913 = ~new_n2910 & new_n2912 ;
  assign new_n2914 = ~new_n2829 & ~new_n2913 ;
  assign new_n2915 = ~lo0297 & ~lo0300 ;
  assign new_n2916 = lo0298 & new_n2915 ;
  assign new_n2917 = lo0846 & new_n2916 ;
  assign new_n2918 = ~lo0299 & new_n2917 ;
  assign new_n2919 = ~new_n2619 & new_n2918 ;
  assign new_n2920 = lo0442 & new_n2490 ;
  assign new_n2921 = lo0441 & new_n2493 ;
  assign new_n2922 = ~new_n2492 & ~new_n2921 ;
  assign new_n2923 = ~new_n2920 & new_n2922 ;
  assign new_n2924 = ~lo0249 & ~new_n2923 ;
  assign new_n2925 = lo0249 & new_n2923 ;
  assign new_n2926 = ~new_n2924 & ~new_n2925 ;
  assign new_n2927 = lo0440 & ~new_n2926 ;
  assign new_n2928 = ~lo0440 & new_n2924 ;
  assign new_n2929 = lo0249 & lo0443 ;
  assign new_n2930 = ~new_n2923 & new_n2929 ;
  assign new_n2931 = ~new_n2928 & ~new_n2930 ;
  assign new_n2932 = ~new_n2927 & new_n2931 ;
  assign new_n2933 = lo0450 & new_n2490 ;
  assign new_n2934 = ~lo0250 & lo0449 ;
  assign new_n2935 = lo0249 & new_n2934 ;
  assign new_n2936 = ~new_n2492 & ~new_n2935 ;
  assign new_n2937 = ~new_n2933 & new_n2936 ;
  assign new_n2938 = ~lo0250 & ~new_n2937 ;
  assign new_n2939 = lo0250 & new_n2937 ;
  assign new_n2940 = ~new_n2938 & ~new_n2939 ;
  assign new_n2941 = lo0448 & ~new_n2940 ;
  assign new_n2942 = ~lo0448 & new_n2938 ;
  assign new_n2943 = lo0250 & lo0451 ;
  assign new_n2944 = ~new_n2937 & new_n2943 ;
  assign new_n2945 = ~new_n2942 & ~new_n2944 ;
  assign new_n2946 = ~new_n2941 & new_n2945 ;
  assign new_n2947 = new_n2506 & ~new_n2946 ;
  assign new_n2948 = lo0446 & new_n2490 ;
  assign new_n2949 = ~lo0250 & lo0445 ;
  assign new_n2950 = lo0249 & new_n2949 ;
  assign new_n2951 = ~new_n2492 & ~new_n2950 ;
  assign new_n2952 = ~new_n2948 & new_n2951 ;
  assign new_n2953 = ~lo0250 & ~new_n2952 ;
  assign new_n2954 = lo0250 & new_n2952 ;
  assign new_n2955 = ~new_n2953 & ~new_n2954 ;
  assign new_n2956 = lo0444 & ~new_n2955 ;
  assign new_n2957 = ~lo0444 & new_n2953 ;
  assign new_n2958 = lo0250 & lo0447 ;
  assign new_n2959 = ~new_n2952 & new_n2958 ;
  assign new_n2960 = ~new_n2957 & ~new_n2959 ;
  assign new_n2961 = ~new_n2956 & new_n2960 ;
  assign new_n2962 = new_n2831 & ~new_n2961 ;
  assign new_n2963 = ~new_n2521 & ~new_n2962 ;
  assign new_n2964 = ~new_n2947 & new_n2963 ;
  assign new_n2965 = ~lo0252 & ~new_n2964 ;
  assign new_n2966 = lo0252 & new_n2964 ;
  assign new_n2967 = ~new_n2965 & ~new_n2966 ;
  assign new_n2968 = ~new_n2932 & ~new_n2967 ;
  assign new_n2969 = new_n2932 & new_n2965 ;
  assign new_n2970 = lo0454 & new_n2490 ;
  assign new_n2971 = lo0453 & new_n2493 ;
  assign new_n2972 = ~new_n2492 & ~new_n2971 ;
  assign new_n2973 = ~new_n2970 & new_n2972 ;
  assign new_n2974 = ~lo0249 & ~new_n2973 ;
  assign new_n2975 = lo0249 & new_n2973 ;
  assign new_n2976 = ~new_n2974 & ~new_n2975 ;
  assign new_n2977 = lo0452 & ~new_n2976 ;
  assign new_n2978 = ~lo0452 & new_n2974 ;
  assign new_n2979 = lo0249 & lo0455 ;
  assign new_n2980 = ~new_n2973 & new_n2979 ;
  assign new_n2981 = ~new_n2978 & ~new_n2980 ;
  assign new_n2982 = ~new_n2977 & new_n2981 ;
  assign new_n2983 = lo0252 & ~new_n2982 ;
  assign new_n2984 = ~new_n2964 & new_n2983 ;
  assign new_n2985 = ~new_n2969 & ~new_n2984 ;
  assign new_n2986 = ~new_n2968 & new_n2985 ;
  assign new_n2987 = new_n2489 & ~new_n2986 ;
  assign new_n2988 = lo0091 & lo0456 ;
  assign new_n2989 = ~new_n2715 & ~new_n2988 ;
  assign new_n2990 = lo0090 & ~new_n2989 ;
  assign new_n2991 = ~new_n2483 & new_n2990 ;
  assign new_n2992 = lo0457 & new_n2601 ;
  assign new_n2993 = lo0459 & new_n2605 ;
  assign new_n2994 = ~new_n2992 & ~new_n2993 ;
  assign new_n2995 = lo0458 & new_n2613 ;
  assign new_n2996 = lo1318 & new_n2610 ;
  assign new_n2997 = ~new_n2995 & ~new_n2996 ;
  assign new_n2998 = new_n2994 & new_n2997 ;
  assign new_n2999 = ~new_n2729 & new_n2998 ;
  assign new_n3000 = ~new_n2991 & new_n2999 ;
  assign new_n3001 = ~new_n2987 & new_n3000 ;
  assign new_n3002 = ~lo0299 & ~lo0300 ;
  assign new_n3003 = new_n2826 & new_n3002 ;
  assign new_n3004 = ~new_n3001 & new_n3003 ;
  assign new_n3005 = ~new_n2919 & ~new_n3004 ;
  assign new_n3006 = new_n2914 & new_n3005 ;
  assign new_n3007 = ~new_n2739 & new_n2916 ;
  assign new_n3008 = lo0299 & ~lo0846 ;
  assign new_n3009 = new_n3007 & new_n3008 ;
  assign new_n3010 = ~lo0298 & new_n2915 ;
  assign new_n3011 = lo0481 & new_n2506 ;
  assign new_n3012 = ~lo0252 & lo0480 ;
  assign new_n3013 = lo0251 & new_n3012 ;
  assign new_n3014 = ~new_n2521 & ~new_n3013 ;
  assign new_n3015 = ~new_n3011 & new_n3014 ;
  assign new_n3016 = ~lo0252 & ~new_n3015 ;
  assign new_n3017 = lo0252 & new_n3015 ;
  assign new_n3018 = ~new_n3016 & ~new_n3017 ;
  assign new_n3019 = lo0479 & ~new_n3018 ;
  assign new_n3020 = ~lo0479 & new_n3016 ;
  assign new_n3021 = lo0252 & lo0482 ;
  assign new_n3022 = ~new_n3015 & new_n3021 ;
  assign new_n3023 = ~new_n3020 & ~new_n3022 ;
  assign new_n3024 = ~new_n3019 & new_n3023 ;
  assign new_n3025 = lo0489 & new_n2506 ;
  assign new_n3026 = ~lo0252 & lo0488 ;
  assign new_n3027 = lo0251 & new_n3026 ;
  assign new_n3028 = ~new_n2521 & ~new_n3027 ;
  assign new_n3029 = ~new_n3025 & new_n3028 ;
  assign new_n3030 = ~lo0252 & ~new_n3029 ;
  assign new_n3031 = lo0252 & new_n3029 ;
  assign new_n3032 = ~new_n3030 & ~new_n3031 ;
  assign new_n3033 = lo0487 & ~new_n3032 ;
  assign new_n3034 = ~lo0487 & new_n3030 ;
  assign new_n3035 = lo0252 & lo0490 ;
  assign new_n3036 = ~new_n3029 & new_n3035 ;
  assign new_n3037 = ~new_n3034 & ~new_n3036 ;
  assign new_n3038 = ~new_n3033 & new_n3037 ;
  assign new_n3039 = new_n2490 & ~new_n3038 ;
  assign new_n3040 = lo0485 & new_n2506 ;
  assign new_n3041 = lo0484 & new_n2522 ;
  assign new_n3042 = ~new_n2521 & ~new_n3041 ;
  assign new_n3043 = ~new_n3040 & new_n3042 ;
  assign new_n3044 = ~lo0251 & ~new_n3043 ;
  assign new_n3045 = lo0251 & new_n3043 ;
  assign new_n3046 = ~new_n3044 & ~new_n3045 ;
  assign new_n3047 = lo0483 & ~new_n3046 ;
  assign new_n3048 = ~lo0483 & new_n3044 ;
  assign new_n3049 = lo0251 & lo0486 ;
  assign new_n3050 = ~new_n3043 & new_n3049 ;
  assign new_n3051 = ~new_n3048 & ~new_n3050 ;
  assign new_n3052 = ~new_n3047 & new_n3051 ;
  assign new_n3053 = new_n2493 & ~new_n3052 ;
  assign new_n3054 = ~new_n2492 & ~new_n3053 ;
  assign new_n3055 = ~new_n3039 & new_n3054 ;
  assign new_n3056 = ~lo0249 & ~new_n3055 ;
  assign new_n3057 = lo0249 & new_n3055 ;
  assign new_n3058 = ~new_n3056 & ~new_n3057 ;
  assign new_n3059 = ~new_n3024 & ~new_n3058 ;
  assign new_n3060 = new_n3024 & new_n3056 ;
  assign new_n3061 = lo0493 & new_n2506 ;
  assign new_n3062 = lo0492 & new_n2522 ;
  assign new_n3063 = ~new_n2521 & ~new_n3062 ;
  assign new_n3064 = ~new_n3061 & new_n3063 ;
  assign new_n3065 = ~lo0251 & ~new_n3064 ;
  assign new_n3066 = lo0251 & new_n3064 ;
  assign new_n3067 = ~new_n3065 & ~new_n3066 ;
  assign new_n3068 = lo0491 & ~new_n3067 ;
  assign new_n3069 = ~lo0491 & new_n3065 ;
  assign new_n3070 = lo0251 & lo0494 ;
  assign new_n3071 = ~new_n3064 & new_n3070 ;
  assign new_n3072 = ~new_n3069 & ~new_n3071 ;
  assign new_n3073 = ~new_n3068 & new_n3072 ;
  assign new_n3074 = lo0249 & ~new_n3073 ;
  assign new_n3075 = ~new_n3055 & new_n3074 ;
  assign new_n3076 = ~new_n3060 & ~new_n3075 ;
  assign new_n3077 = ~new_n3059 & new_n3076 ;
  assign new_n3078 = new_n2489 & ~new_n3077 ;
  assign new_n3079 = lo0091 & lo0436 ;
  assign new_n3080 = ~new_n2715 & ~new_n3079 ;
  assign new_n3081 = lo0090 & ~new_n3080 ;
  assign new_n3082 = ~new_n2483 & new_n3081 ;
  assign new_n3083 = lo0495 & new_n2601 ;
  assign new_n3084 = lo0497 & new_n2605 ;
  assign new_n3085 = ~new_n3083 & ~new_n3084 ;
  assign new_n3086 = lo0496 & new_n2613 ;
  assign new_n3087 = lo1320 & new_n2610 ;
  assign new_n3088 = ~new_n3086 & ~new_n3087 ;
  assign new_n3089 = new_n3085 & new_n3088 ;
  assign new_n3090 = ~new_n2729 & new_n3089 ;
  assign new_n3091 = ~new_n3082 & new_n3090 ;
  assign new_n3092 = ~new_n3078 & new_n3091 ;
  assign new_n3093 = new_n3010 & ~new_n3092 ;
  assign new_n3094 = lo0299 & lo0760 ;
  assign new_n3095 = new_n2917 & new_n3094 ;
  assign new_n3096 = ~new_n3093 & ~new_n3095 ;
  assign new_n3097 = ~new_n3009 & new_n3096 ;
  assign new_n3098 = new_n3006 & new_n3097 ;
  assign new_n3099 = lo0196 & lo0197 ;
  assign new_n3100 = lo0199 & ~lo0200 ;
  assign new_n3101 = lo0198 & new_n3100 ;
  assign new_n3102 = new_n3099 & new_n3101 ;
  assign new_n3103 = ~new_n3098 & new_n3102 ;
  assign new_n3104 = ~new_n2739 & ~new_n3102 ;
  assign new_n3105 = ~new_n3103 & ~new_n3104 ;
  assign new_n3106 = lo0110 & lo0826 ;
  assign new_n3107 = ~lo0110 & ~lo0826 ;
  assign new_n3108 = ~new_n3106 & ~new_n3107 ;
  assign new_n3109 = lo0198 & lo0199 ;
  assign new_n3110 = new_n3099 & new_n3109 ;
  assign new_n3111 = ~new_n3108 & new_n3110 ;
  assign new_n3112 = ~lo0200 & ~new_n3111 ;
  assign new_n3113 = lo0196 & ~lo0197 ;
  assign new_n3114 = lo0198 & new_n3113 ;
  assign new_n3115 = lo0199 & new_n3114 ;
  assign new_n3116 = ~lo0196 & lo0197 ;
  assign new_n3117 = ~new_n3113 & ~new_n3116 ;
  assign new_n3118 = ~lo0197 & ~lo0200 ;
  assign new_n3119 = lo0199 & ~new_n3118 ;
  assign new_n3120 = ~new_n3117 & new_n3119 ;
  assign new_n3121 = new_n3115 & ~new_n3120 ;
  assign new_n3122 = ~lo0062 & ~lo0064 ;
  assign new_n3123 = ~lo0058 & ~lo0060 ;
  assign new_n3124 = lo0057 & new_n3123 ;
  assign new_n3125 = new_n3122 & new_n3124 ;
  assign new_n3126 = new_n3121 & new_n3125 ;
  assign new_n3127 = ~lo0198 & new_n3120 ;
  assign new_n3128 = ~new_n3113 & ~new_n3120 ;
  assign new_n3129 = ~new_n3127 & ~new_n3128 ;
  assign new_n3130 = ~new_n3121 & ~new_n3129 ;
  assign new_n3131 = ~new_n3126 & ~new_n3130 ;
  assign new_n3132 = lo0199 & ~new_n3120 ;
  assign new_n3133 = new_n3131 & ~new_n3132 ;
  assign new_n3134 = ~new_n3121 & ~new_n3133 ;
  assign new_n3135 = ~new_n3131 & ~new_n3134 ;
  assign new_n3136 = new_n3131 & new_n3134 ;
  assign new_n3137 = ~new_n3135 & ~new_n3136 ;
  assign new_n3138 = new_n2728 & ~new_n3137 ;
  assign new_n3139 = ~new_n2728 & new_n3135 ;
  assign new_n3140 = ~new_n3138 & ~new_n3139 ;
  assign new_n3141 = ~new_n3131 & new_n3134 ;
  assign new_n3142 = ~lo0062 & lo0063 ;
  assign new_n3143 = ~lo0058 & lo0059 ;
  assign new_n3144 = lo0060 & ~lo0061 ;
  assign new_n3145 = ~new_n3143 & ~new_n3144 ;
  assign new_n3146 = ~new_n3142 & new_n3145 ;
  assign new_n3147 = ~lo0064 & lo0065 ;
  assign new_n3148 = lo0055 & lo0057 ;
  assign new_n3149 = ~new_n3147 & new_n3148 ;
  assign new_n3150 = lo0058 & ~lo0059 ;
  assign new_n3151 = lo0064 & ~lo0065 ;
  assign new_n3152 = ~new_n3150 & ~new_n3151 ;
  assign new_n3153 = ~lo0060 & lo0061 ;
  assign new_n3154 = lo0062 & ~lo0063 ;
  assign new_n3155 = ~new_n3153 & ~new_n3154 ;
  assign new_n3156 = new_n3152 & new_n3155 ;
  assign new_n3157 = new_n3149 & new_n3156 ;
  assign new_n3158 = new_n3146 & new_n3157 ;
  assign new_n3159 = lo0056 & lo0066 ;
  assign new_n3160 = ~new_n3158 & ~new_n3159 ;
  assign new_n3161 = ~lo0070 & ~lo0071 ;
  assign new_n3162 = ~lo0069 & new_n3161 ;
  assign new_n3163 = ~lo0072 & ~lo0073 ;
  assign new_n3164 = ~lo0068 & new_n3163 ;
  assign new_n3165 = new_n3162 & new_n3164 ;
  assign new_n3166 = ~lo0067 & new_n3165 ;
  assign new_n3167 = lo0055 & ~lo0056 ;
  assign new_n3168 = new_n3166 & new_n3167 ;
  assign new_n3169 = new_n3160 & new_n3168 ;
  assign new_n3170 = ~lo0059 & ~lo0061 ;
  assign new_n3171 = lo0462 & new_n3170 ;
  assign new_n3172 = lo0059 & lo0061 ;
  assign new_n3173 = ~lo0059 & lo0061 ;
  assign new_n3174 = lo0461 & new_n3173 ;
  assign new_n3175 = ~new_n3172 & ~new_n3174 ;
  assign new_n3176 = ~new_n3171 & new_n3175 ;
  assign new_n3177 = ~lo0059 & ~new_n3176 ;
  assign new_n3178 = lo0059 & new_n3176 ;
  assign new_n3179 = ~new_n3177 & ~new_n3178 ;
  assign new_n3180 = lo0460 & ~new_n3179 ;
  assign new_n3181 = ~lo0460 & new_n3177 ;
  assign new_n3182 = lo0059 & lo0463 ;
  assign new_n3183 = ~new_n3176 & new_n3182 ;
  assign new_n3184 = ~new_n3181 & ~new_n3183 ;
  assign new_n3185 = ~new_n3180 & new_n3184 ;
  assign new_n3186 = ~lo0063 & ~lo0065 ;
  assign new_n3187 = lo0470 & new_n3170 ;
  assign new_n3188 = lo0469 & new_n3173 ;
  assign new_n3189 = ~new_n3172 & ~new_n3188 ;
  assign new_n3190 = ~new_n3187 & new_n3189 ;
  assign new_n3191 = ~lo0059 & ~new_n3190 ;
  assign new_n3192 = lo0059 & new_n3190 ;
  assign new_n3193 = ~new_n3191 & ~new_n3192 ;
  assign new_n3194 = lo0468 & ~new_n3193 ;
  assign new_n3195 = ~lo0468 & new_n3191 ;
  assign new_n3196 = lo0059 & lo0471 ;
  assign new_n3197 = ~new_n3190 & new_n3196 ;
  assign new_n3198 = ~new_n3195 & ~new_n3197 ;
  assign new_n3199 = ~new_n3194 & new_n3198 ;
  assign new_n3200 = new_n3186 & ~new_n3199 ;
  assign new_n3201 = lo0063 & lo0065 ;
  assign new_n3202 = ~lo0063 & lo0065 ;
  assign new_n3203 = lo0466 & new_n3170 ;
  assign new_n3204 = lo0059 & ~lo0061 ;
  assign new_n3205 = lo0465 & new_n3204 ;
  assign new_n3206 = ~new_n3172 & ~new_n3205 ;
  assign new_n3207 = ~new_n3203 & new_n3206 ;
  assign new_n3208 = ~lo0061 & ~new_n3207 ;
  assign new_n3209 = lo0061 & new_n3207 ;
  assign new_n3210 = ~new_n3208 & ~new_n3209 ;
  assign new_n3211 = lo0464 & ~new_n3210 ;
  assign new_n3212 = ~lo0464 & new_n3208 ;
  assign new_n3213 = lo0061 & lo0467 ;
  assign new_n3214 = ~new_n3207 & new_n3213 ;
  assign new_n3215 = ~new_n3212 & ~new_n3214 ;
  assign new_n3216 = ~new_n3211 & new_n3215 ;
  assign new_n3217 = new_n3202 & ~new_n3216 ;
  assign new_n3218 = ~new_n3201 & ~new_n3217 ;
  assign new_n3219 = ~new_n3200 & new_n3218 ;
  assign new_n3220 = ~lo0063 & ~new_n3219 ;
  assign new_n3221 = lo0063 & new_n3219 ;
  assign new_n3222 = ~new_n3220 & ~new_n3221 ;
  assign new_n3223 = ~new_n3185 & ~new_n3222 ;
  assign new_n3224 = new_n3185 & new_n3220 ;
  assign new_n3225 = lo0474 & new_n3170 ;
  assign new_n3226 = lo0473 & new_n3204 ;
  assign new_n3227 = ~new_n3172 & ~new_n3226 ;
  assign new_n3228 = ~new_n3225 & new_n3227 ;
  assign new_n3229 = ~lo0061 & ~new_n3228 ;
  assign new_n3230 = lo0061 & new_n3228 ;
  assign new_n3231 = ~new_n3229 & ~new_n3230 ;
  assign new_n3232 = lo0472 & ~new_n3231 ;
  assign new_n3233 = ~lo0472 & new_n3229 ;
  assign new_n3234 = lo0061 & lo0475 ;
  assign new_n3235 = ~new_n3228 & new_n3234 ;
  assign new_n3236 = ~new_n3233 & ~new_n3235 ;
  assign new_n3237 = ~new_n3232 & new_n3236 ;
  assign new_n3238 = lo0063 & ~new_n3237 ;
  assign new_n3239 = ~new_n3219 & new_n3238 ;
  assign new_n3240 = ~new_n3224 & ~new_n3239 ;
  assign new_n3241 = ~new_n3223 & new_n3240 ;
  assign new_n3242 = new_n3169 & ~new_n3241 ;
  assign new_n3243 = new_n2718 & ~new_n3160 ;
  assign new_n3244 = ~lo0055 & ~lo0066 ;
  assign new_n3245 = lo0056 & new_n3244 ;
  assign new_n3246 = new_n3166 & new_n3245 ;
  assign new_n3247 = lo1409 & new_n3246 ;
  assign new_n3248 = ~lo0055 & ~lo0056 ;
  assign new_n3249 = ~lo0067 & new_n3248 ;
  assign new_n3250 = ~lo0068 & ~lo0069 ;
  assign new_n3251 = new_n3249 & new_n3250 ;
  assign new_n3252 = new_n3161 & new_n3251 ;
  assign new_n3253 = ~lo0072 & lo0073 ;
  assign new_n3254 = new_n3252 & new_n3253 ;
  assign new_n3255 = lo1319 & new_n3254 ;
  assign new_n3256 = new_n3163 & new_n3251 ;
  assign new_n3257 = ~lo0070 & lo0071 ;
  assign new_n3258 = new_n3256 & new_n3257 ;
  assign new_n3259 = lo0477 & new_n3258 ;
  assign new_n3260 = ~new_n3255 & ~new_n3259 ;
  assign new_n3261 = ~new_n3247 & new_n3260 ;
  assign new_n3262 = new_n3163 & new_n3249 ;
  assign new_n3263 = lo0068 & new_n3162 ;
  assign new_n3264 = new_n3262 & new_n3263 ;
  assign new_n3265 = new_n2728 & new_n3264 ;
  assign new_n3266 = lo0072 & ~lo0073 ;
  assign new_n3267 = new_n3252 & new_n3266 ;
  assign new_n3268 = lo1408 & new_n3267 ;
  assign new_n3269 = lo0067 & new_n3248 ;
  assign new_n3270 = new_n3165 & new_n3269 ;
  assign new_n3271 = lo1410 & new_n3270 ;
  assign new_n3272 = ~lo0068 & lo0069 ;
  assign new_n3273 = new_n3161 & new_n3272 ;
  assign new_n3274 = new_n3262 & new_n3273 ;
  assign new_n3275 = lo0476 & new_n3274 ;
  assign new_n3276 = ~new_n3271 & ~new_n3275 ;
  assign new_n3277 = ~new_n3268 & new_n3276 ;
  assign new_n3278 = ~new_n3265 & new_n3277 ;
  assign new_n3279 = new_n3261 & new_n3278 ;
  assign new_n3280 = ~new_n3243 & new_n3279 ;
  assign new_n3281 = ~new_n3242 & new_n3280 ;
  assign new_n3282 = new_n3141 & ~new_n3281 ;
  assign new_n3283 = new_n3140 & ~new_n3282 ;
  assign new_n3284 = ~new_n3121 & ~new_n3283 ;
  assign new_n3285 = new_n3121 & new_n3283 ;
  assign new_n3286 = ~new_n3284 & ~new_n3285 ;
  assign new_n3287 = lo0470 & ~new_n3286 ;
  assign new_n3288 = ~lo0470 & new_n3284 ;
  assign new_n3289 = new_n2718 & new_n3121 ;
  assign new_n3290 = ~new_n3283 & new_n3289 ;
  assign new_n3291 = ~new_n3288 & ~new_n3290 ;
  assign new_n3292 = ~new_n3287 & new_n3291 ;
  assign new_n3293 = ~new_n3112 & new_n3292 ;
  assign new_n3294 = new_n3112 & ~new_n3292 ;
  assign new_n3295 = ~new_n3293 & ~new_n3294 ;
  assign new_n3296 = lo0421 & new_n2490 ;
  assign new_n3297 = lo0420 & new_n2493 ;
  assign new_n3298 = ~new_n2492 & ~new_n3297 ;
  assign new_n3299 = ~new_n3296 & new_n3298 ;
  assign new_n3300 = ~lo0249 & ~new_n3299 ;
  assign new_n3301 = lo0249 & new_n3299 ;
  assign new_n3302 = ~new_n3300 & ~new_n3301 ;
  assign new_n3303 = lo0419 & ~new_n3302 ;
  assign new_n3304 = ~lo0419 & new_n3300 ;
  assign new_n3305 = lo0249 & lo0422 ;
  assign new_n3306 = ~new_n3299 & new_n3305 ;
  assign new_n3307 = ~new_n3304 & ~new_n3306 ;
  assign new_n3308 = ~new_n3303 & new_n3307 ;
  assign new_n3309 = lo0429 & new_n2490 ;
  assign new_n3310 = lo0249 & ~lo0250 ;
  assign new_n3311 = lo0428 & new_n3310 ;
  assign new_n3312 = ~new_n2492 & ~new_n3311 ;
  assign new_n3313 = ~new_n3309 & new_n3312 ;
  assign new_n3314 = ~lo0250 & ~new_n3313 ;
  assign new_n3315 = lo0250 & new_n3313 ;
  assign new_n3316 = ~new_n3314 & ~new_n3315 ;
  assign new_n3317 = lo0427 & ~new_n3316 ;
  assign new_n3318 = ~lo0427 & new_n3314 ;
  assign new_n3319 = lo0250 & lo0430 ;
  assign new_n3320 = ~new_n3313 & new_n3319 ;
  assign new_n3321 = ~new_n3318 & ~new_n3320 ;
  assign new_n3322 = ~new_n3317 & new_n3321 ;
  assign new_n3323 = new_n2506 & ~new_n3322 ;
  assign new_n3324 = lo0425 & new_n2490 ;
  assign new_n3325 = lo0424 & new_n3310 ;
  assign new_n3326 = ~new_n2492 & ~new_n3325 ;
  assign new_n3327 = ~new_n3324 & new_n3326 ;
  assign new_n3328 = ~lo0250 & ~new_n3327 ;
  assign new_n3329 = lo0250 & new_n3327 ;
  assign new_n3330 = ~new_n3328 & ~new_n3329 ;
  assign new_n3331 = lo0423 & ~new_n3330 ;
  assign new_n3332 = ~lo0423 & new_n3328 ;
  assign new_n3333 = lo0250 & lo0426 ;
  assign new_n3334 = ~new_n3327 & new_n3333 ;
  assign new_n3335 = ~new_n3332 & ~new_n3334 ;
  assign new_n3336 = ~new_n3331 & new_n3335 ;
  assign new_n3337 = new_n2831 & ~new_n3336 ;
  assign new_n3338 = ~new_n2521 & ~new_n3337 ;
  assign new_n3339 = ~new_n3323 & new_n3338 ;
  assign new_n3340 = ~lo0252 & ~new_n3339 ;
  assign new_n3341 = lo0252 & new_n3339 ;
  assign new_n3342 = ~new_n3340 & ~new_n3341 ;
  assign new_n3343 = ~new_n3308 & ~new_n3342 ;
  assign new_n3344 = new_n3308 & new_n3340 ;
  assign new_n3345 = lo0433 & new_n2490 ;
  assign new_n3346 = lo0432 & new_n2493 ;
  assign new_n3347 = ~new_n2492 & ~new_n3346 ;
  assign new_n3348 = ~new_n3345 & new_n3347 ;
  assign new_n3349 = ~lo0249 & ~new_n3348 ;
  assign new_n3350 = lo0249 & new_n3348 ;
  assign new_n3351 = ~new_n3349 & ~new_n3350 ;
  assign new_n3352 = lo0431 & ~new_n3351 ;
  assign new_n3353 = ~lo0431 & new_n3349 ;
  assign new_n3354 = lo0249 & lo0434 ;
  assign new_n3355 = ~new_n3348 & new_n3354 ;
  assign new_n3356 = ~new_n3353 & ~new_n3355 ;
  assign new_n3357 = ~new_n3352 & new_n3356 ;
  assign new_n3358 = lo0252 & ~new_n3357 ;
  assign new_n3359 = ~new_n3339 & new_n3358 ;
  assign new_n3360 = ~new_n3344 & ~new_n3359 ;
  assign new_n3361 = ~new_n3343 & new_n3360 ;
  assign new_n3362 = new_n2489 & ~new_n3361 ;
  assign new_n3363 = lo0092 & lo0093 ;
  assign new_n3364 = ~lo0091 & ~new_n3363 ;
  assign new_n3365 = lo0090 & new_n3364 ;
  assign new_n3366 = new_n2711 & new_n3365 ;
  assign new_n3367 = lo0090 & ~new_n3364 ;
  assign new_n3368 = lo0435 & new_n3367 ;
  assign new_n3369 = lo0093 & new_n3365 ;
  assign new_n3370 = lo0436 & new_n3369 ;
  assign new_n3371 = ~new_n3368 & ~new_n3370 ;
  assign new_n3372 = ~new_n3366 & new_n3371 ;
  assign new_n3373 = ~new_n2483 & ~new_n3372 ;
  assign new_n3374 = lo0437 & new_n2601 ;
  assign new_n3375 = lo0439 & new_n2605 ;
  assign new_n3376 = ~new_n3374 & ~new_n3375 ;
  assign new_n3377 = lo0438 & new_n2613 ;
  assign new_n3378 = lo1317 & new_n2610 ;
  assign new_n3379 = ~new_n3377 & ~new_n3378 ;
  assign new_n3380 = new_n3376 & new_n3379 ;
  assign new_n3381 = ~new_n2729 & new_n3380 ;
  assign new_n3382 = ~new_n3373 & new_n3381 ;
  assign new_n3383 = ~new_n3362 & new_n3382 ;
  assign new_n3384 = lo0299 & ~new_n3383 ;
  assign new_n3385 = lo0280 & new_n2506 ;
  assign new_n3386 = lo0279 & new_n2831 ;
  assign new_n3387 = ~new_n2521 & ~new_n3386 ;
  assign new_n3388 = ~new_n3385 & new_n3387 ;
  assign new_n3389 = ~lo0252 & ~new_n3388 ;
  assign new_n3390 = lo0252 & new_n3388 ;
  assign new_n3391 = ~new_n3389 & ~new_n3390 ;
  assign new_n3392 = lo0278 & ~new_n3391 ;
  assign new_n3393 = ~lo0278 & new_n3389 ;
  assign new_n3394 = lo0252 & lo0281 ;
  assign new_n3395 = ~new_n3388 & new_n3394 ;
  assign new_n3396 = ~new_n3393 & ~new_n3395 ;
  assign new_n3397 = ~new_n3392 & new_n3396 ;
  assign new_n3398 = lo0288 & new_n2506 ;
  assign new_n3399 = lo0287 & new_n2522 ;
  assign new_n3400 = ~new_n2521 & ~new_n3399 ;
  assign new_n3401 = ~new_n3398 & new_n3400 ;
  assign new_n3402 = ~lo0251 & ~new_n3401 ;
  assign new_n3403 = lo0251 & new_n3401 ;
  assign new_n3404 = ~new_n3402 & ~new_n3403 ;
  assign new_n3405 = lo0286 & ~new_n3404 ;
  assign new_n3406 = ~lo0286 & new_n3402 ;
  assign new_n3407 = lo0251 & lo0289 ;
  assign new_n3408 = ~new_n3401 & new_n3407 ;
  assign new_n3409 = ~new_n3406 & ~new_n3408 ;
  assign new_n3410 = ~new_n3405 & new_n3409 ;
  assign new_n3411 = new_n2490 & ~new_n3410 ;
  assign new_n3412 = lo0284 & new_n2506 ;
  assign new_n3413 = lo0283 & new_n2522 ;
  assign new_n3414 = ~new_n2521 & ~new_n3413 ;
  assign new_n3415 = ~new_n3412 & new_n3414 ;
  assign new_n3416 = ~lo0251 & ~new_n3415 ;
  assign new_n3417 = lo0251 & new_n3415 ;
  assign new_n3418 = ~new_n3416 & ~new_n3417 ;
  assign new_n3419 = lo0282 & ~new_n3418 ;
  assign new_n3420 = ~lo0282 & new_n3416 ;
  assign new_n3421 = lo0251 & lo0285 ;
  assign new_n3422 = ~new_n3415 & new_n3421 ;
  assign new_n3423 = ~new_n3420 & ~new_n3422 ;
  assign new_n3424 = ~new_n3419 & new_n3423 ;
  assign new_n3425 = new_n3310 & ~new_n3424 ;
  assign new_n3426 = ~new_n2492 & ~new_n3425 ;
  assign new_n3427 = ~new_n3411 & new_n3426 ;
  assign new_n3428 = ~lo0250 & ~new_n3427 ;
  assign new_n3429 = lo0250 & new_n3427 ;
  assign new_n3430 = ~new_n3428 & ~new_n3429 ;
  assign new_n3431 = ~new_n3397 & ~new_n3430 ;
  assign new_n3432 = new_n3397 & new_n3428 ;
  assign new_n3433 = lo0292 & new_n2506 ;
  assign new_n3434 = lo0291 & new_n2831 ;
  assign new_n3435 = ~new_n2521 & ~new_n3434 ;
  assign new_n3436 = ~new_n3433 & new_n3435 ;
  assign new_n3437 = ~lo0252 & ~new_n3436 ;
  assign new_n3438 = lo0252 & new_n3436 ;
  assign new_n3439 = ~new_n3437 & ~new_n3438 ;
  assign new_n3440 = lo0290 & ~new_n3439 ;
  assign new_n3441 = ~lo0290 & new_n3437 ;
  assign new_n3442 = lo0252 & lo0293 ;
  assign new_n3443 = ~new_n3436 & new_n3442 ;
  assign new_n3444 = ~new_n3441 & ~new_n3443 ;
  assign new_n3445 = ~new_n3440 & new_n3444 ;
  assign new_n3446 = lo0250 & ~new_n3445 ;
  assign new_n3447 = ~new_n3427 & new_n3446 ;
  assign new_n3448 = ~new_n3432 & ~new_n3447 ;
  assign new_n3449 = ~new_n3431 & new_n3448 ;
  assign new_n3450 = new_n2489 & ~new_n3449 ;
  assign new_n3451 = lo0091 & lo0217 ;
  assign new_n3452 = ~new_n2715 & ~new_n3451 ;
  assign new_n3453 = lo0090 & ~new_n3452 ;
  assign new_n3454 = ~new_n2483 & new_n3453 ;
  assign new_n3455 = lo0294 & new_n2601 ;
  assign new_n3456 = lo0296 & new_n2605 ;
  assign new_n3457 = ~new_n3455 & ~new_n3456 ;
  assign new_n3458 = lo0295 & new_n2613 ;
  assign new_n3459 = lo1304 & new_n2610 ;
  assign new_n3460 = ~new_n3458 & ~new_n3459 ;
  assign new_n3461 = new_n3457 & new_n3460 ;
  assign new_n3462 = ~new_n2729 & new_n3461 ;
  assign new_n3463 = ~new_n3454 & new_n3462 ;
  assign new_n3464 = ~new_n3450 & new_n3463 ;
  assign new_n3465 = ~lo0299 & ~new_n3464 ;
  assign new_n3466 = ~new_n3384 & ~new_n3465 ;
  assign new_n3467 = ~lo0300 & new_n2825 ;
  assign new_n3468 = ~new_n3466 & new_n3467 ;
  assign new_n3469 = ~new_n3001 & new_n3010 ;
  assign new_n3470 = lo0260 & new_n2506 ;
  assign new_n3471 = lo0259 & new_n2831 ;
  assign new_n3472 = ~new_n2521 & ~new_n3471 ;
  assign new_n3473 = ~new_n3470 & new_n3472 ;
  assign new_n3474 = ~lo0252 & ~new_n3473 ;
  assign new_n3475 = lo0252 & new_n3473 ;
  assign new_n3476 = ~new_n3474 & ~new_n3475 ;
  assign new_n3477 = lo0258 & ~new_n3476 ;
  assign new_n3478 = ~lo0258 & new_n3474 ;
  assign new_n3479 = lo0252 & lo0261 ;
  assign new_n3480 = ~new_n3473 & new_n3479 ;
  assign new_n3481 = ~new_n3478 & ~new_n3480 ;
  assign new_n3482 = ~new_n3477 & new_n3481 ;
  assign new_n3483 = lo0268 & new_n2506 ;
  assign new_n3484 = lo0267 & new_n2831 ;
  assign new_n3485 = ~new_n2521 & ~new_n3484 ;
  assign new_n3486 = ~new_n3483 & new_n3485 ;
  assign new_n3487 = ~lo0252 & ~new_n3486 ;
  assign new_n3488 = lo0252 & new_n3486 ;
  assign new_n3489 = ~new_n3487 & ~new_n3488 ;
  assign new_n3490 = lo0266 & ~new_n3489 ;
  assign new_n3491 = ~lo0266 & new_n3487 ;
  assign new_n3492 = lo0252 & lo0269 ;
  assign new_n3493 = ~new_n3486 & new_n3492 ;
  assign new_n3494 = ~new_n3491 & ~new_n3493 ;
  assign new_n3495 = ~new_n3490 & new_n3494 ;
  assign new_n3496 = new_n2490 & ~new_n3495 ;
  assign new_n3497 = lo0264 & new_n2506 ;
  assign new_n3498 = lo0263 & new_n2522 ;
  assign new_n3499 = ~new_n2521 & ~new_n3498 ;
  assign new_n3500 = ~new_n3497 & new_n3499 ;
  assign new_n3501 = ~lo0251 & ~new_n3500 ;
  assign new_n3502 = lo0251 & new_n3500 ;
  assign new_n3503 = ~new_n3501 & ~new_n3502 ;
  assign new_n3504 = lo0262 & ~new_n3503 ;
  assign new_n3505 = ~lo0262 & new_n3501 ;
  assign new_n3506 = lo0251 & lo0265 ;
  assign new_n3507 = ~new_n3500 & new_n3506 ;
  assign new_n3508 = ~new_n3505 & ~new_n3507 ;
  assign new_n3509 = ~new_n3504 & new_n3508 ;
  assign new_n3510 = new_n2493 & ~new_n3509 ;
  assign new_n3511 = ~new_n2492 & ~new_n3510 ;
  assign new_n3512 = ~new_n3496 & new_n3511 ;
  assign new_n3513 = ~lo0249 & ~new_n3512 ;
  assign new_n3514 = lo0249 & new_n3512 ;
  assign new_n3515 = ~new_n3513 & ~new_n3514 ;
  assign new_n3516 = ~new_n3482 & ~new_n3515 ;
  assign new_n3517 = new_n3482 & new_n3513 ;
  assign new_n3518 = lo0272 & new_n2506 ;
  assign new_n3519 = lo0271 & new_n2522 ;
  assign new_n3520 = ~new_n2521 & ~new_n3519 ;
  assign new_n3521 = ~new_n3518 & new_n3520 ;
  assign new_n3522 = ~lo0251 & ~new_n3521 ;
  assign new_n3523 = lo0251 & new_n3521 ;
  assign new_n3524 = ~new_n3522 & ~new_n3523 ;
  assign new_n3525 = lo0270 & ~new_n3524 ;
  assign new_n3526 = ~lo0270 & new_n3522 ;
  assign new_n3527 = lo0251 & lo0273 ;
  assign new_n3528 = ~new_n3521 & new_n3527 ;
  assign new_n3529 = ~new_n3526 & ~new_n3528 ;
  assign new_n3530 = ~new_n3525 & new_n3529 ;
  assign new_n3531 = lo0249 & ~new_n3530 ;
  assign new_n3532 = ~new_n3512 & new_n3531 ;
  assign new_n3533 = ~new_n3517 & ~new_n3532 ;
  assign new_n3534 = ~new_n3516 & new_n3533 ;
  assign new_n3535 = new_n2489 & ~new_n3534 ;
  assign new_n3536 = lo0091 & lo0274 ;
  assign new_n3537 = ~new_n2715 & ~new_n3536 ;
  assign new_n3538 = lo0090 & ~new_n3537 ;
  assign new_n3539 = ~new_n2483 & new_n3538 ;
  assign new_n3540 = lo0275 & new_n2601 ;
  assign new_n3541 = lo0277 & new_n2605 ;
  assign new_n3542 = ~new_n3540 & ~new_n3541 ;
  assign new_n3543 = lo0276 & new_n2613 ;
  assign new_n3544 = lo1303 & new_n2610 ;
  assign new_n3545 = ~new_n3543 & ~new_n3544 ;
  assign new_n3546 = new_n3542 & new_n3545 ;
  assign new_n3547 = ~new_n2729 & new_n3546 ;
  assign new_n3548 = ~new_n3539 & new_n3547 ;
  assign new_n3549 = ~new_n3535 & new_n3548 ;
  assign new_n3550 = new_n2825 & new_n2827 ;
  assign new_n3551 = ~new_n3549 & new_n3550 ;
  assign new_n3552 = ~new_n3469 & ~new_n3551 ;
  assign new_n3553 = ~new_n3007 & new_n3552 ;
  assign new_n3554 = ~new_n3468 & new_n3553 ;
  assign new_n3555 = new_n3102 & ~new_n3554 ;
  assign new_n3556 = ~new_n3092 & ~new_n3102 ;
  assign new_n3557 = ~new_n3555 & ~new_n3556 ;
  assign new_n3558 = lo0481 & new_n3186 ;
  assign new_n3559 = lo0063 & ~lo0065 ;
  assign new_n3560 = lo0480 & new_n3559 ;
  assign new_n3561 = ~new_n3201 & ~new_n3560 ;
  assign new_n3562 = ~new_n3558 & new_n3561 ;
  assign new_n3563 = ~lo0065 & ~new_n3562 ;
  assign new_n3564 = lo0065 & new_n3562 ;
  assign new_n3565 = ~new_n3563 & ~new_n3564 ;
  assign new_n3566 = lo0479 & ~new_n3565 ;
  assign new_n3567 = ~lo0479 & new_n3563 ;
  assign new_n3568 = lo0065 & lo0482 ;
  assign new_n3569 = ~new_n3562 & new_n3568 ;
  assign new_n3570 = ~new_n3567 & ~new_n3569 ;
  assign new_n3571 = ~new_n3566 & new_n3570 ;
  assign new_n3572 = lo0489 & new_n3186 ;
  assign new_n3573 = lo0488 & new_n3559 ;
  assign new_n3574 = ~new_n3201 & ~new_n3573 ;
  assign new_n3575 = ~new_n3572 & new_n3574 ;
  assign new_n3576 = ~lo0065 & ~new_n3575 ;
  assign new_n3577 = lo0065 & new_n3575 ;
  assign new_n3578 = ~new_n3576 & ~new_n3577 ;
  assign new_n3579 = lo0487 & ~new_n3578 ;
  assign new_n3580 = ~lo0487 & new_n3576 ;
  assign new_n3581 = lo0065 & lo0490 ;
  assign new_n3582 = ~new_n3575 & new_n3581 ;
  assign new_n3583 = ~new_n3580 & ~new_n3582 ;
  assign new_n3584 = ~new_n3579 & new_n3583 ;
  assign new_n3585 = new_n3170 & ~new_n3584 ;
  assign new_n3586 = lo0485 & new_n3186 ;
  assign new_n3587 = lo0484 & new_n3202 ;
  assign new_n3588 = ~new_n3201 & ~new_n3587 ;
  assign new_n3589 = ~new_n3586 & new_n3588 ;
  assign new_n3590 = ~lo0063 & ~new_n3589 ;
  assign new_n3591 = lo0063 & new_n3589 ;
  assign new_n3592 = ~new_n3590 & ~new_n3591 ;
  assign new_n3593 = lo0483 & ~new_n3592 ;
  assign new_n3594 = ~lo0483 & new_n3590 ;
  assign new_n3595 = lo0063 & lo0486 ;
  assign new_n3596 = ~new_n3589 & new_n3595 ;
  assign new_n3597 = ~new_n3594 & ~new_n3596 ;
  assign new_n3598 = ~new_n3593 & new_n3597 ;
  assign new_n3599 = new_n3173 & ~new_n3598 ;
  assign new_n3600 = ~new_n3172 & ~new_n3599 ;
  assign new_n3601 = ~new_n3585 & new_n3600 ;
  assign new_n3602 = ~lo0059 & ~new_n3601 ;
  assign new_n3603 = lo0059 & new_n3601 ;
  assign new_n3604 = ~new_n3602 & ~new_n3603 ;
  assign new_n3605 = ~new_n3571 & ~new_n3604 ;
  assign new_n3606 = new_n3571 & new_n3602 ;
  assign new_n3607 = lo0493 & new_n3186 ;
  assign new_n3608 = lo0492 & new_n3202 ;
  assign new_n3609 = ~new_n3201 & ~new_n3608 ;
  assign new_n3610 = ~new_n3607 & new_n3609 ;
  assign new_n3611 = ~lo0063 & ~new_n3610 ;
  assign new_n3612 = lo0063 & new_n3610 ;
  assign new_n3613 = ~new_n3611 & ~new_n3612 ;
  assign new_n3614 = lo0491 & ~new_n3613 ;
  assign new_n3615 = ~lo0491 & new_n3611 ;
  assign new_n3616 = lo0063 & lo0494 ;
  assign new_n3617 = ~new_n3610 & new_n3616 ;
  assign new_n3618 = ~new_n3615 & ~new_n3617 ;
  assign new_n3619 = ~new_n3614 & new_n3618 ;
  assign new_n3620 = lo0059 & ~new_n3619 ;
  assign new_n3621 = ~new_n3601 & new_n3620 ;
  assign new_n3622 = ~new_n3606 & ~new_n3621 ;
  assign new_n3623 = ~new_n3605 & new_n3622 ;
  assign new_n3624 = new_n3169 & ~new_n3623 ;
  assign new_n3625 = new_n3081 & ~new_n3160 ;
  assign new_n3626 = lo1331 & new_n3246 ;
  assign new_n3627 = lo1320 & new_n3254 ;
  assign new_n3628 = lo0496 & new_n3258 ;
  assign new_n3629 = ~new_n3627 & ~new_n3628 ;
  assign new_n3630 = ~new_n3626 & new_n3629 ;
  assign new_n3631 = lo1330 & new_n3267 ;
  assign new_n3632 = lo1332 & new_n3270 ;
  assign new_n3633 = lo0495 & new_n3274 ;
  assign new_n3634 = ~new_n3632 & ~new_n3633 ;
  assign new_n3635 = ~new_n3631 & new_n3634 ;
  assign new_n3636 = ~new_n3265 & new_n3635 ;
  assign new_n3637 = new_n3630 & new_n3636 ;
  assign new_n3638 = ~new_n3625 & new_n3637 ;
  assign new_n3639 = ~new_n3624 & new_n3638 ;
  assign new_n3640 = new_n3141 & ~new_n3639 ;
  assign new_n3641 = new_n3140 & ~new_n3640 ;
  assign new_n3642 = ~new_n3121 & ~new_n3641 ;
  assign new_n3643 = new_n3121 & new_n3641 ;
  assign new_n3644 = ~new_n3642 & ~new_n3643 ;
  assign new_n3645 = lo0489 & ~new_n3644 ;
  assign new_n3646 = ~lo0489 & new_n3642 ;
  assign new_n3647 = new_n3081 & new_n3121 ;
  assign new_n3648 = ~new_n3641 & new_n3647 ;
  assign new_n3649 = ~new_n3646 & ~new_n3648 ;
  assign new_n3650 = ~new_n3645 & new_n3649 ;
  assign new_n3651 = ~new_n3112 & new_n3650 ;
  assign new_n3652 = new_n3112 & ~new_n3650 ;
  assign new_n3653 = ~new_n3651 & ~new_n3652 ;
  assign new_n3654 = lo0520 & new_n2506 ;
  assign new_n3655 = lo0519 & new_n2831 ;
  assign new_n3656 = ~new_n2521 & ~new_n3655 ;
  assign new_n3657 = ~new_n3654 & new_n3656 ;
  assign new_n3658 = ~lo0252 & ~new_n3657 ;
  assign new_n3659 = lo0252 & new_n3657 ;
  assign new_n3660 = ~new_n3658 & ~new_n3659 ;
  assign new_n3661 = lo0518 & ~new_n3660 ;
  assign new_n3662 = ~lo0518 & new_n3658 ;
  assign new_n3663 = lo0252 & lo0521 ;
  assign new_n3664 = ~new_n3657 & new_n3663 ;
  assign new_n3665 = ~new_n3662 & ~new_n3664 ;
  assign new_n3666 = ~new_n3661 & new_n3665 ;
  assign new_n3667 = lo0528 & new_n2506 ;
  assign new_n3668 = lo0527 & new_n2522 ;
  assign new_n3669 = ~new_n2521 & ~new_n3668 ;
  assign new_n3670 = ~new_n3667 & new_n3669 ;
  assign new_n3671 = ~lo0251 & ~new_n3670 ;
  assign new_n3672 = lo0251 & new_n3670 ;
  assign new_n3673 = ~new_n3671 & ~new_n3672 ;
  assign new_n3674 = lo0526 & ~new_n3673 ;
  assign new_n3675 = ~lo0526 & new_n3671 ;
  assign new_n3676 = lo0251 & lo0529 ;
  assign new_n3677 = ~new_n3670 & new_n3676 ;
  assign new_n3678 = ~new_n3675 & ~new_n3677 ;
  assign new_n3679 = ~new_n3674 & new_n3678 ;
  assign new_n3680 = new_n2490 & ~new_n3679 ;
  assign new_n3681 = lo0524 & new_n2506 ;
  assign new_n3682 = lo0523 & new_n2522 ;
  assign new_n3683 = ~new_n2521 & ~new_n3682 ;
  assign new_n3684 = ~new_n3681 & new_n3683 ;
  assign new_n3685 = ~lo0251 & ~new_n3684 ;
  assign new_n3686 = lo0251 & new_n3684 ;
  assign new_n3687 = ~new_n3685 & ~new_n3686 ;
  assign new_n3688 = lo0522 & ~new_n3687 ;
  assign new_n3689 = ~lo0522 & new_n3685 ;
  assign new_n3690 = lo0251 & lo0525 ;
  assign new_n3691 = ~new_n3684 & new_n3690 ;
  assign new_n3692 = ~new_n3689 & ~new_n3691 ;
  assign new_n3693 = ~new_n3688 & new_n3692 ;
  assign new_n3694 = new_n3310 & ~new_n3693 ;
  assign new_n3695 = ~new_n2492 & ~new_n3694 ;
  assign new_n3696 = ~new_n3680 & new_n3695 ;
  assign new_n3697 = ~lo0250 & ~new_n3696 ;
  assign new_n3698 = lo0250 & new_n3696 ;
  assign new_n3699 = ~new_n3697 & ~new_n3698 ;
  assign new_n3700 = ~new_n3666 & ~new_n3699 ;
  assign new_n3701 = new_n3666 & new_n3697 ;
  assign new_n3702 = lo0532 & new_n2506 ;
  assign new_n3703 = lo0531 & new_n2831 ;
  assign new_n3704 = ~new_n2521 & ~new_n3703 ;
  assign new_n3705 = ~new_n3702 & new_n3704 ;
  assign new_n3706 = ~lo0252 & ~new_n3705 ;
  assign new_n3707 = lo0252 & new_n3705 ;
  assign new_n3708 = ~new_n3706 & ~new_n3707 ;
  assign new_n3709 = lo0530 & ~new_n3708 ;
  assign new_n3710 = ~lo0530 & new_n3706 ;
  assign new_n3711 = lo0252 & lo0533 ;
  assign new_n3712 = ~new_n3705 & new_n3711 ;
  assign new_n3713 = ~new_n3710 & ~new_n3712 ;
  assign new_n3714 = ~new_n3709 & new_n3713 ;
  assign new_n3715 = lo0250 & ~new_n3714 ;
  assign new_n3716 = ~new_n3696 & new_n3715 ;
  assign new_n3717 = ~new_n3701 & ~new_n3716 ;
  assign new_n3718 = ~new_n3700 & new_n3717 ;
  assign new_n3719 = new_n2489 & ~new_n3718 ;
  assign new_n3720 = lo0534 & new_n3367 ;
  assign new_n3721 = lo0456 & new_n3369 ;
  assign new_n3722 = ~new_n3720 & ~new_n3721 ;
  assign new_n3723 = ~new_n3366 & new_n3722 ;
  assign new_n3724 = ~new_n2483 & ~new_n3723 ;
  assign new_n3725 = lo0535 & new_n2601 ;
  assign new_n3726 = lo0537 & new_n2605 ;
  assign new_n3727 = ~new_n3725 & ~new_n3726 ;
  assign new_n3728 = lo0536 & new_n2613 ;
  assign new_n3729 = lo1328 & new_n2610 ;
  assign new_n3730 = ~new_n3728 & ~new_n3729 ;
  assign new_n3731 = new_n3727 & new_n3730 ;
  assign new_n3732 = ~new_n2729 & new_n3731 ;
  assign new_n3733 = ~new_n3724 & new_n3732 ;
  assign new_n3734 = ~new_n3719 & new_n3733 ;
  assign new_n3735 = lo0297 & ~new_n3002 ;
  assign new_n3736 = lo0297 & ~lo0300 ;
  assign new_n3737 = ~new_n3735 & new_n3736 ;
  assign new_n3738 = lo0647 & new_n2490 ;
  assign new_n3739 = lo0646 & new_n2493 ;
  assign new_n3740 = ~new_n2492 & ~new_n3739 ;
  assign new_n3741 = ~new_n3738 & new_n3740 ;
  assign new_n3742 = ~lo0249 & ~new_n3741 ;
  assign new_n3743 = lo0249 & new_n3741 ;
  assign new_n3744 = ~new_n3742 & ~new_n3743 ;
  assign new_n3745 = lo0645 & ~new_n3744 ;
  assign new_n3746 = ~lo0645 & new_n3742 ;
  assign new_n3747 = lo0249 & lo0648 ;
  assign new_n3748 = ~new_n3741 & new_n3747 ;
  assign new_n3749 = ~new_n3746 & ~new_n3748 ;
  assign new_n3750 = ~new_n3745 & new_n3749 ;
  assign new_n3751 = lo0655 & new_n2490 ;
  assign new_n3752 = lo0654 & new_n2493 ;
  assign new_n3753 = ~new_n2492 & ~new_n3752 ;
  assign new_n3754 = ~new_n3751 & new_n3753 ;
  assign new_n3755 = ~lo0249 & ~new_n3754 ;
  assign new_n3756 = lo0249 & new_n3754 ;
  assign new_n3757 = ~new_n3755 & ~new_n3756 ;
  assign new_n3758 = lo0653 & ~new_n3757 ;
  assign new_n3759 = ~lo0653 & new_n3755 ;
  assign new_n3760 = lo0249 & lo0656 ;
  assign new_n3761 = ~new_n3754 & new_n3760 ;
  assign new_n3762 = ~new_n3759 & ~new_n3761 ;
  assign new_n3763 = ~new_n3758 & new_n3762 ;
  assign new_n3764 = new_n2506 & ~new_n3763 ;
  assign new_n3765 = lo0651 & new_n2490 ;
  assign new_n3766 = lo0650 & new_n3310 ;
  assign new_n3767 = ~new_n2492 & ~new_n3766 ;
  assign new_n3768 = ~new_n3765 & new_n3767 ;
  assign new_n3769 = ~lo0250 & ~new_n3768 ;
  assign new_n3770 = lo0250 & new_n3768 ;
  assign new_n3771 = ~new_n3769 & ~new_n3770 ;
  assign new_n3772 = lo0649 & ~new_n3771 ;
  assign new_n3773 = ~lo0649 & new_n3769 ;
  assign new_n3774 = lo0250 & lo0652 ;
  assign new_n3775 = ~new_n3768 & new_n3774 ;
  assign new_n3776 = ~new_n3773 & ~new_n3775 ;
  assign new_n3777 = ~new_n3772 & new_n3776 ;
  assign new_n3778 = new_n2522 & ~new_n3777 ;
  assign new_n3779 = ~new_n2521 & ~new_n3778 ;
  assign new_n3780 = ~new_n3764 & new_n3779 ;
  assign new_n3781 = ~lo0251 & ~new_n3780 ;
  assign new_n3782 = lo0251 & new_n3780 ;
  assign new_n3783 = ~new_n3781 & ~new_n3782 ;
  assign new_n3784 = ~new_n3750 & ~new_n3783 ;
  assign new_n3785 = new_n3750 & new_n3781 ;
  assign new_n3786 = lo0659 & new_n2490 ;
  assign new_n3787 = lo0658 & new_n3310 ;
  assign new_n3788 = ~new_n2492 & ~new_n3787 ;
  assign new_n3789 = ~new_n3786 & new_n3788 ;
  assign new_n3790 = ~lo0250 & ~new_n3789 ;
  assign new_n3791 = lo0250 & new_n3789 ;
  assign new_n3792 = ~new_n3790 & ~new_n3791 ;
  assign new_n3793 = lo0657 & ~new_n3792 ;
  assign new_n3794 = ~lo0657 & new_n3790 ;
  assign new_n3795 = lo0250 & lo0660 ;
  assign new_n3796 = ~new_n3789 & new_n3795 ;
  assign new_n3797 = ~new_n3794 & ~new_n3796 ;
  assign new_n3798 = ~new_n3793 & new_n3797 ;
  assign new_n3799 = lo0251 & ~new_n3798 ;
  assign new_n3800 = ~new_n3780 & new_n3799 ;
  assign new_n3801 = ~new_n3785 & ~new_n3800 ;
  assign new_n3802 = ~new_n3784 & new_n3801 ;
  assign new_n3803 = new_n2489 & ~new_n3802 ;
  assign new_n3804 = lo0091 & lo0576 ;
  assign new_n3805 = ~new_n2715 & ~new_n3804 ;
  assign new_n3806 = lo0090 & ~new_n3805 ;
  assign new_n3807 = ~new_n2483 & new_n3806 ;
  assign new_n3808 = lo0661 & new_n2601 ;
  assign new_n3809 = lo0663 & new_n2605 ;
  assign new_n3810 = ~new_n3808 & ~new_n3809 ;
  assign new_n3811 = lo0662 & new_n2613 ;
  assign new_n3812 = lo1349 & new_n2610 ;
  assign new_n3813 = ~new_n3811 & ~new_n3812 ;
  assign new_n3814 = new_n3810 & new_n3813 ;
  assign new_n3815 = ~new_n2729 & new_n3814 ;
  assign new_n3816 = ~new_n3807 & new_n3815 ;
  assign new_n3817 = ~new_n3803 & new_n3816 ;
  assign new_n3818 = new_n3737 & ~new_n3817 ;
  assign new_n3819 = new_n3735 & ~new_n3736 ;
  assign new_n3820 = ~new_n3735 & ~new_n3736 ;
  assign new_n3821 = ~new_n3464 & new_n3820 ;
  assign new_n3822 = ~new_n3819 & ~new_n3821 ;
  assign new_n3823 = ~new_n3818 & new_n3822 ;
  assign new_n3824 = ~new_n3735 & ~new_n3823 ;
  assign new_n3825 = new_n3735 & new_n3823 ;
  assign new_n3826 = ~new_n3824 & ~new_n3825 ;
  assign new_n3827 = ~new_n3734 & ~new_n3826 ;
  assign new_n3828 = new_n3734 & new_n3824 ;
  assign new_n3829 = lo0363 & new_n2490 ;
  assign new_n3830 = lo0362 & new_n2493 ;
  assign new_n3831 = ~new_n2492 & ~new_n3830 ;
  assign new_n3832 = ~new_n3829 & new_n3831 ;
  assign new_n3833 = ~lo0249 & ~new_n3832 ;
  assign new_n3834 = lo0249 & new_n3832 ;
  assign new_n3835 = ~new_n3833 & ~new_n3834 ;
  assign new_n3836 = lo0361 & ~new_n3835 ;
  assign new_n3837 = ~lo0361 & new_n3833 ;
  assign new_n3838 = lo0249 & lo0364 ;
  assign new_n3839 = ~new_n3832 & new_n3838 ;
  assign new_n3840 = ~new_n3837 & ~new_n3839 ;
  assign new_n3841 = ~new_n3836 & new_n3840 ;
  assign new_n3842 = lo0371 & new_n2490 ;
  assign new_n3843 = lo0370 & new_n3310 ;
  assign new_n3844 = ~new_n2492 & ~new_n3843 ;
  assign new_n3845 = ~new_n3842 & new_n3844 ;
  assign new_n3846 = ~lo0250 & ~new_n3845 ;
  assign new_n3847 = lo0250 & new_n3845 ;
  assign new_n3848 = ~new_n3846 & ~new_n3847 ;
  assign new_n3849 = lo0369 & ~new_n3848 ;
  assign new_n3850 = ~lo0369 & new_n3846 ;
  assign new_n3851 = lo0250 & lo0372 ;
  assign new_n3852 = ~new_n3845 & new_n3851 ;
  assign new_n3853 = ~new_n3850 & ~new_n3852 ;
  assign new_n3854 = ~new_n3849 & new_n3853 ;
  assign new_n3855 = new_n2506 & ~new_n3854 ;
  assign new_n3856 = lo0367 & new_n2490 ;
  assign new_n3857 = lo0366 & new_n3310 ;
  assign new_n3858 = ~new_n2492 & ~new_n3857 ;
  assign new_n3859 = ~new_n3856 & new_n3858 ;
  assign new_n3860 = ~lo0250 & ~new_n3859 ;
  assign new_n3861 = lo0250 & new_n3859 ;
  assign new_n3862 = ~new_n3860 & ~new_n3861 ;
  assign new_n3863 = lo0365 & ~new_n3862 ;
  assign new_n3864 = ~lo0365 & new_n3860 ;
  assign new_n3865 = lo0250 & lo0368 ;
  assign new_n3866 = ~new_n3859 & new_n3865 ;
  assign new_n3867 = ~new_n3864 & ~new_n3866 ;
  assign new_n3868 = ~new_n3863 & new_n3867 ;
  assign new_n3869 = new_n2831 & ~new_n3868 ;
  assign new_n3870 = ~new_n2521 & ~new_n3869 ;
  assign new_n3871 = ~new_n3855 & new_n3870 ;
  assign new_n3872 = ~lo0252 & ~new_n3871 ;
  assign new_n3873 = lo0252 & new_n3871 ;
  assign new_n3874 = ~new_n3872 & ~new_n3873 ;
  assign new_n3875 = ~new_n3841 & ~new_n3874 ;
  assign new_n3876 = new_n3841 & new_n3872 ;
  assign new_n3877 = lo0375 & new_n2490 ;
  assign new_n3878 = lo0374 & new_n2493 ;
  assign new_n3879 = ~new_n2492 & ~new_n3878 ;
  assign new_n3880 = ~new_n3877 & new_n3879 ;
  assign new_n3881 = ~lo0249 & ~new_n3880 ;
  assign new_n3882 = lo0249 & new_n3880 ;
  assign new_n3883 = ~new_n3881 & ~new_n3882 ;
  assign new_n3884 = lo0373 & ~new_n3883 ;
  assign new_n3885 = ~lo0373 & new_n3881 ;
  assign new_n3886 = lo0249 & lo0376 ;
  assign new_n3887 = ~new_n3880 & new_n3886 ;
  assign new_n3888 = ~new_n3885 & ~new_n3887 ;
  assign new_n3889 = ~new_n3884 & new_n3888 ;
  assign new_n3890 = lo0252 & ~new_n3889 ;
  assign new_n3891 = ~new_n3871 & new_n3890 ;
  assign new_n3892 = ~new_n3876 & ~new_n3891 ;
  assign new_n3893 = ~new_n3875 & new_n3892 ;
  assign new_n3894 = new_n2489 & ~new_n3893 ;
  assign new_n3895 = lo0091 & lo0377 ;
  assign new_n3896 = ~new_n2715 & ~new_n3895 ;
  assign new_n3897 = lo0090 & ~new_n3896 ;
  assign new_n3898 = ~new_n2483 & new_n3897 ;
  assign new_n3899 = lo0378 & new_n2601 ;
  assign new_n3900 = lo0380 & new_n2605 ;
  assign new_n3901 = ~new_n3899 & ~new_n3900 ;
  assign new_n3902 = lo0379 & new_n2613 ;
  assign new_n3903 = lo1308 & new_n2610 ;
  assign new_n3904 = ~new_n3902 & ~new_n3903 ;
  assign new_n3905 = new_n3901 & new_n3904 ;
  assign new_n3906 = ~new_n2729 & new_n3905 ;
  assign new_n3907 = ~new_n3898 & new_n3906 ;
  assign new_n3908 = ~new_n3894 & new_n3907 ;
  assign new_n3909 = new_n3735 & ~new_n3908 ;
  assign new_n3910 = ~new_n3823 & new_n3909 ;
  assign new_n3911 = ~new_n3828 & ~new_n3910 ;
  assign new_n3912 = ~new_n3827 & new_n3911 ;
  assign new_n3913 = ~lo0298 & ~new_n3912 ;
  assign new_n3914 = lo0297 & new_n3002 ;
  assign new_n3915 = ~new_n2739 & new_n3914 ;
  assign new_n3916 = ~lo0297 & ~new_n3092 ;
  assign new_n3917 = ~new_n3915 & ~new_n3916 ;
  assign new_n3918 = lo0298 & ~new_n3917 ;
  assign new_n3919 = ~new_n3913 & ~new_n3918 ;
  assign new_n3920 = new_n3102 & ~new_n3919 ;
  assign new_n3921 = ~new_n3001 & ~new_n3102 ;
  assign new_n3922 = ~new_n3920 & ~new_n3921 ;
  assign new_n3923 = lo0442 & new_n3170 ;
  assign new_n3924 = lo0441 & new_n3173 ;
  assign new_n3925 = ~new_n3172 & ~new_n3924 ;
  assign new_n3926 = ~new_n3923 & new_n3925 ;
  assign new_n3927 = ~lo0059 & ~new_n3926 ;
  assign new_n3928 = lo0059 & new_n3926 ;
  assign new_n3929 = ~new_n3927 & ~new_n3928 ;
  assign new_n3930 = lo0440 & ~new_n3929 ;
  assign new_n3931 = ~lo0440 & new_n3927 ;
  assign new_n3932 = lo0059 & lo0443 ;
  assign new_n3933 = ~new_n3926 & new_n3932 ;
  assign new_n3934 = ~new_n3931 & ~new_n3933 ;
  assign new_n3935 = ~new_n3930 & new_n3934 ;
  assign new_n3936 = lo0450 & new_n3170 ;
  assign new_n3937 = lo0449 & new_n3204 ;
  assign new_n3938 = ~new_n3172 & ~new_n3937 ;
  assign new_n3939 = ~new_n3936 & new_n3938 ;
  assign new_n3940 = ~lo0061 & ~new_n3939 ;
  assign new_n3941 = lo0061 & new_n3939 ;
  assign new_n3942 = ~new_n3940 & ~new_n3941 ;
  assign new_n3943 = lo0448 & ~new_n3942 ;
  assign new_n3944 = ~lo0448 & new_n3940 ;
  assign new_n3945 = lo0061 & lo0451 ;
  assign new_n3946 = ~new_n3939 & new_n3945 ;
  assign new_n3947 = ~new_n3944 & ~new_n3946 ;
  assign new_n3948 = ~new_n3943 & new_n3947 ;
  assign new_n3949 = new_n3186 & ~new_n3948 ;
  assign new_n3950 = lo0446 & new_n3170 ;
  assign new_n3951 = lo0445 & new_n3204 ;
  assign new_n3952 = ~new_n3172 & ~new_n3951 ;
  assign new_n3953 = ~new_n3950 & new_n3952 ;
  assign new_n3954 = ~lo0061 & ~new_n3953 ;
  assign new_n3955 = lo0061 & new_n3953 ;
  assign new_n3956 = ~new_n3954 & ~new_n3955 ;
  assign new_n3957 = lo0444 & ~new_n3956 ;
  assign new_n3958 = ~lo0444 & new_n3954 ;
  assign new_n3959 = lo0061 & lo0447 ;
  assign new_n3960 = ~new_n3953 & new_n3959 ;
  assign new_n3961 = ~new_n3958 & ~new_n3960 ;
  assign new_n3962 = ~new_n3957 & new_n3961 ;
  assign new_n3963 = new_n3559 & ~new_n3962 ;
  assign new_n3964 = ~new_n3201 & ~new_n3963 ;
  assign new_n3965 = ~new_n3949 & new_n3964 ;
  assign new_n3966 = ~lo0065 & ~new_n3965 ;
  assign new_n3967 = lo0065 & new_n3965 ;
  assign new_n3968 = ~new_n3966 & ~new_n3967 ;
  assign new_n3969 = ~new_n3935 & ~new_n3968 ;
  assign new_n3970 = new_n3935 & new_n3966 ;
  assign new_n3971 = lo0454 & new_n3170 ;
  assign new_n3972 = lo0453 & new_n3173 ;
  assign new_n3973 = ~new_n3172 & ~new_n3972 ;
  assign new_n3974 = ~new_n3971 & new_n3973 ;
  assign new_n3975 = ~lo0059 & ~new_n3974 ;
  assign new_n3976 = lo0059 & new_n3974 ;
  assign new_n3977 = ~new_n3975 & ~new_n3976 ;
  assign new_n3978 = lo0452 & ~new_n3977 ;
  assign new_n3979 = ~lo0452 & new_n3975 ;
  assign new_n3980 = lo0059 & lo0455 ;
  assign new_n3981 = ~new_n3974 & new_n3980 ;
  assign new_n3982 = ~new_n3979 & ~new_n3981 ;
  assign new_n3983 = ~new_n3978 & new_n3982 ;
  assign new_n3984 = lo0065 & ~new_n3983 ;
  assign new_n3985 = ~new_n3965 & new_n3984 ;
  assign new_n3986 = ~new_n3970 & ~new_n3985 ;
  assign new_n3987 = ~new_n3969 & new_n3986 ;
  assign new_n3988 = new_n3169 & ~new_n3987 ;
  assign new_n3989 = new_n2990 & ~new_n3160 ;
  assign new_n3990 = lo1406 & new_n3246 ;
  assign new_n3991 = lo1318 & new_n3254 ;
  assign new_n3992 = lo0458 & new_n3258 ;
  assign new_n3993 = ~new_n3991 & ~new_n3992 ;
  assign new_n3994 = ~new_n3990 & new_n3993 ;
  assign new_n3995 = lo1405 & new_n3267 ;
  assign new_n3996 = lo1407 & new_n3270 ;
  assign new_n3997 = lo0457 & new_n3274 ;
  assign new_n3998 = ~new_n3996 & ~new_n3997 ;
  assign new_n3999 = ~new_n3995 & new_n3998 ;
  assign new_n4000 = ~new_n3265 & new_n3999 ;
  assign new_n4001 = new_n3994 & new_n4000 ;
  assign new_n4002 = ~new_n3989 & new_n4001 ;
  assign new_n4003 = ~new_n3988 & new_n4002 ;
  assign new_n4004 = new_n3141 & ~new_n4003 ;
  assign new_n4005 = new_n3140 & ~new_n4004 ;
  assign new_n4006 = ~new_n3121 & ~new_n4005 ;
  assign new_n4007 = new_n3121 & new_n4005 ;
  assign new_n4008 = ~new_n4006 & ~new_n4007 ;
  assign new_n4009 = lo0450 & ~new_n4008 ;
  assign new_n4010 = ~lo0450 & new_n4006 ;
  assign new_n4011 = new_n2990 & new_n3121 ;
  assign new_n4012 = ~new_n4005 & new_n4011 ;
  assign new_n4013 = ~new_n4010 & ~new_n4012 ;
  assign new_n4014 = ~new_n4009 & new_n4013 ;
  assign new_n4015 = ~new_n3112 & new_n4014 ;
  assign new_n4016 = new_n3112 & ~new_n4014 ;
  assign new_n4017 = ~new_n4015 & ~new_n4016 ;
  assign new_n4018 = lo0666 & new_n2506 ;
  assign new_n4019 = lo0665 & new_n2831 ;
  assign new_n4020 = ~new_n2521 & ~new_n4019 ;
  assign new_n4021 = ~new_n4018 & new_n4020 ;
  assign new_n4022 = ~lo0252 & ~new_n4021 ;
  assign new_n4023 = lo0252 & new_n4021 ;
  assign new_n4024 = ~new_n4022 & ~new_n4023 ;
  assign new_n4025 = lo0664 & ~new_n4024 ;
  assign new_n4026 = ~lo0664 & new_n4022 ;
  assign new_n4027 = lo0252 & lo0667 ;
  assign new_n4028 = ~new_n4021 & new_n4027 ;
  assign new_n4029 = ~new_n4026 & ~new_n4028 ;
  assign new_n4030 = ~new_n4025 & new_n4029 ;
  assign new_n4031 = lo0674 & new_n2506 ;
  assign new_n4032 = lo0673 & new_n2831 ;
  assign new_n4033 = ~new_n2521 & ~new_n4032 ;
  assign new_n4034 = ~new_n4031 & new_n4033 ;
  assign new_n4035 = ~lo0252 & ~new_n4034 ;
  assign new_n4036 = lo0252 & new_n4034 ;
  assign new_n4037 = ~new_n4035 & ~new_n4036 ;
  assign new_n4038 = lo0672 & ~new_n4037 ;
  assign new_n4039 = ~lo0672 & new_n4035 ;
  assign new_n4040 = lo0252 & lo0675 ;
  assign new_n4041 = ~new_n4034 & new_n4040 ;
  assign new_n4042 = ~new_n4039 & ~new_n4041 ;
  assign new_n4043 = ~new_n4038 & new_n4042 ;
  assign new_n4044 = new_n2490 & ~new_n4043 ;
  assign new_n4045 = lo0670 & new_n2506 ;
  assign new_n4046 = lo0669 & new_n2522 ;
  assign new_n4047 = ~new_n2521 & ~new_n4046 ;
  assign new_n4048 = ~new_n4045 & new_n4047 ;
  assign new_n4049 = ~lo0251 & ~new_n4048 ;
  assign new_n4050 = lo0251 & new_n4048 ;
  assign new_n4051 = ~new_n4049 & ~new_n4050 ;
  assign new_n4052 = lo0668 & ~new_n4051 ;
  assign new_n4053 = ~lo0668 & new_n4049 ;
  assign new_n4054 = lo0251 & lo0671 ;
  assign new_n4055 = ~new_n4048 & new_n4054 ;
  assign new_n4056 = ~new_n4053 & ~new_n4055 ;
  assign new_n4057 = ~new_n4052 & new_n4056 ;
  assign new_n4058 = new_n2493 & ~new_n4057 ;
  assign new_n4059 = ~new_n2492 & ~new_n4058 ;
  assign new_n4060 = ~new_n4044 & new_n4059 ;
  assign new_n4061 = ~lo0249 & ~new_n4060 ;
  assign new_n4062 = lo0249 & new_n4060 ;
  assign new_n4063 = ~new_n4061 & ~new_n4062 ;
  assign new_n4064 = ~new_n4030 & ~new_n4063 ;
  assign new_n4065 = new_n4030 & new_n4061 ;
  assign new_n4066 = lo0678 & new_n2506 ;
  assign new_n4067 = lo0677 & new_n2522 ;
  assign new_n4068 = ~new_n2521 & ~new_n4067 ;
  assign new_n4069 = ~new_n4066 & new_n4068 ;
  assign new_n4070 = ~lo0251 & ~new_n4069 ;
  assign new_n4071 = lo0251 & new_n4069 ;
  assign new_n4072 = ~new_n4070 & ~new_n4071 ;
  assign new_n4073 = lo0676 & ~new_n4072 ;
  assign new_n4074 = ~lo0676 & new_n4070 ;
  assign new_n4075 = lo0251 & lo0679 ;
  assign new_n4076 = ~new_n4069 & new_n4075 ;
  assign new_n4077 = ~new_n4074 & ~new_n4076 ;
  assign new_n4078 = ~new_n4073 & new_n4077 ;
  assign new_n4079 = lo0249 & ~new_n4078 ;
  assign new_n4080 = ~new_n4060 & new_n4079 ;
  assign new_n4081 = ~new_n4065 & ~new_n4080 ;
  assign new_n4082 = ~new_n4064 & new_n4081 ;
  assign new_n4083 = new_n2489 & ~new_n4082 ;
  assign new_n4084 = lo0091 & lo0638 ;
  assign new_n4085 = ~new_n2715 & ~new_n4084 ;
  assign new_n4086 = lo0090 & ~new_n4085 ;
  assign new_n4087 = ~new_n2483 & new_n4086 ;
  assign new_n4088 = lo0680 & new_n2601 ;
  assign new_n4089 = lo0682 & new_n2605 ;
  assign new_n4090 = ~new_n4088 & ~new_n4089 ;
  assign new_n4091 = lo0681 & new_n2613 ;
  assign new_n4092 = lo1350 & new_n2610 ;
  assign new_n4093 = ~new_n4091 & ~new_n4092 ;
  assign new_n4094 = new_n4090 & new_n4093 ;
  assign new_n4095 = ~new_n2729 & new_n4094 ;
  assign new_n4096 = ~new_n4087 & new_n4095 ;
  assign new_n4097 = ~new_n4083 & new_n4096 ;
  assign new_n4098 = new_n3737 & ~new_n4097 ;
  assign new_n4099 = lo0344 & new_n2490 ;
  assign new_n4100 = lo0343 & new_n2493 ;
  assign new_n4101 = ~new_n2492 & ~new_n4100 ;
  assign new_n4102 = ~new_n4099 & new_n4101 ;
  assign new_n4103 = ~lo0249 & ~new_n4102 ;
  assign new_n4104 = lo0249 & new_n4102 ;
  assign new_n4105 = ~new_n4103 & ~new_n4104 ;
  assign new_n4106 = lo0342 & ~new_n4105 ;
  assign new_n4107 = ~lo0342 & new_n4103 ;
  assign new_n4108 = lo0249 & lo0345 ;
  assign new_n4109 = ~new_n4102 & new_n4108 ;
  assign new_n4110 = ~new_n4107 & ~new_n4109 ;
  assign new_n4111 = ~new_n4106 & new_n4110 ;
  assign new_n4112 = lo1307 & new_n2490 ;
  assign new_n4113 = lo0351 & new_n2493 ;
  assign new_n4114 = ~new_n2492 & ~new_n4113 ;
  assign new_n4115 = ~new_n4112 & new_n4114 ;
  assign new_n4116 = ~lo0249 & ~new_n4115 ;
  assign new_n4117 = lo0249 & new_n4115 ;
  assign new_n4118 = ~new_n4116 & ~new_n4117 ;
  assign new_n4119 = lo0350 & ~new_n4118 ;
  assign new_n4120 = ~lo0350 & new_n4116 ;
  assign new_n4121 = lo0249 & lo0352 ;
  assign new_n4122 = ~new_n4115 & new_n4121 ;
  assign new_n4123 = ~new_n4120 & ~new_n4122 ;
  assign new_n4124 = ~new_n4119 & new_n4123 ;
  assign new_n4125 = new_n2506 & ~new_n4124 ;
  assign new_n4126 = lo0348 & new_n2490 ;
  assign new_n4127 = lo0347 & new_n3310 ;
  assign new_n4128 = ~new_n2492 & ~new_n4127 ;
  assign new_n4129 = ~new_n4126 & new_n4128 ;
  assign new_n4130 = ~lo0250 & ~new_n4129 ;
  assign new_n4131 = lo0250 & new_n4129 ;
  assign new_n4132 = ~new_n4130 & ~new_n4131 ;
  assign new_n4133 = lo0346 & ~new_n4132 ;
  assign new_n4134 = ~lo0346 & new_n4130 ;
  assign new_n4135 = lo0250 & lo0349 ;
  assign new_n4136 = ~new_n4129 & new_n4135 ;
  assign new_n4137 = ~new_n4134 & ~new_n4136 ;
  assign new_n4138 = ~new_n4133 & new_n4137 ;
  assign new_n4139 = new_n2522 & ~new_n4138 ;
  assign new_n4140 = ~new_n2521 & ~new_n4139 ;
  assign new_n4141 = ~new_n4125 & new_n4140 ;
  assign new_n4142 = ~lo0251 & ~new_n4141 ;
  assign new_n4143 = lo0251 & new_n4141 ;
  assign new_n4144 = ~new_n4142 & ~new_n4143 ;
  assign new_n4145 = ~new_n4111 & ~new_n4144 ;
  assign new_n4146 = new_n4111 & new_n4142 ;
  assign new_n4147 = lo0355 & new_n2490 ;
  assign new_n4148 = lo0354 & new_n3310 ;
  assign new_n4149 = ~new_n2492 & ~new_n4148 ;
  assign new_n4150 = ~new_n4147 & new_n4149 ;
  assign new_n4151 = ~lo0250 & ~new_n4150 ;
  assign new_n4152 = lo0250 & new_n4150 ;
  assign new_n4153 = ~new_n4151 & ~new_n4152 ;
  assign new_n4154 = lo0353 & ~new_n4153 ;
  assign new_n4155 = ~lo0353 & new_n4151 ;
  assign new_n4156 = lo0250 & lo0356 ;
  assign new_n4157 = ~new_n4150 & new_n4156 ;
  assign new_n4158 = ~new_n4155 & ~new_n4157 ;
  assign new_n4159 = ~new_n4154 & new_n4158 ;
  assign new_n4160 = lo0251 & ~new_n4159 ;
  assign new_n4161 = ~new_n4141 & new_n4160 ;
  assign new_n4162 = ~new_n4146 & ~new_n4161 ;
  assign new_n4163 = ~new_n4145 & new_n4162 ;
  assign new_n4164 = new_n2489 & ~new_n4163 ;
  assign new_n4165 = lo0219 & new_n3367 ;
  assign new_n4166 = lo0217 & new_n3369 ;
  assign new_n4167 = ~new_n4165 & ~new_n4166 ;
  assign new_n4168 = ~new_n3366 & new_n4167 ;
  assign new_n4169 = ~new_n2483 & ~new_n4168 ;
  assign new_n4170 = lo0357 & new_n2601 ;
  assign new_n4171 = lo0359 & new_n2605 ;
  assign new_n4172 = ~new_n4170 & ~new_n4171 ;
  assign new_n4173 = lo0358 & new_n2613 ;
  assign new_n4174 = lo0360 & new_n2610 ;
  assign new_n4175 = ~new_n4173 & ~new_n4174 ;
  assign new_n4176 = new_n4172 & new_n4175 ;
  assign new_n4177 = ~new_n2729 & new_n4176 ;
  assign new_n4178 = ~new_n4169 & new_n4177 ;
  assign new_n4179 = ~new_n4164 & new_n4178 ;
  assign new_n4180 = new_n3735 & new_n3736 ;
  assign new_n4181 = ~new_n4179 & new_n4180 ;
  assign new_n4182 = ~new_n3819 & ~new_n4181 ;
  assign new_n4183 = ~new_n4098 & new_n4182 ;
  assign new_n4184 = new_n3736 & ~new_n4183 ;
  assign new_n4185 = ~new_n3736 & new_n4183 ;
  assign new_n4186 = ~new_n4184 & ~new_n4185 ;
  assign new_n4187 = ~new_n3817 & ~new_n4186 ;
  assign new_n4188 = new_n3817 & new_n4184 ;
  assign new_n4189 = lo0232 & new_n2506 ;
  assign new_n4190 = lo0231 & new_n2831 ;
  assign new_n4191 = ~new_n2521 & ~new_n4190 ;
  assign new_n4192 = ~new_n4189 & new_n4191 ;
  assign new_n4193 = ~lo0252 & ~new_n4192 ;
  assign new_n4194 = lo0252 & new_n4192 ;
  assign new_n4195 = ~new_n4193 & ~new_n4194 ;
  assign new_n4196 = lo0230 & ~new_n4195 ;
  assign new_n4197 = ~lo0230 & new_n4193 ;
  assign new_n4198 = lo0233 & lo0252 ;
  assign new_n4199 = ~new_n4192 & new_n4198 ;
  assign new_n4200 = ~new_n4197 & ~new_n4199 ;
  assign new_n4201 = ~new_n4196 & new_n4200 ;
  assign new_n4202 = lo0227 & new_n2506 ;
  assign new_n4203 = lo0239 & new_n2522 ;
  assign new_n4204 = ~new_n2521 & ~new_n4203 ;
  assign new_n4205 = ~new_n4202 & new_n4204 ;
  assign new_n4206 = ~lo0251 & ~new_n4205 ;
  assign new_n4207 = lo0251 & new_n4205 ;
  assign new_n4208 = ~new_n4206 & ~new_n4207 ;
  assign new_n4209 = lo0238 & ~new_n4208 ;
  assign new_n4210 = ~lo0238 & new_n4206 ;
  assign new_n4211 = lo0240 & lo0251 ;
  assign new_n4212 = ~new_n4205 & new_n4211 ;
  assign new_n4213 = ~new_n4210 & ~new_n4212 ;
  assign new_n4214 = ~new_n4209 & new_n4213 ;
  assign new_n4215 = new_n2490 & ~new_n4214 ;
  assign new_n4216 = lo0236 & new_n2506 ;
  assign new_n4217 = lo0235 & new_n2522 ;
  assign new_n4218 = ~new_n2521 & ~new_n4217 ;
  assign new_n4219 = ~new_n4216 & new_n4218 ;
  assign new_n4220 = ~lo0251 & ~new_n4219 ;
  assign new_n4221 = lo0251 & new_n4219 ;
  assign new_n4222 = ~new_n4220 & ~new_n4221 ;
  assign new_n4223 = lo0234 & ~new_n4222 ;
  assign new_n4224 = ~lo0234 & new_n4220 ;
  assign new_n4225 = lo0237 & lo0251 ;
  assign new_n4226 = ~new_n4219 & new_n4225 ;
  assign new_n4227 = ~new_n4224 & ~new_n4226 ;
  assign new_n4228 = ~new_n4223 & new_n4227 ;
  assign new_n4229 = new_n3310 & ~new_n4228 ;
  assign new_n4230 = ~new_n2492 & ~new_n4229 ;
  assign new_n4231 = ~new_n4215 & new_n4230 ;
  assign new_n4232 = ~lo0250 & ~new_n4231 ;
  assign new_n4233 = lo0250 & new_n4231 ;
  assign new_n4234 = ~new_n4232 & ~new_n4233 ;
  assign new_n4235 = ~new_n4201 & ~new_n4234 ;
  assign new_n4236 = new_n4201 & new_n4232 ;
  assign new_n4237 = lo0243 & new_n2506 ;
  assign new_n4238 = lo0242 & new_n2831 ;
  assign new_n4239 = ~new_n2521 & ~new_n4238 ;
  assign new_n4240 = ~new_n4237 & new_n4239 ;
  assign new_n4241 = ~lo0252 & ~new_n4240 ;
  assign new_n4242 = lo0252 & new_n4240 ;
  assign new_n4243 = ~new_n4241 & ~new_n4242 ;
  assign new_n4244 = lo0241 & ~new_n4243 ;
  assign new_n4245 = ~lo0241 & new_n4241 ;
  assign new_n4246 = lo0244 & lo0252 ;
  assign new_n4247 = ~new_n4240 & new_n4246 ;
  assign new_n4248 = ~new_n4245 & ~new_n4247 ;
  assign new_n4249 = ~new_n4244 & new_n4248 ;
  assign new_n4250 = lo0250 & ~new_n4249 ;
  assign new_n4251 = ~new_n4231 & new_n4250 ;
  assign new_n4252 = ~new_n4236 & ~new_n4251 ;
  assign new_n4253 = ~new_n4235 & new_n4252 ;
  assign new_n4254 = new_n2489 & ~new_n4253 ;
  assign new_n4255 = lo0091 & lo0218 ;
  assign new_n4256 = ~new_n2715 & ~new_n4255 ;
  assign new_n4257 = lo0090 & ~new_n4256 ;
  assign new_n4258 = ~new_n2483 & new_n4257 ;
  assign new_n4259 = lo0245 & new_n2601 ;
  assign new_n4260 = lo0381 & new_n2605 ;
  assign new_n4261 = ~new_n4259 & ~new_n4260 ;
  assign new_n4262 = lo0246 & new_n2613 ;
  assign new_n4263 = lo1300 & new_n2610 ;
  assign new_n4264 = ~new_n4262 & ~new_n4263 ;
  assign new_n4265 = new_n4261 & new_n4264 ;
  assign new_n4266 = ~new_n2729 & new_n4265 ;
  assign new_n4267 = ~new_n4258 & new_n4266 ;
  assign new_n4268 = ~new_n4254 & new_n4267 ;
  assign new_n4269 = ~new_n3736 & ~new_n4268 ;
  assign new_n4270 = ~new_n4183 & new_n4269 ;
  assign new_n4271 = ~new_n4188 & ~new_n4270 ;
  assign new_n4272 = ~new_n4187 & new_n4271 ;
  assign new_n4273 = ~lo0298 & ~new_n4272 ;
  assign new_n4274 = ~new_n3092 & new_n3914 ;
  assign new_n4275 = ~lo0297 & ~new_n3001 ;
  assign new_n4276 = ~new_n4274 & ~new_n4275 ;
  assign new_n4277 = lo0298 & ~new_n4276 ;
  assign new_n4278 = ~new_n4273 & ~new_n4277 ;
  assign new_n4279 = new_n3102 & ~new_n4278 ;
  assign new_n4280 = ~new_n3102 & ~new_n3464 ;
  assign new_n4281 = ~new_n4279 & ~new_n4280 ;
  assign new_n4282 = lo0280 & new_n3186 ;
  assign new_n4283 = lo0279 & new_n3559 ;
  assign new_n4284 = ~new_n3201 & ~new_n4283 ;
  assign new_n4285 = ~new_n4282 & new_n4284 ;
  assign new_n4286 = ~lo0065 & ~new_n4285 ;
  assign new_n4287 = lo0065 & new_n4285 ;
  assign new_n4288 = ~new_n4286 & ~new_n4287 ;
  assign new_n4289 = lo0278 & ~new_n4288 ;
  assign new_n4290 = ~lo0278 & new_n4286 ;
  assign new_n4291 = lo0065 & lo0281 ;
  assign new_n4292 = ~new_n4285 & new_n4291 ;
  assign new_n4293 = ~new_n4290 & ~new_n4292 ;
  assign new_n4294 = ~new_n4289 & new_n4293 ;
  assign new_n4295 = lo0288 & new_n3186 ;
  assign new_n4296 = lo0287 & new_n3202 ;
  assign new_n4297 = ~new_n3201 & ~new_n4296 ;
  assign new_n4298 = ~new_n4295 & new_n4297 ;
  assign new_n4299 = ~lo0063 & ~new_n4298 ;
  assign new_n4300 = lo0063 & new_n4298 ;
  assign new_n4301 = ~new_n4299 & ~new_n4300 ;
  assign new_n4302 = lo0286 & ~new_n4301 ;
  assign new_n4303 = ~lo0286 & new_n4299 ;
  assign new_n4304 = lo0063 & lo0289 ;
  assign new_n4305 = ~new_n4298 & new_n4304 ;
  assign new_n4306 = ~new_n4303 & ~new_n4305 ;
  assign new_n4307 = ~new_n4302 & new_n4306 ;
  assign new_n4308 = new_n3170 & ~new_n4307 ;
  assign new_n4309 = lo0284 & new_n3186 ;
  assign new_n4310 = lo0283 & new_n3202 ;
  assign new_n4311 = ~new_n3201 & ~new_n4310 ;
  assign new_n4312 = ~new_n4309 & new_n4311 ;
  assign new_n4313 = ~lo0063 & ~new_n4312 ;
  assign new_n4314 = lo0063 & new_n4312 ;
  assign new_n4315 = ~new_n4313 & ~new_n4314 ;
  assign new_n4316 = lo0282 & ~new_n4315 ;
  assign new_n4317 = ~lo0282 & new_n4313 ;
  assign new_n4318 = lo0063 & lo0285 ;
  assign new_n4319 = ~new_n4312 & new_n4318 ;
  assign new_n4320 = ~new_n4317 & ~new_n4319 ;
  assign new_n4321 = ~new_n4316 & new_n4320 ;
  assign new_n4322 = new_n3204 & ~new_n4321 ;
  assign new_n4323 = ~new_n3172 & ~new_n4322 ;
  assign new_n4324 = ~new_n4308 & new_n4323 ;
  assign new_n4325 = ~lo0061 & ~new_n4324 ;
  assign new_n4326 = lo0061 & new_n4324 ;
  assign new_n4327 = ~new_n4325 & ~new_n4326 ;
  assign new_n4328 = ~new_n4294 & ~new_n4327 ;
  assign new_n4329 = new_n4294 & new_n4325 ;
  assign new_n4330 = lo0292 & new_n3186 ;
  assign new_n4331 = lo0291 & new_n3559 ;
  assign new_n4332 = ~new_n3201 & ~new_n4331 ;
  assign new_n4333 = ~new_n4330 & new_n4332 ;
  assign new_n4334 = ~lo0065 & ~new_n4333 ;
  assign new_n4335 = lo0065 & new_n4333 ;
  assign new_n4336 = ~new_n4334 & ~new_n4335 ;
  assign new_n4337 = lo0290 & ~new_n4336 ;
  assign new_n4338 = ~lo0290 & new_n4334 ;
  assign new_n4339 = lo0065 & lo0293 ;
  assign new_n4340 = ~new_n4333 & new_n4339 ;
  assign new_n4341 = ~new_n4338 & ~new_n4340 ;
  assign new_n4342 = ~new_n4337 & new_n4341 ;
  assign new_n4343 = lo0061 & ~new_n4342 ;
  assign new_n4344 = ~new_n4324 & new_n4343 ;
  assign new_n4345 = ~new_n4329 & ~new_n4344 ;
  assign new_n4346 = ~new_n4328 & new_n4345 ;
  assign new_n4347 = new_n3169 & ~new_n4346 ;
  assign new_n4348 = ~new_n3160 & new_n3453 ;
  assign new_n4349 = lo1354 & new_n3246 ;
  assign new_n4350 = lo1304 & new_n3254 ;
  assign new_n4351 = lo0295 & new_n3258 ;
  assign new_n4352 = ~new_n4350 & ~new_n4351 ;
  assign new_n4353 = ~new_n4349 & new_n4352 ;
  assign new_n4354 = lo1353 & new_n3267 ;
  assign new_n4355 = lo1355 & new_n3270 ;
  assign new_n4356 = lo0294 & new_n3274 ;
  assign new_n4357 = ~new_n4355 & ~new_n4356 ;
  assign new_n4358 = ~new_n4354 & new_n4357 ;
  assign new_n4359 = ~new_n3265 & new_n4358 ;
  assign new_n4360 = new_n4353 & new_n4359 ;
  assign new_n4361 = ~new_n4348 & new_n4360 ;
  assign new_n4362 = ~new_n4347 & new_n4361 ;
  assign new_n4363 = new_n3141 & ~new_n4362 ;
  assign new_n4364 = new_n3140 & ~new_n4363 ;
  assign new_n4365 = ~new_n3121 & ~new_n4364 ;
  assign new_n4366 = new_n3121 & new_n4364 ;
  assign new_n4367 = ~new_n4365 & ~new_n4366 ;
  assign new_n4368 = lo0288 & ~new_n4367 ;
  assign new_n4369 = ~lo0288 & new_n4365 ;
  assign new_n4370 = new_n3121 & new_n3453 ;
  assign new_n4371 = ~new_n4364 & new_n4370 ;
  assign new_n4372 = ~new_n4369 & ~new_n4371 ;
  assign new_n4373 = ~new_n4368 & new_n4372 ;
  assign new_n4374 = ~new_n3112 & new_n4373 ;
  assign new_n4375 = new_n3112 & ~new_n4373 ;
  assign new_n4376 = ~new_n4374 & ~new_n4375 ;
  assign new_n4377 = lo0705 & new_n2506 ;
  assign new_n4378 = lo0704 & new_n2831 ;
  assign new_n4379 = ~new_n2521 & ~new_n4378 ;
  assign new_n4380 = ~new_n4377 & new_n4379 ;
  assign new_n4381 = ~lo0252 & ~new_n4380 ;
  assign new_n4382 = lo0252 & new_n4380 ;
  assign new_n4383 = ~new_n4381 & ~new_n4382 ;
  assign new_n4384 = lo0703 & ~new_n4383 ;
  assign new_n4385 = ~lo0703 & new_n4381 ;
  assign new_n4386 = lo0252 & lo0706 ;
  assign new_n4387 = ~new_n4380 & new_n4386 ;
  assign new_n4388 = ~new_n4385 & ~new_n4387 ;
  assign new_n4389 = ~new_n4384 & new_n4388 ;
  assign new_n4390 = lo0713 & new_n2506 ;
  assign new_n4391 = lo0712 & new_n2831 ;
  assign new_n4392 = ~new_n2521 & ~new_n4391 ;
  assign new_n4393 = ~new_n4390 & new_n4392 ;
  assign new_n4394 = ~lo0252 & ~new_n4393 ;
  assign new_n4395 = lo0252 & new_n4393 ;
  assign new_n4396 = ~new_n4394 & ~new_n4395 ;
  assign new_n4397 = lo0711 & ~new_n4396 ;
  assign new_n4398 = ~lo0711 & new_n4394 ;
  assign new_n4399 = lo0252 & lo0714 ;
  assign new_n4400 = ~new_n4393 & new_n4399 ;
  assign new_n4401 = ~new_n4398 & ~new_n4400 ;
  assign new_n4402 = ~new_n4397 & new_n4401 ;
  assign new_n4403 = new_n2490 & ~new_n4402 ;
  assign new_n4404 = lo0709 & new_n2506 ;
  assign new_n4405 = lo0708 & new_n2522 ;
  assign new_n4406 = ~new_n2521 & ~new_n4405 ;
  assign new_n4407 = ~new_n4404 & new_n4406 ;
  assign new_n4408 = ~lo0251 & ~new_n4407 ;
  assign new_n4409 = lo0251 & new_n4407 ;
  assign new_n4410 = ~new_n4408 & ~new_n4409 ;
  assign new_n4411 = lo0707 & ~new_n4410 ;
  assign new_n4412 = ~lo0707 & new_n4408 ;
  assign new_n4413 = lo0251 & lo0710 ;
  assign new_n4414 = ~new_n4407 & new_n4413 ;
  assign new_n4415 = ~new_n4412 & ~new_n4414 ;
  assign new_n4416 = ~new_n4411 & new_n4415 ;
  assign new_n4417 = new_n2493 & ~new_n4416 ;
  assign new_n4418 = ~new_n2492 & ~new_n4417 ;
  assign new_n4419 = ~new_n4403 & new_n4418 ;
  assign new_n4420 = ~lo0249 & ~new_n4419 ;
  assign new_n4421 = lo0249 & new_n4419 ;
  assign new_n4422 = ~new_n4420 & ~new_n4421 ;
  assign new_n4423 = ~new_n4389 & ~new_n4422 ;
  assign new_n4424 = new_n4389 & new_n4420 ;
  assign new_n4425 = lo0717 & new_n2506 ;
  assign new_n4426 = lo0716 & new_n2522 ;
  assign new_n4427 = ~new_n2521 & ~new_n4426 ;
  assign new_n4428 = ~new_n4425 & new_n4427 ;
  assign new_n4429 = ~lo0251 & ~new_n4428 ;
  assign new_n4430 = lo0251 & new_n4428 ;
  assign new_n4431 = ~new_n4429 & ~new_n4430 ;
  assign new_n4432 = lo0715 & ~new_n4431 ;
  assign new_n4433 = ~lo0715 & new_n4429 ;
  assign new_n4434 = lo0251 & lo0718 ;
  assign new_n4435 = ~new_n4428 & new_n4434 ;
  assign new_n4436 = ~new_n4433 & ~new_n4435 ;
  assign new_n4437 = ~new_n4432 & new_n4436 ;
  assign new_n4438 = lo0249 & ~new_n4437 ;
  assign new_n4439 = ~new_n4419 & new_n4438 ;
  assign new_n4440 = ~new_n4424 & ~new_n4439 ;
  assign new_n4441 = ~new_n4423 & new_n4440 ;
  assign new_n4442 = new_n2489 & ~new_n4441 ;
  assign new_n4443 = lo0577 & new_n3367 ;
  assign new_n4444 = lo0576 & new_n3369 ;
  assign new_n4445 = ~new_n4443 & ~new_n4444 ;
  assign new_n4446 = ~new_n3366 & new_n4445 ;
  assign new_n4447 = ~new_n2483 & ~new_n4446 ;
  assign new_n4448 = lo0719 & new_n2720 ;
  assign new_n4449 = ~new_n2721 & ~new_n4448 ;
  assign new_n4450 = new_n2727 & ~new_n4449 ;
  assign new_n4451 = new_n2591 & new_n4450 ;
  assign new_n4452 = lo0720 & new_n2601 ;
  assign new_n4453 = lo0721 & new_n2605 ;
  assign new_n4454 = ~new_n4452 & ~new_n4453 ;
  assign new_n4455 = lo1352 & new_n2610 ;
  assign new_n4456 = lo0722 & new_n2613 ;
  assign new_n4457 = ~new_n4455 & ~new_n4456 ;
  assign new_n4458 = new_n4454 & new_n4457 ;
  assign new_n4459 = ~new_n4451 & new_n4458 ;
  assign new_n4460 = ~new_n4447 & new_n4459 ;
  assign new_n4461 = ~new_n4442 & new_n4460 ;
  assign new_n4462 = lo0829 & new_n2490 ;
  assign new_n4463 = lo0828 & new_n2493 ;
  assign new_n4464 = ~new_n2492 & ~new_n4463 ;
  assign new_n4465 = ~new_n4462 & new_n4464 ;
  assign new_n4466 = ~lo0249 & ~new_n4465 ;
  assign new_n4467 = lo0249 & new_n4465 ;
  assign new_n4468 = ~new_n4466 & ~new_n4467 ;
  assign new_n4469 = lo0827 & ~new_n4468 ;
  assign new_n4470 = ~lo0827 & new_n4466 ;
  assign new_n4471 = lo0249 & lo0830 ;
  assign new_n4472 = ~new_n4465 & new_n4471 ;
  assign new_n4473 = ~new_n4470 & ~new_n4472 ;
  assign new_n4474 = ~new_n4469 & new_n4473 ;
  assign new_n4475 = lo0837 & new_n2490 ;
  assign new_n4476 = lo0836 & new_n3310 ;
  assign new_n4477 = ~new_n2492 & ~new_n4476 ;
  assign new_n4478 = ~new_n4475 & new_n4477 ;
  assign new_n4479 = ~lo0250 & ~new_n4478 ;
  assign new_n4480 = lo0250 & new_n4478 ;
  assign new_n4481 = ~new_n4479 & ~new_n4480 ;
  assign new_n4482 = lo0835 & ~new_n4481 ;
  assign new_n4483 = ~lo0835 & new_n4479 ;
  assign new_n4484 = lo0250 & lo0838 ;
  assign new_n4485 = ~new_n4478 & new_n4484 ;
  assign new_n4486 = ~new_n4483 & ~new_n4485 ;
  assign new_n4487 = ~new_n4482 & new_n4486 ;
  assign new_n4488 = new_n2506 & ~new_n4487 ;
  assign new_n4489 = lo0833 & new_n2490 ;
  assign new_n4490 = lo0832 & new_n3310 ;
  assign new_n4491 = ~new_n2492 & ~new_n4490 ;
  assign new_n4492 = ~new_n4489 & new_n4491 ;
  assign new_n4493 = ~lo0250 & ~new_n4492 ;
  assign new_n4494 = lo0250 & new_n4492 ;
  assign new_n4495 = ~new_n4493 & ~new_n4494 ;
  assign new_n4496 = lo0831 & ~new_n4495 ;
  assign new_n4497 = ~lo0831 & new_n4493 ;
  assign new_n4498 = lo0250 & lo0834 ;
  assign new_n4499 = ~new_n4492 & new_n4498 ;
  assign new_n4500 = ~new_n4497 & ~new_n4499 ;
  assign new_n4501 = ~new_n4496 & new_n4500 ;
  assign new_n4502 = new_n2831 & ~new_n4501 ;
  assign new_n4503 = ~new_n2521 & ~new_n4502 ;
  assign new_n4504 = ~new_n4488 & new_n4503 ;
  assign new_n4505 = ~lo0252 & ~new_n4504 ;
  assign new_n4506 = lo0252 & new_n4504 ;
  assign new_n4507 = ~new_n4505 & ~new_n4506 ;
  assign new_n4508 = ~new_n4474 & ~new_n4507 ;
  assign new_n4509 = new_n4474 & new_n4505 ;
  assign new_n4510 = lo0841 & new_n2490 ;
  assign new_n4511 = lo0840 & new_n2493 ;
  assign new_n4512 = ~new_n2492 & ~new_n4511 ;
  assign new_n4513 = ~new_n4510 & new_n4512 ;
  assign new_n4514 = ~lo0249 & ~new_n4513 ;
  assign new_n4515 = lo0249 & new_n4513 ;
  assign new_n4516 = ~new_n4514 & ~new_n4515 ;
  assign new_n4517 = lo0839 & ~new_n4516 ;
  assign new_n4518 = ~lo0839 & new_n4514 ;
  assign new_n4519 = lo0249 & lo0842 ;
  assign new_n4520 = ~new_n4513 & new_n4519 ;
  assign new_n4521 = ~new_n4518 & ~new_n4520 ;
  assign new_n4522 = ~new_n4517 & new_n4521 ;
  assign new_n4523 = lo0252 & ~new_n4522 ;
  assign new_n4524 = ~new_n4504 & new_n4523 ;
  assign new_n4525 = ~new_n4509 & ~new_n4524 ;
  assign new_n4526 = ~new_n4508 & new_n4525 ;
  assign new_n4527 = new_n2489 & ~new_n4526 ;
  assign new_n4528 = lo0091 & lo0800 ;
  assign new_n4529 = ~new_n2715 & ~new_n4528 ;
  assign new_n4530 = lo0090 & ~new_n4529 ;
  assign new_n4531 = ~new_n2483 & new_n4530 ;
  assign new_n4532 = lo0843 & new_n2601 ;
  assign new_n4533 = lo0845 & new_n2605 ;
  assign new_n4534 = ~new_n4532 & ~new_n4533 ;
  assign new_n4535 = lo0844 & new_n2613 ;
  assign new_n4536 = lo1392 & new_n2610 ;
  assign new_n4537 = ~new_n4535 & ~new_n4536 ;
  assign new_n4538 = new_n4534 & new_n4537 ;
  assign new_n4539 = ~new_n2729 & new_n4538 ;
  assign new_n4540 = ~new_n4531 & new_n4539 ;
  assign new_n4541 = ~new_n4527 & new_n4540 ;
  assign new_n4542 = new_n3737 & ~new_n4541 ;
  assign new_n4543 = new_n3820 & ~new_n4097 ;
  assign new_n4544 = ~new_n3819 & ~new_n4543 ;
  assign new_n4545 = ~new_n4542 & new_n4544 ;
  assign new_n4546 = ~new_n3735 & ~new_n4545 ;
  assign new_n4547 = new_n3735 & new_n4545 ;
  assign new_n4548 = ~new_n4546 & ~new_n4547 ;
  assign new_n4549 = ~new_n4461 & ~new_n4548 ;
  assign new_n4550 = new_n4461 & new_n4546 ;
  assign new_n4551 = lo0303 & new_n2490 ;
  assign new_n4552 = lo0302 & new_n2493 ;
  assign new_n4553 = ~new_n2492 & ~new_n4552 ;
  assign new_n4554 = ~new_n4551 & new_n4553 ;
  assign new_n4555 = ~lo0249 & ~new_n4554 ;
  assign new_n4556 = lo0249 & new_n4554 ;
  assign new_n4557 = ~new_n4555 & ~new_n4556 ;
  assign new_n4558 = lo0301 & ~new_n4557 ;
  assign new_n4559 = ~lo0301 & new_n4555 ;
  assign new_n4560 = lo0249 & lo0304 ;
  assign new_n4561 = ~new_n4554 & new_n4560 ;
  assign new_n4562 = ~new_n4559 & ~new_n4561 ;
  assign new_n4563 = ~new_n4558 & new_n4562 ;
  assign new_n4564 = lo0311 & new_n2490 ;
  assign new_n4565 = lo0310 & new_n2493 ;
  assign new_n4566 = ~new_n2492 & ~new_n4565 ;
  assign new_n4567 = ~new_n4564 & new_n4566 ;
  assign new_n4568 = ~lo0249 & ~new_n4567 ;
  assign new_n4569 = lo0249 & new_n4567 ;
  assign new_n4570 = ~new_n4568 & ~new_n4569 ;
  assign new_n4571 = lo0309 & ~new_n4570 ;
  assign new_n4572 = ~lo0309 & new_n4568 ;
  assign new_n4573 = lo0249 & lo0312 ;
  assign new_n4574 = ~new_n4567 & new_n4573 ;
  assign new_n4575 = ~new_n4572 & ~new_n4574 ;
  assign new_n4576 = ~new_n4571 & new_n4575 ;
  assign new_n4577 = new_n2506 & ~new_n4576 ;
  assign new_n4578 = lo0307 & new_n2490 ;
  assign new_n4579 = lo0306 & new_n3310 ;
  assign new_n4580 = ~new_n2492 & ~new_n4579 ;
  assign new_n4581 = ~new_n4578 & new_n4580 ;
  assign new_n4582 = ~lo0250 & ~new_n4581 ;
  assign new_n4583 = lo0250 & new_n4581 ;
  assign new_n4584 = ~new_n4582 & ~new_n4583 ;
  assign new_n4585 = lo0305 & ~new_n4584 ;
  assign new_n4586 = ~lo0305 & new_n4582 ;
  assign new_n4587 = lo0250 & lo0308 ;
  assign new_n4588 = ~new_n4581 & new_n4587 ;
  assign new_n4589 = ~new_n4586 & ~new_n4588 ;
  assign new_n4590 = ~new_n4585 & new_n4589 ;
  assign new_n4591 = new_n2522 & ~new_n4590 ;
  assign new_n4592 = ~new_n2521 & ~new_n4591 ;
  assign new_n4593 = ~new_n4577 & new_n4592 ;
  assign new_n4594 = ~lo0251 & ~new_n4593 ;
  assign new_n4595 = lo0251 & new_n4593 ;
  assign new_n4596 = ~new_n4594 & ~new_n4595 ;
  assign new_n4597 = ~new_n4563 & ~new_n4596 ;
  assign new_n4598 = new_n4563 & new_n4594 ;
  assign new_n4599 = lo0315 & new_n2490 ;
  assign new_n4600 = lo0314 & new_n3310 ;
  assign new_n4601 = ~new_n2492 & ~new_n4600 ;
  assign new_n4602 = ~new_n4599 & new_n4601 ;
  assign new_n4603 = ~lo0250 & ~new_n4602 ;
  assign new_n4604 = lo0250 & new_n4602 ;
  assign new_n4605 = ~new_n4603 & ~new_n4604 ;
  assign new_n4606 = lo0313 & ~new_n4605 ;
  assign new_n4607 = ~lo0313 & new_n4603 ;
  assign new_n4608 = lo0250 & lo0316 ;
  assign new_n4609 = ~new_n4602 & new_n4608 ;
  assign new_n4610 = ~new_n4607 & ~new_n4609 ;
  assign new_n4611 = ~new_n4606 & new_n4610 ;
  assign new_n4612 = lo0251 & ~new_n4611 ;
  assign new_n4613 = ~new_n4593 & new_n4612 ;
  assign new_n4614 = ~new_n4598 & ~new_n4613 ;
  assign new_n4615 = ~new_n4597 & new_n4614 ;
  assign new_n4616 = new_n2489 & ~new_n4615 ;
  assign new_n4617 = lo0091 & lo0317 ;
  assign new_n4618 = ~new_n2715 & ~new_n4617 ;
  assign new_n4619 = lo0090 & ~new_n4618 ;
  assign new_n4620 = ~new_n2483 & new_n4619 ;
  assign new_n4621 = lo0318 & new_n2601 ;
  assign new_n4622 = lo0320 & new_n2605 ;
  assign new_n4623 = ~new_n4621 & ~new_n4622 ;
  assign new_n4624 = lo0319 & new_n2613 ;
  assign new_n4625 = lo1305 & new_n2610 ;
  assign new_n4626 = ~new_n4624 & ~new_n4625 ;
  assign new_n4627 = new_n4623 & new_n4626 ;
  assign new_n4628 = ~new_n2729 & new_n4627 ;
  assign new_n4629 = ~new_n4620 & new_n4628 ;
  assign new_n4630 = ~new_n4616 & new_n4629 ;
  assign new_n4631 = new_n3735 & ~new_n4630 ;
  assign new_n4632 = ~new_n4545 & new_n4631 ;
  assign new_n4633 = ~new_n4550 & ~new_n4632 ;
  assign new_n4634 = ~new_n4549 & new_n4633 ;
  assign new_n4635 = ~lo0298 & ~new_n4634 ;
  assign new_n4636 = ~new_n3001 & new_n3914 ;
  assign new_n4637 = ~lo0297 & ~new_n3464 ;
  assign new_n4638 = ~new_n4636 & ~new_n4637 ;
  assign new_n4639 = lo0298 & ~new_n4638 ;
  assign new_n4640 = ~new_n4635 & ~new_n4639 ;
  assign new_n4641 = new_n3102 & ~new_n4640 ;
  assign new_n4642 = ~new_n3102 & ~new_n3817 ;
  assign new_n4643 = ~new_n4641 & ~new_n4642 ;
  assign new_n4644 = lo0647 & new_n3170 ;
  assign new_n4645 = lo0646 & new_n3173 ;
  assign new_n4646 = ~new_n3172 & ~new_n4645 ;
  assign new_n4647 = ~new_n4644 & new_n4646 ;
  assign new_n4648 = ~lo0059 & ~new_n4647 ;
  assign new_n4649 = lo0059 & new_n4647 ;
  assign new_n4650 = ~new_n4648 & ~new_n4649 ;
  assign new_n4651 = lo0645 & ~new_n4650 ;
  assign new_n4652 = ~lo0645 & new_n4648 ;
  assign new_n4653 = lo0059 & lo0648 ;
  assign new_n4654 = ~new_n4647 & new_n4653 ;
  assign new_n4655 = ~new_n4652 & ~new_n4654 ;
  assign new_n4656 = ~new_n4651 & new_n4655 ;
  assign new_n4657 = lo0655 & new_n3170 ;
  assign new_n4658 = lo0654 & new_n3173 ;
  assign new_n4659 = ~new_n3172 & ~new_n4658 ;
  assign new_n4660 = ~new_n4657 & new_n4659 ;
  assign new_n4661 = ~lo0059 & ~new_n4660 ;
  assign new_n4662 = lo0059 & new_n4660 ;
  assign new_n4663 = ~new_n4661 & ~new_n4662 ;
  assign new_n4664 = lo0653 & ~new_n4663 ;
  assign new_n4665 = ~lo0653 & new_n4661 ;
  assign new_n4666 = lo0059 & lo0656 ;
  assign new_n4667 = ~new_n4660 & new_n4666 ;
  assign new_n4668 = ~new_n4665 & ~new_n4667 ;
  assign new_n4669 = ~new_n4664 & new_n4668 ;
  assign new_n4670 = new_n3186 & ~new_n4669 ;
  assign new_n4671 = lo0651 & new_n3170 ;
  assign new_n4672 = lo0650 & new_n3204 ;
  assign new_n4673 = ~new_n3172 & ~new_n4672 ;
  assign new_n4674 = ~new_n4671 & new_n4673 ;
  assign new_n4675 = ~lo0061 & ~new_n4674 ;
  assign new_n4676 = lo0061 & new_n4674 ;
  assign new_n4677 = ~new_n4675 & ~new_n4676 ;
  assign new_n4678 = lo0649 & ~new_n4677 ;
  assign new_n4679 = ~lo0649 & new_n4675 ;
  assign new_n4680 = lo0061 & lo0652 ;
  assign new_n4681 = ~new_n4674 & new_n4680 ;
  assign new_n4682 = ~new_n4679 & ~new_n4681 ;
  assign new_n4683 = ~new_n4678 & new_n4682 ;
  assign new_n4684 = new_n3202 & ~new_n4683 ;
  assign new_n4685 = ~new_n3201 & ~new_n4684 ;
  assign new_n4686 = ~new_n4670 & new_n4685 ;
  assign new_n4687 = ~lo0063 & ~new_n4686 ;
  assign new_n4688 = lo0063 & new_n4686 ;
  assign new_n4689 = ~new_n4687 & ~new_n4688 ;
  assign new_n4690 = ~new_n4656 & ~new_n4689 ;
  assign new_n4691 = new_n4656 & new_n4687 ;
  assign new_n4692 = lo0659 & new_n3170 ;
  assign new_n4693 = lo0658 & new_n3204 ;
  assign new_n4694 = ~new_n3172 & ~new_n4693 ;
  assign new_n4695 = ~new_n4692 & new_n4694 ;
  assign new_n4696 = ~lo0061 & ~new_n4695 ;
  assign new_n4697 = lo0061 & new_n4695 ;
  assign new_n4698 = ~new_n4696 & ~new_n4697 ;
  assign new_n4699 = lo0657 & ~new_n4698 ;
  assign new_n4700 = ~lo0657 & new_n4696 ;
  assign new_n4701 = lo0061 & lo0660 ;
  assign new_n4702 = ~new_n4695 & new_n4701 ;
  assign new_n4703 = ~new_n4700 & ~new_n4702 ;
  assign new_n4704 = ~new_n4699 & new_n4703 ;
  assign new_n4705 = lo0063 & ~new_n4704 ;
  assign new_n4706 = ~new_n4686 & new_n4705 ;
  assign new_n4707 = ~new_n4691 & ~new_n4706 ;
  assign new_n4708 = ~new_n4690 & new_n4707 ;
  assign new_n4709 = new_n3169 & ~new_n4708 ;
  assign new_n4710 = ~new_n3160 & new_n3806 ;
  assign new_n4711 = lo1400 & new_n3246 ;
  assign new_n4712 = lo1349 & new_n3254 ;
  assign new_n4713 = lo0662 & new_n3258 ;
  assign new_n4714 = ~new_n4712 & ~new_n4713 ;
  assign new_n4715 = ~new_n4711 & new_n4714 ;
  assign new_n4716 = lo1399 & new_n3267 ;
  assign new_n4717 = lo1401 & new_n3270 ;
  assign new_n4718 = lo0661 & new_n3274 ;
  assign new_n4719 = ~new_n4717 & ~new_n4718 ;
  assign new_n4720 = ~new_n4716 & new_n4719 ;
  assign new_n4721 = ~new_n3265 & new_n4720 ;
  assign new_n4722 = new_n4715 & new_n4721 ;
  assign new_n4723 = ~new_n4710 & new_n4722 ;
  assign new_n4724 = ~new_n4709 & new_n4723 ;
  assign new_n4725 = new_n3141 & ~new_n4724 ;
  assign new_n4726 = new_n3140 & ~new_n4725 ;
  assign new_n4727 = ~new_n3121 & ~new_n4726 ;
  assign new_n4728 = new_n3121 & new_n4726 ;
  assign new_n4729 = ~new_n4727 & ~new_n4728 ;
  assign new_n4730 = lo0655 & ~new_n4729 ;
  assign new_n4731 = ~lo0655 & new_n4727 ;
  assign new_n4732 = new_n3121 & new_n3806 ;
  assign new_n4733 = ~new_n4726 & new_n4732 ;
  assign new_n4734 = ~new_n4731 & ~new_n4733 ;
  assign new_n4735 = ~new_n4730 & new_n4734 ;
  assign new_n4736 = ~new_n3112 & new_n4735 ;
  assign new_n4737 = new_n3112 & ~new_n4735 ;
  assign new_n4738 = ~new_n4736 & ~new_n4737 ;
  assign new_n4739 = lo0725 & new_n2506 ;
  assign new_n4740 = lo0724 & new_n2831 ;
  assign new_n4741 = ~new_n2521 & ~new_n4740 ;
  assign new_n4742 = ~new_n4739 & new_n4741 ;
  assign new_n4743 = ~lo0252 & ~new_n4742 ;
  assign new_n4744 = lo0252 & new_n4742 ;
  assign new_n4745 = ~new_n4743 & ~new_n4744 ;
  assign new_n4746 = lo0723 & ~new_n4745 ;
  assign new_n4747 = ~lo0723 & new_n4743 ;
  assign new_n4748 = lo0252 & lo0726 ;
  assign new_n4749 = ~new_n4742 & new_n4748 ;
  assign new_n4750 = ~new_n4747 & ~new_n4749 ;
  assign new_n4751 = ~new_n4746 & new_n4750 ;
  assign new_n4752 = lo0733 & new_n2506 ;
  assign new_n4753 = lo0732 & new_n2522 ;
  assign new_n4754 = ~new_n2521 & ~new_n4753 ;
  assign new_n4755 = ~new_n4752 & new_n4754 ;
  assign new_n4756 = ~lo0251 & ~new_n4755 ;
  assign new_n4757 = lo0251 & new_n4755 ;
  assign new_n4758 = ~new_n4756 & ~new_n4757 ;
  assign new_n4759 = lo0731 & ~new_n4758 ;
  assign new_n4760 = ~lo0731 & new_n4756 ;
  assign new_n4761 = lo0251 & lo0734 ;
  assign new_n4762 = ~new_n4755 & new_n4761 ;
  assign new_n4763 = ~new_n4760 & ~new_n4762 ;
  assign new_n4764 = ~new_n4759 & new_n4763 ;
  assign new_n4765 = new_n2490 & ~new_n4764 ;
  assign new_n4766 = lo0729 & new_n2506 ;
  assign new_n4767 = lo0728 & new_n2522 ;
  assign new_n4768 = ~new_n2521 & ~new_n4767 ;
  assign new_n4769 = ~new_n4766 & new_n4768 ;
  assign new_n4770 = ~lo0251 & ~new_n4769 ;
  assign new_n4771 = lo0251 & new_n4769 ;
  assign new_n4772 = ~new_n4770 & ~new_n4771 ;
  assign new_n4773 = lo0727 & ~new_n4772 ;
  assign new_n4774 = ~lo0727 & new_n4770 ;
  assign new_n4775 = lo0251 & lo0730 ;
  assign new_n4776 = ~new_n4769 & new_n4775 ;
  assign new_n4777 = ~new_n4774 & ~new_n4776 ;
  assign new_n4778 = ~new_n4773 & new_n4777 ;
  assign new_n4779 = new_n3310 & ~new_n4778 ;
  assign new_n4780 = ~new_n2492 & ~new_n4779 ;
  assign new_n4781 = ~new_n4765 & new_n4780 ;
  assign new_n4782 = ~lo0250 & ~new_n4781 ;
  assign new_n4783 = lo0250 & new_n4781 ;
  assign new_n4784 = ~new_n4782 & ~new_n4783 ;
  assign new_n4785 = ~new_n4751 & ~new_n4784 ;
  assign new_n4786 = new_n4751 & new_n4782 ;
  assign new_n4787 = lo0737 & new_n2506 ;
  assign new_n4788 = lo0736 & new_n2831 ;
  assign new_n4789 = ~new_n2521 & ~new_n4788 ;
  assign new_n4790 = ~new_n4787 & new_n4789 ;
  assign new_n4791 = ~lo0252 & ~new_n4790 ;
  assign new_n4792 = lo0252 & new_n4790 ;
  assign new_n4793 = ~new_n4791 & ~new_n4792 ;
  assign new_n4794 = lo0735 & ~new_n4793 ;
  assign new_n4795 = ~lo0735 & new_n4791 ;
  assign new_n4796 = lo0252 & lo0738 ;
  assign new_n4797 = ~new_n4790 & new_n4796 ;
  assign new_n4798 = ~new_n4795 & ~new_n4797 ;
  assign new_n4799 = ~new_n4794 & new_n4798 ;
  assign new_n4800 = lo0250 & ~new_n4799 ;
  assign new_n4801 = ~new_n4781 & new_n4800 ;
  assign new_n4802 = ~new_n4786 & ~new_n4801 ;
  assign new_n4803 = ~new_n4785 & new_n4802 ;
  assign new_n4804 = new_n2489 & ~new_n4803 ;
  assign new_n4805 = lo0091 & lo0100 ;
  assign new_n4806 = ~new_n2715 & ~new_n4805 ;
  assign new_n4807 = lo0090 & ~new_n4806 ;
  assign new_n4808 = ~new_n2483 & new_n4807 ;
  assign new_n4809 = lo0739 & new_n2601 ;
  assign new_n4810 = lo0741 & new_n2605 ;
  assign new_n4811 = ~new_n4809 & ~new_n4810 ;
  assign new_n4812 = lo0740 & new_n2613 ;
  assign new_n4813 = lo1359 & new_n2610 ;
  assign new_n4814 = ~new_n4812 & ~new_n4813 ;
  assign new_n4815 = new_n4811 & new_n4814 ;
  assign new_n4816 = ~new_n2729 & new_n4815 ;
  assign new_n4817 = ~new_n4808 & new_n4816 ;
  assign new_n4818 = ~new_n4804 & new_n4817 ;
  assign new_n4819 = new_n3737 & ~new_n4818 ;
  assign new_n4820 = lo0685 & new_n2490 ;
  assign new_n4821 = lo0684 & new_n2493 ;
  assign new_n4822 = ~new_n2492 & ~new_n4821 ;
  assign new_n4823 = ~new_n4820 & new_n4822 ;
  assign new_n4824 = ~lo0249 & ~new_n4823 ;
  assign new_n4825 = lo0249 & new_n4823 ;
  assign new_n4826 = ~new_n4824 & ~new_n4825 ;
  assign new_n4827 = lo0683 & ~new_n4826 ;
  assign new_n4828 = ~lo0683 & new_n4824 ;
  assign new_n4829 = lo0249 & lo0686 ;
  assign new_n4830 = ~new_n4823 & new_n4829 ;
  assign new_n4831 = ~new_n4828 & ~new_n4830 ;
  assign new_n4832 = ~new_n4827 & new_n4831 ;
  assign new_n4833 = lo1351 & new_n2490 ;
  assign new_n4834 = lo0692 & new_n3310 ;
  assign new_n4835 = ~new_n2492 & ~new_n4834 ;
  assign new_n4836 = ~new_n4833 & new_n4835 ;
  assign new_n4837 = ~lo0250 & ~new_n4836 ;
  assign new_n4838 = lo0250 & new_n4836 ;
  assign new_n4839 = ~new_n4837 & ~new_n4838 ;
  assign new_n4840 = lo0691 & ~new_n4839 ;
  assign new_n4841 = ~lo0691 & new_n4837 ;
  assign new_n4842 = lo0250 & lo0693 ;
  assign new_n4843 = ~new_n4836 & new_n4842 ;
  assign new_n4844 = ~new_n4841 & ~new_n4843 ;
  assign new_n4845 = ~new_n4840 & new_n4844 ;
  assign new_n4846 = new_n2506 & ~new_n4845 ;
  assign new_n4847 = lo0689 & new_n2490 ;
  assign new_n4848 = lo0688 & new_n3310 ;
  assign new_n4849 = ~new_n2492 & ~new_n4848 ;
  assign new_n4850 = ~new_n4847 & new_n4849 ;
  assign new_n4851 = ~lo0250 & ~new_n4850 ;
  assign new_n4852 = lo0250 & new_n4850 ;
  assign new_n4853 = ~new_n4851 & ~new_n4852 ;
  assign new_n4854 = lo0687 & ~new_n4853 ;
  assign new_n4855 = ~lo0687 & new_n4851 ;
  assign new_n4856 = lo0250 & lo0690 ;
  assign new_n4857 = ~new_n4850 & new_n4856 ;
  assign new_n4858 = ~new_n4855 & ~new_n4857 ;
  assign new_n4859 = ~new_n4854 & new_n4858 ;
  assign new_n4860 = new_n2831 & ~new_n4859 ;
  assign new_n4861 = ~new_n2521 & ~new_n4860 ;
  assign new_n4862 = ~new_n4846 & new_n4861 ;
  assign new_n4863 = ~lo0252 & ~new_n4862 ;
  assign new_n4864 = lo0252 & new_n4862 ;
  assign new_n4865 = ~new_n4863 & ~new_n4864 ;
  assign new_n4866 = ~new_n4832 & ~new_n4865 ;
  assign new_n4867 = new_n4832 & new_n4863 ;
  assign new_n4868 = lo0696 & new_n2490 ;
  assign new_n4869 = lo0695 & new_n2493 ;
  assign new_n4870 = ~new_n2492 & ~new_n4869 ;
  assign new_n4871 = ~new_n4868 & new_n4870 ;
  assign new_n4872 = ~lo0249 & ~new_n4871 ;
  assign new_n4873 = lo0249 & new_n4871 ;
  assign new_n4874 = ~new_n4872 & ~new_n4873 ;
  assign new_n4875 = lo0694 & ~new_n4874 ;
  assign new_n4876 = ~lo0694 & new_n4872 ;
  assign new_n4877 = lo0249 & lo0697 ;
  assign new_n4878 = ~new_n4871 & new_n4877 ;
  assign new_n4879 = ~new_n4876 & ~new_n4878 ;
  assign new_n4880 = ~new_n4875 & new_n4879 ;
  assign new_n4881 = lo0252 & ~new_n4880 ;
  assign new_n4882 = ~new_n4862 & new_n4881 ;
  assign new_n4883 = ~new_n4867 & ~new_n4882 ;
  assign new_n4884 = ~new_n4866 & new_n4883 ;
  assign new_n4885 = new_n2489 & ~new_n4884 ;
  assign new_n4886 = lo0639 & new_n3367 ;
  assign new_n4887 = lo0638 & new_n3369 ;
  assign new_n4888 = ~new_n4886 & ~new_n4887 ;
  assign new_n4889 = ~new_n3366 & new_n4888 ;
  assign new_n4890 = ~new_n2483 & ~new_n4889 ;
  assign new_n4891 = lo0698 & new_n2720 ;
  assign new_n4892 = ~new_n2721 & ~new_n4891 ;
  assign new_n4893 = new_n2727 & ~new_n4892 ;
  assign new_n4894 = new_n2591 & new_n4893 ;
  assign new_n4895 = lo0699 & new_n2601 ;
  assign new_n4896 = lo0701 & new_n2605 ;
  assign new_n4897 = ~new_n4895 & ~new_n4896 ;
  assign new_n4898 = lo0700 & new_n2610 ;
  assign new_n4899 = lo0702 & new_n2613 ;
  assign new_n4900 = ~new_n4898 & ~new_n4899 ;
  assign new_n4901 = new_n4897 & new_n4900 ;
  assign new_n4902 = ~new_n4894 & new_n4901 ;
  assign new_n4903 = ~new_n4890 & new_n4902 ;
  assign new_n4904 = ~new_n4885 & new_n4903 ;
  assign new_n4905 = new_n4180 & ~new_n4904 ;
  assign new_n4906 = ~new_n3819 & ~new_n4905 ;
  assign new_n4907 = ~new_n4819 & new_n4906 ;
  assign new_n4908 = new_n3736 & ~new_n4907 ;
  assign new_n4909 = ~new_n3736 & new_n4907 ;
  assign new_n4910 = ~new_n4908 & ~new_n4909 ;
  assign new_n4911 = ~new_n4541 & ~new_n4910 ;
  assign new_n4912 = new_n4541 & new_n4908 ;
  assign new_n4913 = lo0324 & new_n2506 ;
  assign new_n4914 = lo0323 & new_n2831 ;
  assign new_n4915 = ~new_n2521 & ~new_n4914 ;
  assign new_n4916 = ~new_n4913 & new_n4915 ;
  assign new_n4917 = ~lo0252 & ~new_n4916 ;
  assign new_n4918 = lo0252 & new_n4916 ;
  assign new_n4919 = ~new_n4917 & ~new_n4918 ;
  assign new_n4920 = lo0322 & ~new_n4919 ;
  assign new_n4921 = ~lo0322 & new_n4917 ;
  assign new_n4922 = lo0252 & lo0325 ;
  assign new_n4923 = ~new_n4916 & new_n4922 ;
  assign new_n4924 = ~new_n4921 & ~new_n4923 ;
  assign new_n4925 = ~new_n4920 & new_n4924 ;
  assign new_n4926 = lo0332 & new_n2506 ;
  assign new_n4927 = lo0331 & new_n2831 ;
  assign new_n4928 = ~new_n2521 & ~new_n4927 ;
  assign new_n4929 = ~new_n4926 & new_n4928 ;
  assign new_n4930 = ~lo0252 & ~new_n4929 ;
  assign new_n4931 = lo0252 & new_n4929 ;
  assign new_n4932 = ~new_n4930 & ~new_n4931 ;
  assign new_n4933 = lo0330 & ~new_n4932 ;
  assign new_n4934 = ~lo0330 & new_n4930 ;
  assign new_n4935 = lo0252 & lo0333 ;
  assign new_n4936 = ~new_n4929 & new_n4935 ;
  assign new_n4937 = ~new_n4934 & ~new_n4936 ;
  assign new_n4938 = ~new_n4933 & new_n4937 ;
  assign new_n4939 = new_n2490 & ~new_n4938 ;
  assign new_n4940 = lo0328 & new_n2506 ;
  assign new_n4941 = lo0327 & new_n2522 ;
  assign new_n4942 = ~new_n2521 & ~new_n4941 ;
  assign new_n4943 = ~new_n4940 & new_n4942 ;
  assign new_n4944 = ~lo0251 & ~new_n4943 ;
  assign new_n4945 = lo0251 & new_n4943 ;
  assign new_n4946 = ~new_n4944 & ~new_n4945 ;
  assign new_n4947 = lo0326 & ~new_n4946 ;
  assign new_n4948 = ~lo0326 & new_n4944 ;
  assign new_n4949 = lo0251 & lo0329 ;
  assign new_n4950 = ~new_n4943 & new_n4949 ;
  assign new_n4951 = ~new_n4948 & ~new_n4950 ;
  assign new_n4952 = ~new_n4947 & new_n4951 ;
  assign new_n4953 = new_n2493 & ~new_n4952 ;
  assign new_n4954 = ~new_n2492 & ~new_n4953 ;
  assign new_n4955 = ~new_n4939 & new_n4954 ;
  assign new_n4956 = ~lo0249 & ~new_n4955 ;
  assign new_n4957 = lo0249 & new_n4955 ;
  assign new_n4958 = ~new_n4956 & ~new_n4957 ;
  assign new_n4959 = ~new_n4925 & ~new_n4958 ;
  assign new_n4960 = new_n4925 & new_n4956 ;
  assign new_n4961 = lo0336 & new_n2506 ;
  assign new_n4962 = lo0335 & new_n2522 ;
  assign new_n4963 = ~new_n2521 & ~new_n4962 ;
  assign new_n4964 = ~new_n4961 & new_n4963 ;
  assign new_n4965 = ~lo0251 & ~new_n4964 ;
  assign new_n4966 = lo0251 & new_n4964 ;
  assign new_n4967 = ~new_n4965 & ~new_n4966 ;
  assign new_n4968 = lo0334 & ~new_n4967 ;
  assign new_n4969 = ~lo0334 & new_n4965 ;
  assign new_n4970 = lo0251 & lo0337 ;
  assign new_n4971 = ~new_n4964 & new_n4970 ;
  assign new_n4972 = ~new_n4969 & ~new_n4971 ;
  assign new_n4973 = ~new_n4968 & new_n4972 ;
  assign new_n4974 = lo0249 & ~new_n4973 ;
  assign new_n4975 = ~new_n4955 & new_n4974 ;
  assign new_n4976 = ~new_n4960 & ~new_n4975 ;
  assign new_n4977 = ~new_n4959 & new_n4976 ;
  assign new_n4978 = new_n2489 & ~new_n4977 ;
  assign new_n4979 = lo0091 & lo0338 ;
  assign new_n4980 = ~new_n2715 & ~new_n4979 ;
  assign new_n4981 = lo0090 & ~new_n4980 ;
  assign new_n4982 = ~new_n2483 & new_n4981 ;
  assign new_n4983 = lo0339 & new_n2601 ;
  assign new_n4984 = lo0341 & new_n2605 ;
  assign new_n4985 = ~new_n4983 & ~new_n4984 ;
  assign new_n4986 = lo0340 & new_n2613 ;
  assign new_n4987 = lo1306 & new_n2610 ;
  assign new_n4988 = ~new_n4986 & ~new_n4987 ;
  assign new_n4989 = new_n4985 & new_n4988 ;
  assign new_n4990 = ~new_n2729 & new_n4989 ;
  assign new_n4991 = ~new_n4982 & new_n4990 ;
  assign new_n4992 = ~new_n4978 & new_n4991 ;
  assign new_n4993 = ~new_n3736 & ~new_n4992 ;
  assign new_n4994 = ~new_n4907 & new_n4993 ;
  assign new_n4995 = ~new_n4912 & ~new_n4994 ;
  assign new_n4996 = ~new_n4911 & new_n4995 ;
  assign new_n4997 = ~lo0298 & ~new_n4996 ;
  assign new_n4998 = ~new_n3464 & new_n3914 ;
  assign new_n4999 = ~lo0297 & ~new_n3817 ;
  assign new_n5000 = ~new_n4998 & ~new_n4999 ;
  assign new_n5001 = lo0298 & ~new_n5000 ;
  assign new_n5002 = ~new_n4997 & ~new_n5001 ;
  assign new_n5003 = new_n3102 & ~new_n5002 ;
  assign new_n5004 = ~new_n3102 & ~new_n4097 ;
  assign new_n5005 = ~new_n5003 & ~new_n5004 ;
  assign new_n5006 = lo0666 & new_n3186 ;
  assign new_n5007 = lo0665 & new_n3559 ;
  assign new_n5008 = ~new_n3201 & ~new_n5007 ;
  assign new_n5009 = ~new_n5006 & new_n5008 ;
  assign new_n5010 = ~lo0065 & ~new_n5009 ;
  assign new_n5011 = lo0065 & new_n5009 ;
  assign new_n5012 = ~new_n5010 & ~new_n5011 ;
  assign new_n5013 = lo0664 & ~new_n5012 ;
  assign new_n5014 = ~lo0664 & new_n5010 ;
  assign new_n5015 = lo0065 & lo0667 ;
  assign new_n5016 = ~new_n5009 & new_n5015 ;
  assign new_n5017 = ~new_n5014 & ~new_n5016 ;
  assign new_n5018 = ~new_n5013 & new_n5017 ;
  assign new_n5019 = lo0674 & new_n3186 ;
  assign new_n5020 = lo0673 & new_n3559 ;
  assign new_n5021 = ~new_n3201 & ~new_n5020 ;
  assign new_n5022 = ~new_n5019 & new_n5021 ;
  assign new_n5023 = ~lo0065 & ~new_n5022 ;
  assign new_n5024 = lo0065 & new_n5022 ;
  assign new_n5025 = ~new_n5023 & ~new_n5024 ;
  assign new_n5026 = lo0672 & ~new_n5025 ;
  assign new_n5027 = ~lo0672 & new_n5023 ;
  assign new_n5028 = lo0065 & lo0675 ;
  assign new_n5029 = ~new_n5022 & new_n5028 ;
  assign new_n5030 = ~new_n5027 & ~new_n5029 ;
  assign new_n5031 = ~new_n5026 & new_n5030 ;
  assign new_n5032 = new_n3170 & ~new_n5031 ;
  assign new_n5033 = lo0670 & new_n3186 ;
  assign new_n5034 = lo0669 & new_n3202 ;
  assign new_n5035 = ~new_n3201 & ~new_n5034 ;
  assign new_n5036 = ~new_n5033 & new_n5035 ;
  assign new_n5037 = ~lo0063 & ~new_n5036 ;
  assign new_n5038 = lo0063 & new_n5036 ;
  assign new_n5039 = ~new_n5037 & ~new_n5038 ;
  assign new_n5040 = lo0668 & ~new_n5039 ;
  assign new_n5041 = ~lo0668 & new_n5037 ;
  assign new_n5042 = lo0063 & lo0671 ;
  assign new_n5043 = ~new_n5036 & new_n5042 ;
  assign new_n5044 = ~new_n5041 & ~new_n5043 ;
  assign new_n5045 = ~new_n5040 & new_n5044 ;
  assign new_n5046 = new_n3173 & ~new_n5045 ;
  assign new_n5047 = ~new_n3172 & ~new_n5046 ;
  assign new_n5048 = ~new_n5032 & new_n5047 ;
  assign new_n5049 = ~lo0059 & ~new_n5048 ;
  assign new_n5050 = lo0059 & new_n5048 ;
  assign new_n5051 = ~new_n5049 & ~new_n5050 ;
  assign new_n5052 = ~new_n5018 & ~new_n5051 ;
  assign new_n5053 = new_n5018 & new_n5049 ;
  assign new_n5054 = lo0678 & new_n3186 ;
  assign new_n5055 = lo0677 & new_n3202 ;
  assign new_n5056 = ~new_n3201 & ~new_n5055 ;
  assign new_n5057 = ~new_n5054 & new_n5056 ;
  assign new_n5058 = ~lo0063 & ~new_n5057 ;
  assign new_n5059 = lo0063 & new_n5057 ;
  assign new_n5060 = ~new_n5058 & ~new_n5059 ;
  assign new_n5061 = lo0676 & ~new_n5060 ;
  assign new_n5062 = ~lo0676 & new_n5058 ;
  assign new_n5063 = lo0063 & lo0679 ;
  assign new_n5064 = ~new_n5057 & new_n5063 ;
  assign new_n5065 = ~new_n5062 & ~new_n5064 ;
  assign new_n5066 = ~new_n5061 & new_n5065 ;
  assign new_n5067 = lo0059 & ~new_n5066 ;
  assign new_n5068 = ~new_n5048 & new_n5067 ;
  assign new_n5069 = ~new_n5053 & ~new_n5068 ;
  assign new_n5070 = ~new_n5052 & new_n5069 ;
  assign new_n5071 = new_n3169 & ~new_n5070 ;
  assign new_n5072 = ~new_n3160 & new_n4086 ;
  assign new_n5073 = lo1415 & new_n3246 ;
  assign new_n5074 = lo1350 & new_n3254 ;
  assign new_n5075 = lo0681 & new_n3258 ;
  assign new_n5076 = ~new_n5074 & ~new_n5075 ;
  assign new_n5077 = ~new_n5073 & new_n5076 ;
  assign new_n5078 = lo1414 & new_n3267 ;
  assign new_n5079 = lo1416 & new_n3270 ;
  assign new_n5080 = lo0680 & new_n3274 ;
  assign new_n5081 = ~new_n5079 & ~new_n5080 ;
  assign new_n5082 = ~new_n5078 & new_n5081 ;
  assign new_n5083 = ~new_n3265 & new_n5082 ;
  assign new_n5084 = new_n5077 & new_n5083 ;
  assign new_n5085 = ~new_n5072 & new_n5084 ;
  assign new_n5086 = ~new_n5071 & new_n5085 ;
  assign new_n5087 = new_n3141 & ~new_n5086 ;
  assign new_n5088 = new_n3140 & ~new_n5087 ;
  assign new_n5089 = ~new_n3121 & ~new_n5088 ;
  assign new_n5090 = new_n3121 & new_n5088 ;
  assign new_n5091 = ~new_n5089 & ~new_n5090 ;
  assign new_n5092 = lo0674 & ~new_n5091 ;
  assign new_n5093 = ~lo0674 & new_n5089 ;
  assign new_n5094 = new_n3121 & new_n4086 ;
  assign new_n5095 = ~new_n5088 & new_n5094 ;
  assign new_n5096 = ~new_n5093 & ~new_n5095 ;
  assign new_n5097 = ~new_n5092 & new_n5096 ;
  assign new_n5098 = ~new_n3112 & new_n5097 ;
  assign new_n5099 = new_n3112 & ~new_n5097 ;
  assign new_n5100 = ~new_n5098 & ~new_n5099 ;
  assign new_n5101 = lo0808 & new_n2506 ;
  assign new_n5102 = lo0807 & new_n2831 ;
  assign new_n5103 = ~new_n2521 & ~new_n5102 ;
  assign new_n5104 = ~new_n5101 & new_n5103 ;
  assign new_n5105 = ~lo0252 & ~new_n5104 ;
  assign new_n5106 = lo0252 & new_n5104 ;
  assign new_n5107 = ~new_n5105 & ~new_n5106 ;
  assign new_n5108 = lo0806 & ~new_n5107 ;
  assign new_n5109 = ~lo0806 & new_n5105 ;
  assign new_n5110 = lo0252 & lo0809 ;
  assign new_n5111 = ~new_n5104 & new_n5110 ;
  assign new_n5112 = ~new_n5109 & ~new_n5111 ;
  assign new_n5113 = ~new_n5108 & new_n5112 ;
  assign new_n5114 = lo0816 & new_n2506 ;
  assign new_n5115 = lo0815 & new_n2522 ;
  assign new_n5116 = ~new_n2521 & ~new_n5115 ;
  assign new_n5117 = ~new_n5114 & new_n5116 ;
  assign new_n5118 = ~lo0251 & ~new_n5117 ;
  assign new_n5119 = lo0251 & new_n5117 ;
  assign new_n5120 = ~new_n5118 & ~new_n5119 ;
  assign new_n5121 = lo0814 & ~new_n5120 ;
  assign new_n5122 = ~lo0814 & new_n5118 ;
  assign new_n5123 = lo0251 & lo0817 ;
  assign new_n5124 = ~new_n5117 & new_n5123 ;
  assign new_n5125 = ~new_n5122 & ~new_n5124 ;
  assign new_n5126 = ~new_n5121 & new_n5125 ;
  assign new_n5127 = new_n2490 & ~new_n5126 ;
  assign new_n5128 = lo0812 & new_n2506 ;
  assign new_n5129 = lo0811 & new_n2522 ;
  assign new_n5130 = ~new_n2521 & ~new_n5129 ;
  assign new_n5131 = ~new_n5128 & new_n5130 ;
  assign new_n5132 = ~lo0251 & ~new_n5131 ;
  assign new_n5133 = lo0251 & new_n5131 ;
  assign new_n5134 = ~new_n5132 & ~new_n5133 ;
  assign new_n5135 = lo0810 & ~new_n5134 ;
  assign new_n5136 = ~lo0810 & new_n5132 ;
  assign new_n5137 = lo0251 & lo0813 ;
  assign new_n5138 = ~new_n5131 & new_n5137 ;
  assign new_n5139 = ~new_n5136 & ~new_n5138 ;
  assign new_n5140 = ~new_n5135 & new_n5139 ;
  assign new_n5141 = new_n3310 & ~new_n5140 ;
  assign new_n5142 = ~new_n2492 & ~new_n5141 ;
  assign new_n5143 = ~new_n5127 & new_n5142 ;
  assign new_n5144 = ~lo0250 & ~new_n5143 ;
  assign new_n5145 = lo0250 & new_n5143 ;
  assign new_n5146 = ~new_n5144 & ~new_n5145 ;
  assign new_n5147 = ~new_n5113 & ~new_n5146 ;
  assign new_n5148 = new_n5113 & new_n5144 ;
  assign new_n5149 = lo0820 & new_n2506 ;
  assign new_n5150 = lo0819 & new_n2831 ;
  assign new_n5151 = ~new_n2521 & ~new_n5150 ;
  assign new_n5152 = ~new_n5149 & new_n5151 ;
  assign new_n5153 = ~lo0252 & ~new_n5152 ;
  assign new_n5154 = lo0252 & new_n5152 ;
  assign new_n5155 = ~new_n5153 & ~new_n5154 ;
  assign new_n5156 = lo0818 & ~new_n5155 ;
  assign new_n5157 = ~lo0818 & new_n5153 ;
  assign new_n5158 = lo0252 & lo0821 ;
  assign new_n5159 = ~new_n5152 & new_n5158 ;
  assign new_n5160 = ~new_n5157 & ~new_n5159 ;
  assign new_n5161 = ~new_n5156 & new_n5160 ;
  assign new_n5162 = lo0250 & ~new_n5161 ;
  assign new_n5163 = ~new_n5143 & new_n5162 ;
  assign new_n5164 = ~new_n5148 & ~new_n5163 ;
  assign new_n5165 = ~new_n5147 & new_n5164 ;
  assign new_n5166 = new_n2489 & ~new_n5165 ;
  assign new_n5167 = lo0801 & new_n3367 ;
  assign new_n5168 = lo0800 & new_n3369 ;
  assign new_n5169 = ~new_n5167 & ~new_n5168 ;
  assign new_n5170 = ~new_n3366 & new_n5169 ;
  assign new_n5171 = ~new_n2483 & ~new_n5170 ;
  assign new_n5172 = ~lo0102 & new_n2720 ;
  assign new_n5173 = lo0822 & new_n5172 ;
  assign new_n5174 = lo0104 & ~new_n5172 ;
  assign new_n5175 = ~new_n5173 & ~new_n5174 ;
  assign new_n5176 = new_n2726 & ~new_n5175 ;
  assign new_n5177 = new_n2591 & new_n5176 ;
  assign new_n5178 = lo0824 & new_n2613 ;
  assign new_n5179 = lo0823 & new_n2605 ;
  assign new_n5180 = ~new_n5178 & ~new_n5179 ;
  assign new_n5181 = lo0825 & new_n2601 ;
  assign new_n5182 = lo1381 & new_n2610 ;
  assign new_n5183 = ~new_n5181 & ~new_n5182 ;
  assign new_n5184 = new_n5180 & new_n5183 ;
  assign new_n5185 = ~new_n5177 & new_n5184 ;
  assign new_n5186 = ~new_n5171 & new_n5185 ;
  assign new_n5187 = ~new_n5166 & new_n5186 ;
  assign new_n5188 = ~new_n2824 & new_n3737 ;
  assign new_n5189 = new_n3820 & ~new_n4818 ;
  assign new_n5190 = ~new_n3819 & ~new_n5189 ;
  assign new_n5191 = ~new_n5188 & new_n5190 ;
  assign new_n5192 = ~new_n3735 & ~new_n5191 ;
  assign new_n5193 = new_n3735 & new_n5191 ;
  assign new_n5194 = ~new_n5192 & ~new_n5193 ;
  assign new_n5195 = ~new_n5187 & ~new_n5194 ;
  assign new_n5196 = new_n5187 & new_n5192 ;
  assign new_n5197 = lo0766 & new_n2490 ;
  assign new_n5198 = lo0765 & new_n2493 ;
  assign new_n5199 = ~new_n2492 & ~new_n5198 ;
  assign new_n5200 = ~new_n5197 & new_n5199 ;
  assign new_n5201 = ~lo0249 & ~new_n5200 ;
  assign new_n5202 = lo0249 & new_n5200 ;
  assign new_n5203 = ~new_n5201 & ~new_n5202 ;
  assign new_n5204 = lo0764 & ~new_n5203 ;
  assign new_n5205 = ~lo0764 & new_n5201 ;
  assign new_n5206 = lo0249 & lo0767 ;
  assign new_n5207 = ~new_n5200 & new_n5206 ;
  assign new_n5208 = ~new_n5205 & ~new_n5207 ;
  assign new_n5209 = ~new_n5204 & new_n5208 ;
  assign new_n5210 = lo0774 & new_n2490 ;
  assign new_n5211 = lo0773 & new_n3310 ;
  assign new_n5212 = ~new_n2492 & ~new_n5211 ;
  assign new_n5213 = ~new_n5210 & new_n5212 ;
  assign new_n5214 = ~lo0250 & ~new_n5213 ;
  assign new_n5215 = lo0250 & new_n5213 ;
  assign new_n5216 = ~new_n5214 & ~new_n5215 ;
  assign new_n5217 = lo0772 & ~new_n5216 ;
  assign new_n5218 = ~lo0772 & new_n5214 ;
  assign new_n5219 = lo0250 & lo0775 ;
  assign new_n5220 = ~new_n5213 & new_n5219 ;
  assign new_n5221 = ~new_n5218 & ~new_n5220 ;
  assign new_n5222 = ~new_n5217 & new_n5221 ;
  assign new_n5223 = new_n2506 & ~new_n5222 ;
  assign new_n5224 = lo0770 & new_n2490 ;
  assign new_n5225 = lo0769 & new_n3310 ;
  assign new_n5226 = ~new_n2492 & ~new_n5225 ;
  assign new_n5227 = ~new_n5224 & new_n5226 ;
  assign new_n5228 = ~lo0250 & ~new_n5227 ;
  assign new_n5229 = lo0250 & new_n5227 ;
  assign new_n5230 = ~new_n5228 & ~new_n5229 ;
  assign new_n5231 = lo0768 & ~new_n5230 ;
  assign new_n5232 = ~lo0768 & new_n5228 ;
  assign new_n5233 = lo0250 & lo0771 ;
  assign new_n5234 = ~new_n5227 & new_n5233 ;
  assign new_n5235 = ~new_n5232 & ~new_n5234 ;
  assign new_n5236 = ~new_n5231 & new_n5235 ;
  assign new_n5237 = new_n2831 & ~new_n5236 ;
  assign new_n5238 = ~new_n2521 & ~new_n5237 ;
  assign new_n5239 = ~new_n5223 & new_n5238 ;
  assign new_n5240 = ~lo0252 & ~new_n5239 ;
  assign new_n5241 = lo0252 & new_n5239 ;
  assign new_n5242 = ~new_n5240 & ~new_n5241 ;
  assign new_n5243 = ~new_n5209 & ~new_n5242 ;
  assign new_n5244 = new_n5209 & new_n5240 ;
  assign new_n5245 = lo0778 & new_n2490 ;
  assign new_n5246 = lo0777 & new_n2493 ;
  assign new_n5247 = ~new_n2492 & ~new_n5246 ;
  assign new_n5248 = ~new_n5245 & new_n5247 ;
  assign new_n5249 = ~lo0249 & ~new_n5248 ;
  assign new_n5250 = lo0249 & new_n5248 ;
  assign new_n5251 = ~new_n5249 & ~new_n5250 ;
  assign new_n5252 = lo0776 & ~new_n5251 ;
  assign new_n5253 = ~lo0776 & new_n5249 ;
  assign new_n5254 = lo0249 & lo0779 ;
  assign new_n5255 = ~new_n5248 & new_n5254 ;
  assign new_n5256 = ~new_n5253 & ~new_n5255 ;
  assign new_n5257 = ~new_n5252 & new_n5256 ;
  assign new_n5258 = lo0252 & ~new_n5257 ;
  assign new_n5259 = ~new_n5239 & new_n5258 ;
  assign new_n5260 = ~new_n5244 & ~new_n5259 ;
  assign new_n5261 = ~new_n5243 & new_n5260 ;
  assign new_n5262 = new_n2489 & ~new_n5261 ;
  assign new_n5263 = lo0091 & lo0780 ;
  assign new_n5264 = ~new_n2715 & ~new_n5263 ;
  assign new_n5265 = lo0090 & ~new_n5264 ;
  assign new_n5266 = ~new_n2483 & new_n5265 ;
  assign new_n5267 = lo0781 & new_n2601 ;
  assign new_n5268 = lo0783 & new_n2605 ;
  assign new_n5269 = ~new_n5267 & ~new_n5268 ;
  assign new_n5270 = lo0782 & new_n2613 ;
  assign new_n5271 = lo1367 & new_n2610 ;
  assign new_n5272 = ~new_n5270 & ~new_n5271 ;
  assign new_n5273 = new_n5269 & new_n5272 ;
  assign new_n5274 = ~new_n2729 & new_n5273 ;
  assign new_n5275 = ~new_n5266 & new_n5274 ;
  assign new_n5276 = ~new_n5262 & new_n5275 ;
  assign new_n5277 = new_n3735 & ~new_n5276 ;
  assign new_n5278 = ~new_n5191 & new_n5277 ;
  assign new_n5279 = ~new_n5196 & ~new_n5278 ;
  assign new_n5280 = ~new_n5195 & new_n5279 ;
  assign new_n5281 = ~lo0298 & ~new_n5280 ;
  assign new_n5282 = ~new_n3817 & new_n3914 ;
  assign new_n5283 = ~lo0297 & ~new_n4097 ;
  assign new_n5284 = ~new_n5282 & ~new_n5283 ;
  assign new_n5285 = lo0298 & ~new_n5284 ;
  assign new_n5286 = ~new_n5281 & ~new_n5285 ;
  assign new_n5287 = new_n3102 & ~new_n5286 ;
  assign new_n5288 = ~new_n3102 & ~new_n4541 ;
  assign new_n5289 = ~new_n5287 & ~new_n5288 ;
  assign new_n5290 = lo0829 & new_n3170 ;
  assign new_n5291 = lo0828 & new_n3173 ;
  assign new_n5292 = ~new_n3172 & ~new_n5291 ;
  assign new_n5293 = ~new_n5290 & new_n5292 ;
  assign new_n5294 = ~lo0059 & ~new_n5293 ;
  assign new_n5295 = lo0059 & new_n5293 ;
  assign new_n5296 = ~new_n5294 & ~new_n5295 ;
  assign new_n5297 = lo0827 & ~new_n5296 ;
  assign new_n5298 = ~lo0827 & new_n5294 ;
  assign new_n5299 = lo0059 & lo0830 ;
  assign new_n5300 = ~new_n5293 & new_n5299 ;
  assign new_n5301 = ~new_n5298 & ~new_n5300 ;
  assign new_n5302 = ~new_n5297 & new_n5301 ;
  assign new_n5303 = lo0837 & new_n3170 ;
  assign new_n5304 = lo0836 & new_n3204 ;
  assign new_n5305 = ~new_n3172 & ~new_n5304 ;
  assign new_n5306 = ~new_n5303 & new_n5305 ;
  assign new_n5307 = ~lo0061 & ~new_n5306 ;
  assign new_n5308 = lo0061 & new_n5306 ;
  assign new_n5309 = ~new_n5307 & ~new_n5308 ;
  assign new_n5310 = lo0835 & ~new_n5309 ;
  assign new_n5311 = ~lo0835 & new_n5307 ;
  assign new_n5312 = lo0061 & lo0838 ;
  assign new_n5313 = ~new_n5306 & new_n5312 ;
  assign new_n5314 = ~new_n5311 & ~new_n5313 ;
  assign new_n5315 = ~new_n5310 & new_n5314 ;
  assign new_n5316 = new_n3186 & ~new_n5315 ;
  assign new_n5317 = lo0833 & new_n3170 ;
  assign new_n5318 = lo0832 & new_n3204 ;
  assign new_n5319 = ~new_n3172 & ~new_n5318 ;
  assign new_n5320 = ~new_n5317 & new_n5319 ;
  assign new_n5321 = ~lo0061 & ~new_n5320 ;
  assign new_n5322 = lo0061 & new_n5320 ;
  assign new_n5323 = ~new_n5321 & ~new_n5322 ;
  assign new_n5324 = lo0831 & ~new_n5323 ;
  assign new_n5325 = ~lo0831 & new_n5321 ;
  assign new_n5326 = lo0061 & lo0834 ;
  assign new_n5327 = ~new_n5320 & new_n5326 ;
  assign new_n5328 = ~new_n5325 & ~new_n5327 ;
  assign new_n5329 = ~new_n5324 & new_n5328 ;
  assign new_n5330 = new_n3559 & ~new_n5329 ;
  assign new_n5331 = ~new_n3201 & ~new_n5330 ;
  assign new_n5332 = ~new_n5316 & new_n5331 ;
  assign new_n5333 = ~lo0065 & ~new_n5332 ;
  assign new_n5334 = lo0065 & new_n5332 ;
  assign new_n5335 = ~new_n5333 & ~new_n5334 ;
  assign new_n5336 = ~new_n5302 & ~new_n5335 ;
  assign new_n5337 = new_n5302 & new_n5333 ;
  assign new_n5338 = lo0841 & new_n3170 ;
  assign new_n5339 = lo0840 & new_n3173 ;
  assign new_n5340 = ~new_n3172 & ~new_n5339 ;
  assign new_n5341 = ~new_n5338 & new_n5340 ;
  assign new_n5342 = ~lo0059 & ~new_n5341 ;
  assign new_n5343 = lo0059 & new_n5341 ;
  assign new_n5344 = ~new_n5342 & ~new_n5343 ;
  assign new_n5345 = lo0839 & ~new_n5344 ;
  assign new_n5346 = ~lo0839 & new_n5342 ;
  assign new_n5347 = lo0059 & lo0842 ;
  assign new_n5348 = ~new_n5341 & new_n5347 ;
  assign new_n5349 = ~new_n5346 & ~new_n5348 ;
  assign new_n5350 = ~new_n5345 & new_n5349 ;
  assign new_n5351 = lo0065 & ~new_n5350 ;
  assign new_n5352 = ~new_n5332 & new_n5351 ;
  assign new_n5353 = ~new_n5337 & ~new_n5352 ;
  assign new_n5354 = ~new_n5336 & new_n5353 ;
  assign new_n5355 = new_n3169 & ~new_n5354 ;
  assign new_n5356 = ~new_n3160 & new_n4530 ;
  assign new_n5357 = lo1403 & new_n3246 ;
  assign new_n5358 = lo1392 & new_n3254 ;
  assign new_n5359 = lo0844 & new_n3258 ;
  assign new_n5360 = ~new_n5358 & ~new_n5359 ;
  assign new_n5361 = ~new_n5357 & new_n5360 ;
  assign new_n5362 = lo1402 & new_n3267 ;
  assign new_n5363 = lo1404 & new_n3270 ;
  assign new_n5364 = lo0843 & new_n3274 ;
  assign new_n5365 = ~new_n5363 & ~new_n5364 ;
  assign new_n5366 = ~new_n5362 & new_n5365 ;
  assign new_n5367 = ~new_n3265 & new_n5366 ;
  assign new_n5368 = new_n5361 & new_n5367 ;
  assign new_n5369 = ~new_n5356 & new_n5368 ;
  assign new_n5370 = ~new_n5355 & new_n5369 ;
  assign new_n5371 = new_n3141 & ~new_n5370 ;
  assign new_n5372 = new_n3140 & ~new_n5371 ;
  assign new_n5373 = ~new_n3121 & ~new_n5372 ;
  assign new_n5374 = new_n3121 & new_n5372 ;
  assign new_n5375 = ~new_n5373 & ~new_n5374 ;
  assign new_n5376 = lo0837 & ~new_n5375 ;
  assign new_n5377 = ~lo0837 & new_n5373 ;
  assign new_n5378 = new_n3121 & new_n4530 ;
  assign new_n5379 = ~new_n5372 & new_n5378 ;
  assign new_n5380 = ~new_n5377 & ~new_n5379 ;
  assign new_n5381 = ~new_n5376 & new_n5380 ;
  assign new_n5382 = ~new_n3112 & new_n5381 ;
  assign new_n5383 = new_n3112 & ~new_n5381 ;
  assign new_n5384 = ~new_n5382 & ~new_n5383 ;
  assign new_n5385 = ~new_n3549 & new_n3737 ;
  assign new_n5386 = lo0076 & new_n2490 ;
  assign new_n5387 = lo0075 & new_n2493 ;
  assign new_n5388 = ~new_n2492 & ~new_n5387 ;
  assign new_n5389 = ~new_n5386 & new_n5388 ;
  assign new_n5390 = ~lo0249 & ~new_n5389 ;
  assign new_n5391 = lo0249 & new_n5389 ;
  assign new_n5392 = ~new_n5390 & ~new_n5391 ;
  assign new_n5393 = lo0074 & ~new_n5392 ;
  assign new_n5394 = ~lo0074 & new_n5390 ;
  assign new_n5395 = lo0077 & lo0249 ;
  assign new_n5396 = ~new_n5389 & new_n5395 ;
  assign new_n5397 = ~new_n5394 & ~new_n5396 ;
  assign new_n5398 = ~new_n5393 & new_n5397 ;
  assign new_n5399 = lo0084 & new_n2490 ;
  assign new_n5400 = lo0083 & new_n2493 ;
  assign new_n5401 = ~new_n2492 & ~new_n5400 ;
  assign new_n5402 = ~new_n5399 & new_n5401 ;
  assign new_n5403 = ~lo0249 & ~new_n5402 ;
  assign new_n5404 = lo0249 & new_n5402 ;
  assign new_n5405 = ~new_n5403 & ~new_n5404 ;
  assign new_n5406 = lo0082 & ~new_n5405 ;
  assign new_n5407 = ~lo0082 & new_n5403 ;
  assign new_n5408 = lo0085 & lo0249 ;
  assign new_n5409 = ~new_n5402 & new_n5408 ;
  assign new_n5410 = ~new_n5407 & ~new_n5409 ;
  assign new_n5411 = ~new_n5406 & new_n5410 ;
  assign new_n5412 = new_n2506 & ~new_n5411 ;
  assign new_n5413 = lo0080 & new_n2490 ;
  assign new_n5414 = lo0079 & new_n3310 ;
  assign new_n5415 = ~new_n2492 & ~new_n5414 ;
  assign new_n5416 = ~new_n5413 & new_n5415 ;
  assign new_n5417 = ~lo0250 & ~new_n5416 ;
  assign new_n5418 = lo0250 & new_n5416 ;
  assign new_n5419 = ~new_n5417 & ~new_n5418 ;
  assign new_n5420 = lo0078 & ~new_n5419 ;
  assign new_n5421 = ~lo0078 & new_n5417 ;
  assign new_n5422 = lo0081 & lo0250 ;
  assign new_n5423 = ~new_n5416 & new_n5422 ;
  assign new_n5424 = ~new_n5421 & ~new_n5423 ;
  assign new_n5425 = ~new_n5420 & new_n5424 ;
  assign new_n5426 = new_n2522 & ~new_n5425 ;
  assign new_n5427 = ~new_n2521 & ~new_n5426 ;
  assign new_n5428 = ~new_n5412 & new_n5427 ;
  assign new_n5429 = ~lo0251 & ~new_n5428 ;
  assign new_n5430 = lo0251 & new_n5428 ;
  assign new_n5431 = ~new_n5429 & ~new_n5430 ;
  assign new_n5432 = ~new_n5398 & ~new_n5431 ;
  assign new_n5433 = new_n5398 & new_n5429 ;
  assign new_n5434 = lo0088 & new_n2490 ;
  assign new_n5435 = lo0087 & new_n3310 ;
  assign new_n5436 = ~new_n2492 & ~new_n5435 ;
  assign new_n5437 = ~new_n5434 & new_n5436 ;
  assign new_n5438 = ~lo0250 & ~new_n5437 ;
  assign new_n5439 = lo0250 & new_n5437 ;
  assign new_n5440 = ~new_n5438 & ~new_n5439 ;
  assign new_n5441 = lo0086 & ~new_n5440 ;
  assign new_n5442 = ~lo0086 & new_n5438 ;
  assign new_n5443 = lo0089 & lo0250 ;
  assign new_n5444 = ~new_n5437 & new_n5443 ;
  assign new_n5445 = ~new_n5442 & ~new_n5444 ;
  assign new_n5446 = ~new_n5441 & new_n5445 ;
  assign new_n5447 = lo0251 & ~new_n5446 ;
  assign new_n5448 = ~new_n5428 & new_n5447 ;
  assign new_n5449 = ~new_n5433 & ~new_n5448 ;
  assign new_n5450 = ~new_n5432 & new_n5449 ;
  assign new_n5451 = new_n2489 & ~new_n5450 ;
  assign new_n5452 = lo0099 & new_n3367 ;
  assign new_n5453 = lo0100 & new_n3369 ;
  assign new_n5454 = ~new_n5452 & ~new_n5453 ;
  assign new_n5455 = ~new_n3366 & new_n5454 ;
  assign new_n5456 = ~new_n2483 & ~new_n5455 ;
  assign new_n5457 = lo1288 & new_n2610 ;
  assign new_n5458 = lo0763 & new_n2605 ;
  assign new_n5459 = ~new_n5457 & ~new_n5458 ;
  assign new_n5460 = lo0109 & new_n2613 ;
  assign new_n5461 = lo0102 & ~lo0103 ;
  assign new_n5462 = lo0101 & new_n5461 ;
  assign new_n5463 = lo0104 & ~new_n5461 ;
  assign new_n5464 = ~new_n5462 & ~new_n5463 ;
  assign new_n5465 = new_n2725 & ~new_n5464 ;
  assign new_n5466 = new_n2591 & new_n5465 ;
  assign new_n5467 = lo0111 & new_n2601 ;
  assign new_n5468 = ~new_n5466 & ~new_n5467 ;
  assign new_n5469 = ~new_n5460 & new_n5468 ;
  assign new_n5470 = new_n5459 & new_n5469 ;
  assign new_n5471 = ~new_n5456 & new_n5470 ;
  assign new_n5472 = ~new_n5451 & new_n5471 ;
  assign new_n5473 = new_n4180 & ~new_n5472 ;
  assign new_n5474 = ~new_n3819 & ~new_n5473 ;
  assign new_n5475 = ~new_n5385 & new_n5474 ;
  assign new_n5476 = new_n3736 & ~new_n5475 ;
  assign new_n5477 = ~new_n3736 & new_n5475 ;
  assign new_n5478 = ~new_n5476 & ~new_n5477 ;
  assign new_n5479 = ~new_n2824 & ~new_n5478 ;
  assign new_n5480 = new_n2824 & new_n5476 ;
  assign new_n5481 = lo0541 & new_n2506 ;
  assign new_n5482 = lo0540 & new_n2831 ;
  assign new_n5483 = ~new_n2521 & ~new_n5482 ;
  assign new_n5484 = ~new_n5481 & new_n5483 ;
  assign new_n5485 = ~lo0252 & ~new_n5484 ;
  assign new_n5486 = lo0252 & new_n5484 ;
  assign new_n5487 = ~new_n5485 & ~new_n5486 ;
  assign new_n5488 = lo0539 & ~new_n5487 ;
  assign new_n5489 = ~lo0539 & new_n5485 ;
  assign new_n5490 = lo0252 & lo0542 ;
  assign new_n5491 = ~new_n5484 & new_n5490 ;
  assign new_n5492 = ~new_n5489 & ~new_n5491 ;
  assign new_n5493 = ~new_n5488 & new_n5492 ;
  assign new_n5494 = lo0549 & new_n2506 ;
  assign new_n5495 = lo0548 & new_n2522 ;
  assign new_n5496 = ~new_n2521 & ~new_n5495 ;
  assign new_n5497 = ~new_n5494 & new_n5496 ;
  assign new_n5498 = ~lo0251 & ~new_n5497 ;
  assign new_n5499 = lo0251 & new_n5497 ;
  assign new_n5500 = ~new_n5498 & ~new_n5499 ;
  assign new_n5501 = lo0547 & ~new_n5500 ;
  assign new_n5502 = ~lo0547 & new_n5498 ;
  assign new_n5503 = lo0251 & lo0550 ;
  assign new_n5504 = ~new_n5497 & new_n5503 ;
  assign new_n5505 = ~new_n5502 & ~new_n5504 ;
  assign new_n5506 = ~new_n5501 & new_n5505 ;
  assign new_n5507 = new_n2490 & ~new_n5506 ;
  assign new_n5508 = lo0545 & new_n2506 ;
  assign new_n5509 = lo0544 & new_n2522 ;
  assign new_n5510 = ~new_n2521 & ~new_n5509 ;
  assign new_n5511 = ~new_n5508 & new_n5510 ;
  assign new_n5512 = ~lo0251 & ~new_n5511 ;
  assign new_n5513 = lo0251 & new_n5511 ;
  assign new_n5514 = ~new_n5512 & ~new_n5513 ;
  assign new_n5515 = lo0543 & ~new_n5514 ;
  assign new_n5516 = ~lo0543 & new_n5512 ;
  assign new_n5517 = lo0251 & lo0546 ;
  assign new_n5518 = ~new_n5511 & new_n5517 ;
  assign new_n5519 = ~new_n5516 & ~new_n5518 ;
  assign new_n5520 = ~new_n5515 & new_n5519 ;
  assign new_n5521 = new_n3310 & ~new_n5520 ;
  assign new_n5522 = ~new_n2492 & ~new_n5521 ;
  assign new_n5523 = ~new_n5507 & new_n5522 ;
  assign new_n5524 = ~lo0250 & ~new_n5523 ;
  assign new_n5525 = lo0250 & new_n5523 ;
  assign new_n5526 = ~new_n5524 & ~new_n5525 ;
  assign new_n5527 = ~new_n5493 & ~new_n5526 ;
  assign new_n5528 = new_n5493 & new_n5524 ;
  assign new_n5529 = lo0553 & new_n2506 ;
  assign new_n5530 = lo0552 & new_n2831 ;
  assign new_n5531 = ~new_n2521 & ~new_n5530 ;
  assign new_n5532 = ~new_n5529 & new_n5531 ;
  assign new_n5533 = ~lo0252 & ~new_n5532 ;
  assign new_n5534 = lo0252 & new_n5532 ;
  assign new_n5535 = ~new_n5533 & ~new_n5534 ;
  assign new_n5536 = lo0551 & ~new_n5535 ;
  assign new_n5537 = ~lo0551 & new_n5533 ;
  assign new_n5538 = lo0252 & lo0554 ;
  assign new_n5539 = ~new_n5532 & new_n5538 ;
  assign new_n5540 = ~new_n5537 & ~new_n5539 ;
  assign new_n5541 = ~new_n5536 & new_n5540 ;
  assign new_n5542 = lo0250 & ~new_n5541 ;
  assign new_n5543 = ~new_n5523 & new_n5542 ;
  assign new_n5544 = ~new_n5528 & ~new_n5543 ;
  assign new_n5545 = ~new_n5527 & new_n5544 ;
  assign new_n5546 = new_n2489 & ~new_n5545 ;
  assign new_n5547 = lo0091 & lo0555 ;
  assign new_n5548 = ~new_n2715 & ~new_n5547 ;
  assign new_n5549 = lo0090 & ~new_n5548 ;
  assign new_n5550 = ~new_n2483 & new_n5549 ;
  assign new_n5551 = lo0556 & new_n2601 ;
  assign new_n5552 = lo0558 & new_n2605 ;
  assign new_n5553 = ~new_n5551 & ~new_n5552 ;
  assign new_n5554 = lo0557 & new_n2613 ;
  assign new_n5555 = lo1329 & new_n2610 ;
  assign new_n5556 = ~new_n5554 & ~new_n5555 ;
  assign new_n5557 = new_n5553 & new_n5556 ;
  assign new_n5558 = ~new_n2729 & new_n5557 ;
  assign new_n5559 = ~new_n5550 & new_n5558 ;
  assign new_n5560 = ~new_n5546 & new_n5559 ;
  assign new_n5561 = ~new_n3736 & ~new_n5560 ;
  assign new_n5562 = ~new_n5475 & new_n5561 ;
  assign new_n5563 = ~new_n5480 & ~new_n5562 ;
  assign new_n5564 = ~new_n5479 & new_n5563 ;
  assign new_n5565 = ~lo0298 & ~new_n5564 ;
  assign new_n5566 = new_n3914 & ~new_n4097 ;
  assign new_n5567 = ~lo0297 & ~new_n4541 ;
  assign new_n5568 = ~new_n5566 & ~new_n5567 ;
  assign new_n5569 = lo0298 & ~new_n5568 ;
  assign new_n5570 = ~new_n5565 & ~new_n5569 ;
  assign new_n5571 = new_n3102 & ~new_n5570 ;
  assign new_n5572 = ~new_n3102 & ~new_n4818 ;
  assign new_n5573 = ~new_n5571 & ~new_n5572 ;
  assign new_n5574 = lo0725 & new_n3186 ;
  assign new_n5575 = lo0724 & new_n3559 ;
  assign new_n5576 = ~new_n3201 & ~new_n5575 ;
  assign new_n5577 = ~new_n5574 & new_n5576 ;
  assign new_n5578 = ~lo0065 & ~new_n5577 ;
  assign new_n5579 = lo0065 & new_n5577 ;
  assign new_n5580 = ~new_n5578 & ~new_n5579 ;
  assign new_n5581 = lo0723 & ~new_n5580 ;
  assign new_n5582 = ~lo0723 & new_n5578 ;
  assign new_n5583 = lo0065 & lo0726 ;
  assign new_n5584 = ~new_n5577 & new_n5583 ;
  assign new_n5585 = ~new_n5582 & ~new_n5584 ;
  assign new_n5586 = ~new_n5581 & new_n5585 ;
  assign new_n5587 = lo0733 & new_n3186 ;
  assign new_n5588 = lo0732 & new_n3202 ;
  assign new_n5589 = ~new_n3201 & ~new_n5588 ;
  assign new_n5590 = ~new_n5587 & new_n5589 ;
  assign new_n5591 = ~lo0063 & ~new_n5590 ;
  assign new_n5592 = lo0063 & new_n5590 ;
  assign new_n5593 = ~new_n5591 & ~new_n5592 ;
  assign new_n5594 = lo0731 & ~new_n5593 ;
  assign new_n5595 = ~lo0731 & new_n5591 ;
  assign new_n5596 = lo0063 & lo0734 ;
  assign new_n5597 = ~new_n5590 & new_n5596 ;
  assign new_n5598 = ~new_n5595 & ~new_n5597 ;
  assign new_n5599 = ~new_n5594 & new_n5598 ;
  assign new_n5600 = new_n3170 & ~new_n5599 ;
  assign new_n5601 = lo0729 & new_n3186 ;
  assign new_n5602 = lo0728 & new_n3202 ;
  assign new_n5603 = ~new_n3201 & ~new_n5602 ;
  assign new_n5604 = ~new_n5601 & new_n5603 ;
  assign new_n5605 = ~lo0063 & ~new_n5604 ;
  assign new_n5606 = lo0063 & new_n5604 ;
  assign new_n5607 = ~new_n5605 & ~new_n5606 ;
  assign new_n5608 = lo0727 & ~new_n5607 ;
  assign new_n5609 = ~lo0727 & new_n5605 ;
  assign new_n5610 = lo0063 & lo0730 ;
  assign new_n5611 = ~new_n5604 & new_n5610 ;
  assign new_n5612 = ~new_n5609 & ~new_n5611 ;
  assign new_n5613 = ~new_n5608 & new_n5612 ;
  assign new_n5614 = new_n3204 & ~new_n5613 ;
  assign new_n5615 = ~new_n3172 & ~new_n5614 ;
  assign new_n5616 = ~new_n5600 & new_n5615 ;
  assign new_n5617 = ~lo0061 & ~new_n5616 ;
  assign new_n5618 = lo0061 & new_n5616 ;
  assign new_n5619 = ~new_n5617 & ~new_n5618 ;
  assign new_n5620 = ~new_n5586 & ~new_n5619 ;
  assign new_n5621 = new_n5586 & new_n5617 ;
  assign new_n5622 = lo0737 & new_n3186 ;
  assign new_n5623 = lo0736 & new_n3559 ;
  assign new_n5624 = ~new_n3201 & ~new_n5623 ;
  assign new_n5625 = ~new_n5622 & new_n5624 ;
  assign new_n5626 = ~lo0065 & ~new_n5625 ;
  assign new_n5627 = lo0065 & new_n5625 ;
  assign new_n5628 = ~new_n5626 & ~new_n5627 ;
  assign new_n5629 = lo0735 & ~new_n5628 ;
  assign new_n5630 = ~lo0735 & new_n5626 ;
  assign new_n5631 = lo0065 & lo0738 ;
  assign new_n5632 = ~new_n5625 & new_n5631 ;
  assign new_n5633 = ~new_n5630 & ~new_n5632 ;
  assign new_n5634 = ~new_n5629 & new_n5633 ;
  assign new_n5635 = lo0061 & ~new_n5634 ;
  assign new_n5636 = ~new_n5616 & new_n5635 ;
  assign new_n5637 = ~new_n5621 & ~new_n5636 ;
  assign new_n5638 = ~new_n5620 & new_n5637 ;
  assign new_n5639 = new_n3169 & ~new_n5638 ;
  assign new_n5640 = ~new_n3160 & new_n4807 ;
  assign new_n5641 = lo1418 & new_n3246 ;
  assign new_n5642 = lo1359 & new_n3254 ;
  assign new_n5643 = lo0740 & new_n3258 ;
  assign new_n5644 = ~new_n5642 & ~new_n5643 ;
  assign new_n5645 = ~new_n5641 & new_n5644 ;
  assign new_n5646 = lo1417 & new_n3267 ;
  assign new_n5647 = lo1419 & new_n3270 ;
  assign new_n5648 = lo0739 & new_n3274 ;
  assign new_n5649 = ~new_n5647 & ~new_n5648 ;
  assign new_n5650 = ~new_n5646 & new_n5649 ;
  assign new_n5651 = ~new_n3265 & new_n5650 ;
  assign new_n5652 = new_n5645 & new_n5651 ;
  assign new_n5653 = ~new_n5640 & new_n5652 ;
  assign new_n5654 = ~new_n5639 & new_n5653 ;
  assign new_n5655 = new_n3141 & ~new_n5654 ;
  assign new_n5656 = new_n3140 & ~new_n5655 ;
  assign new_n5657 = ~new_n3121 & ~new_n5656 ;
  assign new_n5658 = new_n3121 & new_n5656 ;
  assign new_n5659 = ~new_n5657 & ~new_n5658 ;
  assign new_n5660 = lo0733 & ~new_n5659 ;
  assign new_n5661 = ~lo0733 & new_n5657 ;
  assign new_n5662 = new_n3121 & new_n4807 ;
  assign new_n5663 = ~new_n5656 & new_n5662 ;
  assign new_n5664 = ~new_n5661 & ~new_n5663 ;
  assign new_n5665 = ~new_n5660 & new_n5664 ;
  assign new_n5666 = ~new_n3112 & new_n5665 ;
  assign new_n5667 = new_n3112 & ~new_n5665 ;
  assign new_n5668 = ~new_n5666 & ~new_n5667 ;
  assign new_n5669 = lo0297 & lo0298 ;
  assign new_n5670 = lo0298 & ~new_n3736 ;
  assign new_n5671 = lo0299 & ~new_n5670 ;
  assign new_n5672 = new_n5669 & ~new_n5671 ;
  assign new_n5673 = new_n5669 & new_n5670 ;
  assign new_n5674 = lo0384 & new_n2506 ;
  assign new_n5675 = lo0383 & new_n2831 ;
  assign new_n5676 = ~new_n2521 & ~new_n5675 ;
  assign new_n5677 = ~new_n5674 & new_n5676 ;
  assign new_n5678 = ~lo0252 & ~new_n5677 ;
  assign new_n5679 = lo0252 & new_n5677 ;
  assign new_n5680 = ~new_n5678 & ~new_n5679 ;
  assign new_n5681 = lo0382 & ~new_n5680 ;
  assign new_n5682 = ~lo0382 & new_n5678 ;
  assign new_n5683 = lo0252 & lo0385 ;
  assign new_n5684 = ~new_n5677 & new_n5683 ;
  assign new_n5685 = ~new_n5682 & ~new_n5684 ;
  assign new_n5686 = ~new_n5681 & new_n5685 ;
  assign new_n5687 = lo0392 & new_n2506 ;
  assign new_n5688 = lo0391 & new_n2831 ;
  assign new_n5689 = ~new_n2521 & ~new_n5688 ;
  assign new_n5690 = ~new_n5687 & new_n5689 ;
  assign new_n5691 = ~lo0252 & ~new_n5690 ;
  assign new_n5692 = lo0252 & new_n5690 ;
  assign new_n5693 = ~new_n5691 & ~new_n5692 ;
  assign new_n5694 = lo0390 & ~new_n5693 ;
  assign new_n5695 = ~lo0390 & new_n5691 ;
  assign new_n5696 = lo0252 & lo0393 ;
  assign new_n5697 = ~new_n5690 & new_n5696 ;
  assign new_n5698 = ~new_n5695 & ~new_n5697 ;
  assign new_n5699 = ~new_n5694 & new_n5698 ;
  assign new_n5700 = new_n2490 & ~new_n5699 ;
  assign new_n5701 = lo0388 & new_n2506 ;
  assign new_n5702 = lo0387 & new_n2522 ;
  assign new_n5703 = ~new_n2521 & ~new_n5702 ;
  assign new_n5704 = ~new_n5701 & new_n5703 ;
  assign new_n5705 = ~lo0251 & ~new_n5704 ;
  assign new_n5706 = lo0251 & new_n5704 ;
  assign new_n5707 = ~new_n5705 & ~new_n5706 ;
  assign new_n5708 = lo0386 & ~new_n5707 ;
  assign new_n5709 = ~lo0386 & new_n5705 ;
  assign new_n5710 = lo0251 & lo0389 ;
  assign new_n5711 = ~new_n5704 & new_n5710 ;
  assign new_n5712 = ~new_n5709 & ~new_n5711 ;
  assign new_n5713 = ~new_n5708 & new_n5712 ;
  assign new_n5714 = new_n2493 & ~new_n5713 ;
  assign new_n5715 = ~new_n2492 & ~new_n5714 ;
  assign new_n5716 = ~new_n5700 & new_n5715 ;
  assign new_n5717 = ~lo0249 & ~new_n5716 ;
  assign new_n5718 = lo0249 & new_n5716 ;
  assign new_n5719 = ~new_n5717 & ~new_n5718 ;
  assign new_n5720 = ~new_n5686 & ~new_n5719 ;
  assign new_n5721 = new_n5686 & new_n5717 ;
  assign new_n5722 = lo0396 & new_n2506 ;
  assign new_n5723 = lo0395 & new_n2522 ;
  assign new_n5724 = ~new_n2521 & ~new_n5723 ;
  assign new_n5725 = ~new_n5722 & new_n5724 ;
  assign new_n5726 = ~lo0251 & ~new_n5725 ;
  assign new_n5727 = lo0251 & new_n5725 ;
  assign new_n5728 = ~new_n5726 & ~new_n5727 ;
  assign new_n5729 = lo0394 & ~new_n5728 ;
  assign new_n5730 = ~lo0394 & new_n5726 ;
  assign new_n5731 = lo0251 & lo0397 ;
  assign new_n5732 = ~new_n5725 & new_n5731 ;
  assign new_n5733 = ~new_n5730 & ~new_n5732 ;
  assign new_n5734 = ~new_n5729 & new_n5733 ;
  assign new_n5735 = lo0249 & ~new_n5734 ;
  assign new_n5736 = ~new_n5716 & new_n5735 ;
  assign new_n5737 = ~new_n5721 & ~new_n5736 ;
  assign new_n5738 = ~new_n5720 & new_n5737 ;
  assign new_n5739 = new_n2489 & ~new_n5738 ;
  assign new_n5740 = lo0098 & new_n3367 ;
  assign new_n5741 = lo0094 & new_n3369 ;
  assign new_n5742 = ~new_n5740 & ~new_n5741 ;
  assign new_n5743 = ~new_n3366 & new_n5742 ;
  assign new_n5744 = ~new_n2483 & ~new_n5743 ;
  assign new_n5745 = ~lo0102 & ~lo0222 ;
  assign new_n5746 = ~lo0103 & ~new_n5745 ;
  assign new_n5747 = ~lo0102 & new_n5746 ;
  assign new_n5748 = ~lo0105 & ~new_n5747 ;
  assign new_n5749 = lo0104 & ~new_n5748 ;
  assign new_n5750 = lo0101 & ~new_n5746 ;
  assign new_n5751 = lo0398 & new_n5746 ;
  assign new_n5752 = ~new_n5750 & ~new_n5751 ;
  assign new_n5753 = new_n5748 & ~new_n5752 ;
  assign new_n5754 = ~new_n5749 & ~new_n5753 ;
  assign new_n5755 = new_n2724 & ~new_n5754 ;
  assign new_n5756 = new_n2591 & new_n5755 ;
  assign new_n5757 = lo0399 & new_n2601 ;
  assign new_n5758 = lo0559 & new_n2605 ;
  assign new_n5759 = ~new_n5757 & ~new_n5758 ;
  assign new_n5760 = lo1309 & new_n2610 ;
  assign new_n5761 = lo0400 & new_n2613 ;
  assign new_n5762 = ~new_n5760 & ~new_n5761 ;
  assign new_n5763 = new_n5759 & new_n5762 ;
  assign new_n5764 = ~new_n5756 & new_n5763 ;
  assign new_n5765 = ~new_n5744 & new_n5764 ;
  assign new_n5766 = ~new_n5739 & new_n5765 ;
  assign new_n5767 = new_n3737 & ~new_n3908 ;
  assign new_n5768 = ~new_n3549 & new_n3820 ;
  assign new_n5769 = ~new_n3819 & ~new_n5768 ;
  assign new_n5770 = ~new_n5767 & new_n5769 ;
  assign new_n5771 = ~new_n3735 & ~new_n5770 ;
  assign new_n5772 = new_n3735 & new_n5770 ;
  assign new_n5773 = ~new_n5771 & ~new_n5772 ;
  assign new_n5774 = ~new_n5766 & ~new_n5773 ;
  assign new_n5775 = new_n5766 & new_n5771 ;
  assign new_n5776 = ~new_n2910 & new_n3735 ;
  assign new_n5777 = ~new_n5770 & new_n5776 ;
  assign new_n5778 = ~new_n5775 & ~new_n5777 ;
  assign new_n5779 = ~new_n5774 & new_n5778 ;
  assign new_n5780 = new_n5673 & new_n5779 ;
  assign new_n5781 = ~new_n5669 & ~new_n5670 ;
  assign new_n5782 = ~new_n5673 & ~new_n5781 ;
  assign new_n5783 = ~new_n5779 & ~new_n5782 ;
  assign new_n5784 = ~new_n5669 & new_n5670 ;
  assign new_n5785 = ~new_n4818 & new_n5784 ;
  assign new_n5786 = ~new_n5783 & ~new_n5785 ;
  assign new_n5787 = ~new_n5780 & new_n5786 ;
  assign new_n5788 = ~new_n5672 & ~new_n5787 ;
  assign new_n5789 = new_n5672 & new_n5787 ;
  assign new_n5790 = ~new_n5788 & ~new_n5789 ;
  assign new_n5791 = ~new_n4541 & ~new_n5790 ;
  assign new_n5792 = new_n4541 & new_n5788 ;
  assign new_n5793 = ~new_n2739 & new_n5672 ;
  assign new_n5794 = ~new_n5787 & new_n5793 ;
  assign new_n5795 = ~new_n5792 & ~new_n5794 ;
  assign new_n5796 = ~new_n5791 & new_n5795 ;
  assign new_n5797 = new_n3102 & ~new_n5796 ;
  assign new_n5798 = ~new_n2824 & ~new_n3102 ;
  assign new_n5799 = ~new_n5797 & ~new_n5798 ;
  assign new_n5800 = lo0605 & new_n3170 ;
  assign new_n5801 = lo0604 & new_n3173 ;
  assign new_n5802 = ~new_n3172 & ~new_n5801 ;
  assign new_n5803 = ~new_n5800 & new_n5802 ;
  assign new_n5804 = ~lo0059 & ~new_n5803 ;
  assign new_n5805 = lo0059 & new_n5803 ;
  assign new_n5806 = ~new_n5804 & ~new_n5805 ;
  assign new_n5807 = lo0603 & ~new_n5806 ;
  assign new_n5808 = ~lo0603 & new_n5804 ;
  assign new_n5809 = lo0059 & lo0606 ;
  assign new_n5810 = ~new_n5803 & new_n5809 ;
  assign new_n5811 = ~new_n5808 & ~new_n5810 ;
  assign new_n5812 = ~new_n5807 & new_n5811 ;
  assign new_n5813 = lo0613 & new_n3170 ;
  assign new_n5814 = lo0612 & new_n3173 ;
  assign new_n5815 = ~new_n3172 & ~new_n5814 ;
  assign new_n5816 = ~new_n5813 & new_n5815 ;
  assign new_n5817 = ~lo0059 & ~new_n5816 ;
  assign new_n5818 = lo0059 & new_n5816 ;
  assign new_n5819 = ~new_n5817 & ~new_n5818 ;
  assign new_n5820 = lo0611 & ~new_n5819 ;
  assign new_n5821 = ~lo0611 & new_n5817 ;
  assign new_n5822 = lo0059 & lo0614 ;
  assign new_n5823 = ~new_n5816 & new_n5822 ;
  assign new_n5824 = ~new_n5821 & ~new_n5823 ;
  assign new_n5825 = ~new_n5820 & new_n5824 ;
  assign new_n5826 = new_n3186 & ~new_n5825 ;
  assign new_n5827 = lo0609 & new_n3170 ;
  assign new_n5828 = lo0608 & new_n3204 ;
  assign new_n5829 = ~new_n3172 & ~new_n5828 ;
  assign new_n5830 = ~new_n5827 & new_n5829 ;
  assign new_n5831 = ~lo0061 & ~new_n5830 ;
  assign new_n5832 = lo0061 & new_n5830 ;
  assign new_n5833 = ~new_n5831 & ~new_n5832 ;
  assign new_n5834 = lo0607 & ~new_n5833 ;
  assign new_n5835 = ~lo0607 & new_n5831 ;
  assign new_n5836 = lo0061 & lo0610 ;
  assign new_n5837 = ~new_n5830 & new_n5836 ;
  assign new_n5838 = ~new_n5835 & ~new_n5837 ;
  assign new_n5839 = ~new_n5834 & new_n5838 ;
  assign new_n5840 = new_n3202 & ~new_n5839 ;
  assign new_n5841 = ~new_n3201 & ~new_n5840 ;
  assign new_n5842 = ~new_n5826 & new_n5841 ;
  assign new_n5843 = ~lo0063 & ~new_n5842 ;
  assign new_n5844 = lo0063 & new_n5842 ;
  assign new_n5845 = ~new_n5843 & ~new_n5844 ;
  assign new_n5846 = ~new_n5812 & ~new_n5845 ;
  assign new_n5847 = new_n5812 & new_n5843 ;
  assign new_n5848 = lo0617 & new_n3170 ;
  assign new_n5849 = lo0616 & new_n3204 ;
  assign new_n5850 = ~new_n3172 & ~new_n5849 ;
  assign new_n5851 = ~new_n5848 & new_n5850 ;
  assign new_n5852 = ~lo0061 & ~new_n5851 ;
  assign new_n5853 = lo0061 & new_n5851 ;
  assign new_n5854 = ~new_n5852 & ~new_n5853 ;
  assign new_n5855 = lo0615 & ~new_n5854 ;
  assign new_n5856 = ~lo0615 & new_n5852 ;
  assign new_n5857 = lo0061 & lo0618 ;
  assign new_n5858 = ~new_n5851 & new_n5857 ;
  assign new_n5859 = ~new_n5856 & ~new_n5858 ;
  assign new_n5860 = ~new_n5855 & new_n5859 ;
  assign new_n5861 = lo0063 & ~new_n5860 ;
  assign new_n5862 = ~new_n5842 & new_n5861 ;
  assign new_n5863 = ~new_n5847 & ~new_n5862 ;
  assign new_n5864 = ~new_n5846 & new_n5863 ;
  assign new_n5865 = new_n3169 & ~new_n5864 ;
  assign new_n5866 = new_n2813 & ~new_n3160 ;
  assign new_n5867 = lo1394 & new_n3246 ;
  assign new_n5868 = lo1344 & new_n3254 ;
  assign new_n5869 = lo0620 & new_n3258 ;
  assign new_n5870 = ~new_n5868 & ~new_n5869 ;
  assign new_n5871 = ~new_n5867 & new_n5870 ;
  assign new_n5872 = lo1393 & new_n3267 ;
  assign new_n5873 = lo1395 & new_n3270 ;
  assign new_n5874 = lo0619 & new_n3274 ;
  assign new_n5875 = ~new_n5873 & ~new_n5874 ;
  assign new_n5876 = ~new_n5872 & new_n5875 ;
  assign new_n5877 = ~new_n3265 & new_n5876 ;
  assign new_n5878 = new_n5871 & new_n5877 ;
  assign new_n5879 = ~new_n5866 & new_n5878 ;
  assign new_n5880 = ~new_n5865 & new_n5879 ;
  assign new_n5881 = new_n3141 & ~new_n5880 ;
  assign new_n5882 = new_n3140 & ~new_n5881 ;
  assign new_n5883 = ~new_n3121 & ~new_n5882 ;
  assign new_n5884 = new_n3121 & new_n5882 ;
  assign new_n5885 = ~new_n5883 & ~new_n5884 ;
  assign new_n5886 = lo0613 & ~new_n5885 ;
  assign new_n5887 = ~lo0613 & new_n5883 ;
  assign new_n5888 = new_n2813 & new_n3121 ;
  assign new_n5889 = ~new_n5882 & new_n5888 ;
  assign new_n5890 = ~new_n5887 & ~new_n5889 ;
  assign new_n5891 = ~new_n5886 & new_n5890 ;
  assign new_n5892 = ~new_n3112 & new_n5891 ;
  assign new_n5893 = new_n3112 & ~new_n5891 ;
  assign new_n5894 = ~new_n5892 & ~new_n5893 ;
  assign new_n5895 = new_n3737 & ~new_n4268 ;
  assign new_n5896 = lo0501 & new_n2490 ;
  assign new_n5897 = lo0500 & new_n2493 ;
  assign new_n5898 = ~new_n2492 & ~new_n5897 ;
  assign new_n5899 = ~new_n5896 & new_n5898 ;
  assign new_n5900 = ~lo0249 & ~new_n5899 ;
  assign new_n5901 = lo0249 & new_n5899 ;
  assign new_n5902 = ~new_n5900 & ~new_n5901 ;
  assign new_n5903 = lo0499 & ~new_n5902 ;
  assign new_n5904 = ~lo0499 & new_n5900 ;
  assign new_n5905 = lo0249 & lo0502 ;
  assign new_n5906 = ~new_n5899 & new_n5905 ;
  assign new_n5907 = ~new_n5904 & ~new_n5906 ;
  assign new_n5908 = ~new_n5903 & new_n5907 ;
  assign new_n5909 = lo0498 & new_n2490 ;
  assign new_n5910 = lo0508 & new_n3310 ;
  assign new_n5911 = ~new_n2492 & ~new_n5910 ;
  assign new_n5912 = ~new_n5909 & new_n5911 ;
  assign new_n5913 = ~lo0250 & ~new_n5912 ;
  assign new_n5914 = lo0250 & new_n5912 ;
  assign new_n5915 = ~new_n5913 & ~new_n5914 ;
  assign new_n5916 = lo0507 & ~new_n5915 ;
  assign new_n5917 = ~lo0507 & new_n5913 ;
  assign new_n5918 = lo0250 & lo0509 ;
  assign new_n5919 = ~new_n5912 & new_n5918 ;
  assign new_n5920 = ~new_n5917 & ~new_n5919 ;
  assign new_n5921 = ~new_n5916 & new_n5920 ;
  assign new_n5922 = new_n2506 & ~new_n5921 ;
  assign new_n5923 = lo0505 & new_n2490 ;
  assign new_n5924 = lo0504 & new_n3310 ;
  assign new_n5925 = ~new_n2492 & ~new_n5924 ;
  assign new_n5926 = ~new_n5923 & new_n5925 ;
  assign new_n5927 = ~lo0250 & ~new_n5926 ;
  assign new_n5928 = lo0250 & new_n5926 ;
  assign new_n5929 = ~new_n5927 & ~new_n5928 ;
  assign new_n5930 = lo0503 & ~new_n5929 ;
  assign new_n5931 = ~lo0503 & new_n5927 ;
  assign new_n5932 = lo0250 & lo0506 ;
  assign new_n5933 = ~new_n5926 & new_n5932 ;
  assign new_n5934 = ~new_n5931 & ~new_n5933 ;
  assign new_n5935 = ~new_n5930 & new_n5934 ;
  assign new_n5936 = new_n2831 & ~new_n5935 ;
  assign new_n5937 = ~new_n2521 & ~new_n5936 ;
  assign new_n5938 = ~new_n5922 & new_n5937 ;
  assign new_n5939 = ~lo0252 & ~new_n5938 ;
  assign new_n5940 = lo0252 & new_n5938 ;
  assign new_n5941 = ~new_n5939 & ~new_n5940 ;
  assign new_n5942 = ~new_n5908 & ~new_n5941 ;
  assign new_n5943 = new_n5908 & new_n5939 ;
  assign new_n5944 = lo0512 & new_n2490 ;
  assign new_n5945 = lo0511 & new_n2493 ;
  assign new_n5946 = ~new_n2492 & ~new_n5945 ;
  assign new_n5947 = ~new_n5944 & new_n5946 ;
  assign new_n5948 = ~lo0249 & ~new_n5947 ;
  assign new_n5949 = lo0249 & new_n5947 ;
  assign new_n5950 = ~new_n5948 & ~new_n5949 ;
  assign new_n5951 = lo0510 & ~new_n5950 ;
  assign new_n5952 = ~lo0510 & new_n5948 ;
  assign new_n5953 = lo0249 & lo0513 ;
  assign new_n5954 = ~new_n5947 & new_n5953 ;
  assign new_n5955 = ~new_n5952 & ~new_n5954 ;
  assign new_n5956 = ~new_n5951 & new_n5955 ;
  assign new_n5957 = lo0252 & ~new_n5956 ;
  assign new_n5958 = ~new_n5938 & new_n5957 ;
  assign new_n5959 = ~new_n5943 & ~new_n5958 ;
  assign new_n5960 = ~new_n5942 & new_n5959 ;
  assign new_n5961 = new_n2489 & ~new_n5960 ;
  assign new_n5962 = lo0435 & new_n2565 ;
  assign new_n5963 = new_n2569 & new_n5962 ;
  assign new_n5964 = lo0274 & ~new_n2565 ;
  assign new_n5965 = new_n2569 & new_n5964 ;
  assign new_n5966 = ~new_n2572 & ~new_n5965 ;
  assign new_n5967 = ~new_n5963 & new_n5966 ;
  assign new_n5968 = new_n2569 & ~new_n5967 ;
  assign new_n5969 = ~new_n2569 & new_n5967 ;
  assign new_n5970 = ~new_n5968 & ~new_n5969 ;
  assign new_n5971 = lo0436 & ~new_n5970 ;
  assign new_n5972 = ~lo0436 & new_n5968 ;
  assign new_n5973 = lo0514 & ~new_n2569 ;
  assign new_n5974 = ~new_n5967 & new_n5973 ;
  assign new_n5975 = ~new_n5972 & ~new_n5974 ;
  assign new_n5976 = ~new_n5971 & new_n5975 ;
  assign new_n5977 = lo0090 & ~new_n5976 ;
  assign new_n5978 = ~new_n2483 & new_n5977 ;
  assign new_n5979 = lo0101 & ~new_n5748 ;
  assign new_n5980 = lo0398 & ~new_n5746 ;
  assign new_n5981 = lo0224 & new_n5746 ;
  assign new_n5982 = ~new_n5980 & ~new_n5981 ;
  assign new_n5983 = new_n5748 & ~new_n5982 ;
  assign new_n5984 = ~new_n5979 & ~new_n5983 ;
  assign new_n5985 = new_n2724 & ~new_n5984 ;
  assign new_n5986 = new_n2591 & new_n5985 ;
  assign new_n5987 = lo0516 & new_n2601 ;
  assign new_n5988 = lo0517 & new_n2605 ;
  assign new_n5989 = ~new_n5987 & ~new_n5988 ;
  assign new_n5990 = lo1322 & new_n2610 ;
  assign new_n5991 = lo0515 & new_n2613 ;
  assign new_n5992 = ~new_n5990 & ~new_n5991 ;
  assign new_n5993 = new_n5989 & new_n5992 ;
  assign new_n5994 = ~new_n5986 & new_n5993 ;
  assign new_n5995 = ~new_n5978 & new_n5994 ;
  assign new_n5996 = ~new_n5961 & new_n5995 ;
  assign new_n5997 = new_n4180 & ~new_n5996 ;
  assign new_n5998 = ~new_n3819 & ~new_n5997 ;
  assign new_n5999 = ~new_n5895 & new_n5998 ;
  assign new_n6000 = new_n3736 & ~new_n5999 ;
  assign new_n6001 = ~new_n3736 & new_n5999 ;
  assign new_n6002 = ~new_n6000 & ~new_n6001 ;
  assign new_n6003 = ~new_n3908 & ~new_n6002 ;
  assign new_n6004 = new_n3908 & new_n6000 ;
  assign new_n6005 = ~new_n3383 & ~new_n3736 ;
  assign new_n6006 = ~new_n5999 & new_n6005 ;
  assign new_n6007 = ~new_n6004 & ~new_n6006 ;
  assign new_n6008 = ~new_n6003 & new_n6007 ;
  assign new_n6009 = new_n5673 & new_n6008 ;
  assign new_n6010 = ~new_n5782 & ~new_n6008 ;
  assign new_n6011 = ~new_n2824 & new_n5784 ;
  assign new_n6012 = ~new_n6010 & ~new_n6011 ;
  assign new_n6013 = ~new_n6009 & new_n6012 ;
  assign new_n6014 = ~new_n5672 & ~new_n6013 ;
  assign new_n6015 = new_n5672 & new_n6013 ;
  assign new_n6016 = ~new_n6014 & ~new_n6015 ;
  assign new_n6017 = ~new_n4818 & ~new_n6016 ;
  assign new_n6018 = new_n4818 & new_n6014 ;
  assign new_n6019 = ~new_n3092 & new_n5672 ;
  assign new_n6020 = ~new_n6013 & new_n6019 ;
  assign new_n6021 = ~new_n6018 & ~new_n6020 ;
  assign new_n6022 = ~new_n6017 & new_n6021 ;
  assign new_n6023 = new_n3102 & ~new_n6022 ;
  assign new_n6024 = ~new_n3102 & ~new_n3549 ;
  assign new_n6025 = ~new_n6023 & ~new_n6024 ;
  assign new_n6026 = lo0260 & new_n3186 ;
  assign new_n6027 = lo0259 & new_n3559 ;
  assign new_n6028 = ~new_n3201 & ~new_n6027 ;
  assign new_n6029 = ~new_n6026 & new_n6028 ;
  assign new_n6030 = ~lo0065 & ~new_n6029 ;
  assign new_n6031 = lo0065 & new_n6029 ;
  assign new_n6032 = ~new_n6030 & ~new_n6031 ;
  assign new_n6033 = lo0258 & ~new_n6032 ;
  assign new_n6034 = ~lo0258 & new_n6030 ;
  assign new_n6035 = lo0065 & lo0261 ;
  assign new_n6036 = ~new_n6029 & new_n6035 ;
  assign new_n6037 = ~new_n6034 & ~new_n6036 ;
  assign new_n6038 = ~new_n6033 & new_n6037 ;
  assign new_n6039 = lo0268 & new_n3186 ;
  assign new_n6040 = lo0267 & new_n3559 ;
  assign new_n6041 = ~new_n3201 & ~new_n6040 ;
  assign new_n6042 = ~new_n6039 & new_n6041 ;
  assign new_n6043 = ~lo0065 & ~new_n6042 ;
  assign new_n6044 = lo0065 & new_n6042 ;
  assign new_n6045 = ~new_n6043 & ~new_n6044 ;
  assign new_n6046 = lo0266 & ~new_n6045 ;
  assign new_n6047 = ~lo0266 & new_n6043 ;
  assign new_n6048 = lo0065 & lo0269 ;
  assign new_n6049 = ~new_n6042 & new_n6048 ;
  assign new_n6050 = ~new_n6047 & ~new_n6049 ;
  assign new_n6051 = ~new_n6046 & new_n6050 ;
  assign new_n6052 = new_n3170 & ~new_n6051 ;
  assign new_n6053 = lo0264 & new_n3186 ;
  assign new_n6054 = lo0263 & new_n3202 ;
  assign new_n6055 = ~new_n3201 & ~new_n6054 ;
  assign new_n6056 = ~new_n6053 & new_n6055 ;
  assign new_n6057 = ~lo0063 & ~new_n6056 ;
  assign new_n6058 = lo0063 & new_n6056 ;
  assign new_n6059 = ~new_n6057 & ~new_n6058 ;
  assign new_n6060 = lo0262 & ~new_n6059 ;
  assign new_n6061 = ~lo0262 & new_n6057 ;
  assign new_n6062 = lo0063 & lo0265 ;
  assign new_n6063 = ~new_n6056 & new_n6062 ;
  assign new_n6064 = ~new_n6061 & ~new_n6063 ;
  assign new_n6065 = ~new_n6060 & new_n6064 ;
  assign new_n6066 = new_n3173 & ~new_n6065 ;
  assign new_n6067 = ~new_n3172 & ~new_n6066 ;
  assign new_n6068 = ~new_n6052 & new_n6067 ;
  assign new_n6069 = ~lo0059 & ~new_n6068 ;
  assign new_n6070 = lo0059 & new_n6068 ;
  assign new_n6071 = ~new_n6069 & ~new_n6070 ;
  assign new_n6072 = ~new_n6038 & ~new_n6071 ;
  assign new_n6073 = new_n6038 & new_n6069 ;
  assign new_n6074 = lo0272 & new_n3186 ;
  assign new_n6075 = lo0271 & new_n3202 ;
  assign new_n6076 = ~new_n3201 & ~new_n6075 ;
  assign new_n6077 = ~new_n6074 & new_n6076 ;
  assign new_n6078 = ~lo0063 & ~new_n6077 ;
  assign new_n6079 = lo0063 & new_n6077 ;
  assign new_n6080 = ~new_n6078 & ~new_n6079 ;
  assign new_n6081 = lo0270 & ~new_n6080 ;
  assign new_n6082 = ~lo0270 & new_n6078 ;
  assign new_n6083 = lo0063 & lo0273 ;
  assign new_n6084 = ~new_n6077 & new_n6083 ;
  assign new_n6085 = ~new_n6082 & ~new_n6084 ;
  assign new_n6086 = ~new_n6081 & new_n6085 ;
  assign new_n6087 = lo0059 & ~new_n6086 ;
  assign new_n6088 = ~new_n6068 & new_n6087 ;
  assign new_n6089 = ~new_n6073 & ~new_n6088 ;
  assign new_n6090 = ~new_n6072 & new_n6089 ;
  assign new_n6091 = new_n3169 & ~new_n6090 ;
  assign new_n6092 = ~new_n3160 & new_n3538 ;
  assign new_n6093 = lo1357 & new_n3246 ;
  assign new_n6094 = lo1303 & new_n3254 ;
  assign new_n6095 = lo0276 & new_n3258 ;
  assign new_n6096 = ~new_n6094 & ~new_n6095 ;
  assign new_n6097 = ~new_n6093 & new_n6096 ;
  assign new_n6098 = lo1356 & new_n3267 ;
  assign new_n6099 = lo1358 & new_n3270 ;
  assign new_n6100 = lo0275 & new_n3274 ;
  assign new_n6101 = ~new_n6099 & ~new_n6100 ;
  assign new_n6102 = ~new_n6098 & new_n6101 ;
  assign new_n6103 = ~new_n3265 & new_n6102 ;
  assign new_n6104 = new_n6097 & new_n6103 ;
  assign new_n6105 = ~new_n6092 & new_n6104 ;
  assign new_n6106 = ~new_n6091 & new_n6105 ;
  assign new_n6107 = new_n3141 & ~new_n6106 ;
  assign new_n6108 = new_n3140 & ~new_n6107 ;
  assign new_n6109 = ~new_n3121 & ~new_n6108 ;
  assign new_n6110 = new_n3121 & new_n6108 ;
  assign new_n6111 = ~new_n6109 & ~new_n6110 ;
  assign new_n6112 = lo0268 & ~new_n6111 ;
  assign new_n6113 = ~lo0268 & new_n6109 ;
  assign new_n6114 = new_n3121 & new_n3538 ;
  assign new_n6115 = ~new_n6108 & new_n6114 ;
  assign new_n6116 = ~new_n6113 & ~new_n6115 ;
  assign new_n6117 = ~new_n6112 & new_n6116 ;
  assign new_n6118 = ~new_n3112 & new_n6117 ;
  assign new_n6119 = new_n3112 & ~new_n6117 ;
  assign new_n6120 = ~new_n6118 & ~new_n6119 ;
  assign new_n6121 = lo0585 & new_n2506 ;
  assign new_n6122 = lo0584 & new_n2831 ;
  assign new_n6123 = ~new_n2521 & ~new_n6122 ;
  assign new_n6124 = ~new_n6121 & new_n6123 ;
  assign new_n6125 = ~lo0252 & ~new_n6124 ;
  assign new_n6126 = lo0252 & new_n6124 ;
  assign new_n6127 = ~new_n6125 & ~new_n6126 ;
  assign new_n6128 = lo0583 & ~new_n6127 ;
  assign new_n6129 = ~lo0583 & new_n6125 ;
  assign new_n6130 = lo0252 & lo0586 ;
  assign new_n6131 = ~new_n6124 & new_n6130 ;
  assign new_n6132 = ~new_n6129 & ~new_n6131 ;
  assign new_n6133 = ~new_n6128 & new_n6132 ;
  assign new_n6134 = lo0593 & new_n2506 ;
  assign new_n6135 = lo0592 & new_n2522 ;
  assign new_n6136 = ~new_n2521 & ~new_n6135 ;
  assign new_n6137 = ~new_n6134 & new_n6136 ;
  assign new_n6138 = ~lo0251 & ~new_n6137 ;
  assign new_n6139 = lo0251 & new_n6137 ;
  assign new_n6140 = ~new_n6138 & ~new_n6139 ;
  assign new_n6141 = lo0591 & ~new_n6140 ;
  assign new_n6142 = ~lo0591 & new_n6138 ;
  assign new_n6143 = lo0251 & lo0594 ;
  assign new_n6144 = ~new_n6137 & new_n6143 ;
  assign new_n6145 = ~new_n6142 & ~new_n6144 ;
  assign new_n6146 = ~new_n6141 & new_n6145 ;
  assign new_n6147 = new_n2490 & ~new_n6146 ;
  assign new_n6148 = lo0589 & new_n2506 ;
  assign new_n6149 = lo0588 & new_n2522 ;
  assign new_n6150 = ~new_n2521 & ~new_n6149 ;
  assign new_n6151 = ~new_n6148 & new_n6150 ;
  assign new_n6152 = ~lo0251 & ~new_n6151 ;
  assign new_n6153 = lo0251 & new_n6151 ;
  assign new_n6154 = ~new_n6152 & ~new_n6153 ;
  assign new_n6155 = lo0587 & ~new_n6154 ;
  assign new_n6156 = ~lo0587 & new_n6152 ;
  assign new_n6157 = lo0251 & lo0590 ;
  assign new_n6158 = ~new_n6151 & new_n6157 ;
  assign new_n6159 = ~new_n6156 & ~new_n6158 ;
  assign new_n6160 = ~new_n6155 & new_n6159 ;
  assign new_n6161 = new_n3310 & ~new_n6160 ;
  assign new_n6162 = ~new_n2492 & ~new_n6161 ;
  assign new_n6163 = ~new_n6147 & new_n6162 ;
  assign new_n6164 = ~lo0250 & ~new_n6163 ;
  assign new_n6165 = lo0250 & new_n6163 ;
  assign new_n6166 = ~new_n6164 & ~new_n6165 ;
  assign new_n6167 = ~new_n6133 & ~new_n6166 ;
  assign new_n6168 = new_n6133 & new_n6164 ;
  assign new_n6169 = lo0597 & new_n2506 ;
  assign new_n6170 = lo0596 & new_n2831 ;
  assign new_n6171 = ~new_n2521 & ~new_n6170 ;
  assign new_n6172 = ~new_n6169 & new_n6171 ;
  assign new_n6173 = ~lo0252 & ~new_n6172 ;
  assign new_n6174 = lo0252 & new_n6172 ;
  assign new_n6175 = ~new_n6173 & ~new_n6174 ;
  assign new_n6176 = lo0595 & ~new_n6175 ;
  assign new_n6177 = ~lo0595 & new_n6173 ;
  assign new_n6178 = lo0252 & lo0598 ;
  assign new_n6179 = ~new_n6172 & new_n6178 ;
  assign new_n6180 = ~new_n6177 & ~new_n6179 ;
  assign new_n6181 = ~new_n6176 & new_n6180 ;
  assign new_n6182 = lo0250 & ~new_n6181 ;
  assign new_n6183 = ~new_n6163 & new_n6182 ;
  assign new_n6184 = ~new_n6168 & ~new_n6183 ;
  assign new_n6185 = ~new_n6167 & new_n6184 ;
  assign new_n6186 = new_n2489 & ~new_n6185 ;
  assign new_n6187 = lo0534 & new_n2565 ;
  assign new_n6188 = new_n2569 & new_n6187 ;
  assign new_n6189 = lo0456 & new_n2565 ;
  assign new_n6190 = ~new_n2569 & new_n6189 ;
  assign new_n6191 = ~new_n2572 & ~new_n6190 ;
  assign new_n6192 = ~new_n6188 & new_n6191 ;
  assign new_n6193 = new_n2565 & ~new_n6192 ;
  assign new_n6194 = ~new_n2565 & new_n6192 ;
  assign new_n6195 = ~new_n6193 & ~new_n6194 ;
  assign new_n6196 = lo0377 & ~new_n6195 ;
  assign new_n6197 = ~lo0377 & new_n6193 ;
  assign new_n6198 = lo0599 & ~new_n2565 ;
  assign new_n6199 = ~new_n6192 & new_n6198 ;
  assign new_n6200 = ~new_n6197 & ~new_n6199 ;
  assign new_n6201 = ~new_n6196 & new_n6200 ;
  assign new_n6202 = lo0090 & ~new_n6201 ;
  assign new_n6203 = ~new_n2483 & new_n6202 ;
  assign new_n6204 = lo0108 & lo0221 ;
  assign new_n6205 = lo0398 & ~new_n2595 ;
  assign new_n6206 = lo0221 & new_n5461 ;
  assign new_n6207 = lo0224 & ~new_n5746 ;
  assign new_n6208 = ~new_n6206 & ~new_n6207 ;
  assign new_n6209 = ~lo0105 & ~new_n6208 ;
  assign new_n6210 = ~new_n6205 & ~new_n6209 ;
  assign new_n6211 = ~lo0108 & ~new_n6210 ;
  assign new_n6212 = ~new_n6204 & ~new_n6211 ;
  assign new_n6213 = ~lo0106 & ~lo0107 ;
  assign new_n6214 = ~new_n6212 & new_n6213 ;
  assign new_n6215 = new_n2591 & new_n6214 ;
  assign new_n6216 = lo0600 & new_n2601 ;
  assign new_n6217 = lo0601 & new_n2605 ;
  assign new_n6218 = ~new_n6216 & ~new_n6217 ;
  assign new_n6219 = lo1334 & new_n2610 ;
  assign new_n6220 = lo0602 & new_n2613 ;
  assign new_n6221 = ~new_n6219 & ~new_n6220 ;
  assign new_n6222 = new_n6218 & new_n6221 ;
  assign new_n6223 = ~new_n6215 & new_n6222 ;
  assign new_n6224 = ~new_n6203 & new_n6223 ;
  assign new_n6225 = ~new_n6186 & new_n6224 ;
  assign new_n6226 = new_n3737 & ~new_n4630 ;
  assign new_n6227 = new_n3820 & ~new_n4268 ;
  assign new_n6228 = ~new_n3819 & ~new_n6227 ;
  assign new_n6229 = ~new_n6226 & new_n6228 ;
  assign new_n6230 = ~new_n3735 & ~new_n6229 ;
  assign new_n6231 = new_n3735 & new_n6229 ;
  assign new_n6232 = ~new_n6230 & ~new_n6231 ;
  assign new_n6233 = ~new_n6225 & ~new_n6232 ;
  assign new_n6234 = new_n6225 & new_n6230 ;
  assign new_n6235 = ~new_n3734 & new_n3735 ;
  assign new_n6236 = ~new_n6229 & new_n6235 ;
  assign new_n6237 = ~new_n6234 & ~new_n6236 ;
  assign new_n6238 = ~new_n6233 & new_n6237 ;
  assign new_n6239 = new_n5673 & new_n6238 ;
  assign new_n6240 = ~new_n5782 & ~new_n6238 ;
  assign new_n6241 = ~new_n3549 & new_n5784 ;
  assign new_n6242 = ~new_n6240 & ~new_n6241 ;
  assign new_n6243 = ~new_n6239 & new_n6242 ;
  assign new_n6244 = ~new_n5672 & ~new_n6243 ;
  assign new_n6245 = new_n5672 & new_n6243 ;
  assign new_n6246 = ~new_n6244 & ~new_n6245 ;
  assign new_n6247 = ~new_n2824 & ~new_n6246 ;
  assign new_n6248 = new_n2824 & new_n6244 ;
  assign new_n6249 = ~new_n3001 & new_n5672 ;
  assign new_n6250 = ~new_n6243 & new_n6249 ;
  assign new_n6251 = ~new_n6248 & ~new_n6250 ;
  assign new_n6252 = ~new_n6247 & new_n6251 ;
  assign new_n6253 = new_n3102 & ~new_n6252 ;
  assign new_n6254 = ~new_n3102 & ~new_n3908 ;
  assign new_n6255 = ~new_n6253 & ~new_n6254 ;
  assign new_n6256 = lo0363 & new_n3170 ;
  assign new_n6257 = lo0362 & new_n3173 ;
  assign new_n6258 = ~new_n3172 & ~new_n6257 ;
  assign new_n6259 = ~new_n6256 & new_n6258 ;
  assign new_n6260 = ~lo0059 & ~new_n6259 ;
  assign new_n6261 = lo0059 & new_n6259 ;
  assign new_n6262 = ~new_n6260 & ~new_n6261 ;
  assign new_n6263 = lo0361 & ~new_n6262 ;
  assign new_n6264 = ~lo0361 & new_n6260 ;
  assign new_n6265 = lo0059 & lo0364 ;
  assign new_n6266 = ~new_n6259 & new_n6265 ;
  assign new_n6267 = ~new_n6264 & ~new_n6266 ;
  assign new_n6268 = ~new_n6263 & new_n6267 ;
  assign new_n6269 = lo0371 & new_n3170 ;
  assign new_n6270 = lo0370 & new_n3204 ;
  assign new_n6271 = ~new_n3172 & ~new_n6270 ;
  assign new_n6272 = ~new_n6269 & new_n6271 ;
  assign new_n6273 = ~lo0061 & ~new_n6272 ;
  assign new_n6274 = lo0061 & new_n6272 ;
  assign new_n6275 = ~new_n6273 & ~new_n6274 ;
  assign new_n6276 = lo0369 & ~new_n6275 ;
  assign new_n6277 = ~lo0369 & new_n6273 ;
  assign new_n6278 = lo0061 & lo0372 ;
  assign new_n6279 = ~new_n6272 & new_n6278 ;
  assign new_n6280 = ~new_n6277 & ~new_n6279 ;
  assign new_n6281 = ~new_n6276 & new_n6280 ;
  assign new_n6282 = new_n3186 & ~new_n6281 ;
  assign new_n6283 = lo0367 & new_n3170 ;
  assign new_n6284 = lo0366 & new_n3204 ;
  assign new_n6285 = ~new_n3172 & ~new_n6284 ;
  assign new_n6286 = ~new_n6283 & new_n6285 ;
  assign new_n6287 = ~lo0061 & ~new_n6286 ;
  assign new_n6288 = lo0061 & new_n6286 ;
  assign new_n6289 = ~new_n6287 & ~new_n6288 ;
  assign new_n6290 = lo0365 & ~new_n6289 ;
  assign new_n6291 = ~lo0365 & new_n6287 ;
  assign new_n6292 = lo0061 & lo0368 ;
  assign new_n6293 = ~new_n6286 & new_n6292 ;
  assign new_n6294 = ~new_n6291 & ~new_n6293 ;
  assign new_n6295 = ~new_n6290 & new_n6294 ;
  assign new_n6296 = new_n3559 & ~new_n6295 ;
  assign new_n6297 = ~new_n3201 & ~new_n6296 ;
  assign new_n6298 = ~new_n6282 & new_n6297 ;
  assign new_n6299 = ~lo0065 & ~new_n6298 ;
  assign new_n6300 = lo0065 & new_n6298 ;
  assign new_n6301 = ~new_n6299 & ~new_n6300 ;
  assign new_n6302 = ~new_n6268 & ~new_n6301 ;
  assign new_n6303 = new_n6268 & new_n6299 ;
  assign new_n6304 = lo0375 & new_n3170 ;
  assign new_n6305 = lo0374 & new_n3173 ;
  assign new_n6306 = ~new_n3172 & ~new_n6305 ;
  assign new_n6307 = ~new_n6304 & new_n6306 ;
  assign new_n6308 = ~lo0059 & ~new_n6307 ;
  assign new_n6309 = lo0059 & new_n6307 ;
  assign new_n6310 = ~new_n6308 & ~new_n6309 ;
  assign new_n6311 = lo0373 & ~new_n6310 ;
  assign new_n6312 = ~lo0373 & new_n6308 ;
  assign new_n6313 = lo0059 & lo0376 ;
  assign new_n6314 = ~new_n6307 & new_n6313 ;
  assign new_n6315 = ~new_n6312 & ~new_n6314 ;
  assign new_n6316 = ~new_n6311 & new_n6315 ;
  assign new_n6317 = lo0065 & ~new_n6316 ;
  assign new_n6318 = ~new_n6298 & new_n6317 ;
  assign new_n6319 = ~new_n6303 & ~new_n6318 ;
  assign new_n6320 = ~new_n6302 & new_n6319 ;
  assign new_n6321 = new_n3169 & ~new_n6320 ;
  assign new_n6322 = ~new_n3160 & new_n3897 ;
  assign new_n6323 = lo1342 & new_n3246 ;
  assign new_n6324 = lo1308 & new_n3254 ;
  assign new_n6325 = lo0379 & new_n3258 ;
  assign new_n6326 = ~new_n6324 & ~new_n6325 ;
  assign new_n6327 = ~new_n6323 & new_n6326 ;
  assign new_n6328 = lo1341 & new_n3267 ;
  assign new_n6329 = lo1343 & new_n3270 ;
  assign new_n6330 = lo0378 & new_n3274 ;
  assign new_n6331 = ~new_n6329 & ~new_n6330 ;
  assign new_n6332 = ~new_n6328 & new_n6331 ;
  assign new_n6333 = ~new_n3265 & new_n6332 ;
  assign new_n6334 = new_n6327 & new_n6333 ;
  assign new_n6335 = ~new_n6322 & new_n6334 ;
  assign new_n6336 = ~new_n6321 & new_n6335 ;
  assign new_n6337 = new_n3141 & ~new_n6336 ;
  assign new_n6338 = new_n3140 & ~new_n6337 ;
  assign new_n6339 = ~new_n3121 & ~new_n6338 ;
  assign new_n6340 = new_n3121 & new_n6338 ;
  assign new_n6341 = ~new_n6339 & ~new_n6340 ;
  assign new_n6342 = lo0371 & ~new_n6341 ;
  assign new_n6343 = ~lo0371 & new_n6339 ;
  assign new_n6344 = new_n3121 & new_n3897 ;
  assign new_n6345 = ~new_n6338 & new_n6344 ;
  assign new_n6346 = ~new_n6343 & ~new_n6345 ;
  assign new_n6347 = ~new_n6342 & new_n6346 ;
  assign new_n6348 = ~new_n3112 & new_n6347 ;
  assign new_n6349 = new_n3112 & ~new_n6347 ;
  assign new_n6350 = ~new_n6348 & ~new_n6349 ;
  assign new_n6351 = new_n3737 & ~new_n4992 ;
  assign new_n6352 = lo0204 & new_n2490 ;
  assign new_n6353 = lo0203 & new_n2493 ;
  assign new_n6354 = ~new_n2492 & ~new_n6353 ;
  assign new_n6355 = ~new_n6352 & new_n6354 ;
  assign new_n6356 = ~lo0249 & ~new_n6355 ;
  assign new_n6357 = lo0249 & new_n6355 ;
  assign new_n6358 = ~new_n6356 & ~new_n6357 ;
  assign new_n6359 = lo0202 & ~new_n6358 ;
  assign new_n6360 = ~lo0202 & new_n6356 ;
  assign new_n6361 = lo0205 & lo0249 ;
  assign new_n6362 = ~new_n6355 & new_n6361 ;
  assign new_n6363 = ~new_n6360 & ~new_n6362 ;
  assign new_n6364 = ~new_n6359 & new_n6363 ;
  assign new_n6365 = lo0201 & new_n2490 ;
  assign new_n6366 = lo0211 & new_n2493 ;
  assign new_n6367 = ~new_n2492 & ~new_n6366 ;
  assign new_n6368 = ~new_n6365 & new_n6367 ;
  assign new_n6369 = ~lo0249 & ~new_n6368 ;
  assign new_n6370 = lo0249 & new_n6368 ;
  assign new_n6371 = ~new_n6369 & ~new_n6370 ;
  assign new_n6372 = lo0210 & ~new_n6371 ;
  assign new_n6373 = ~lo0210 & new_n6369 ;
  assign new_n6374 = lo0212 & lo0249 ;
  assign new_n6375 = ~new_n6368 & new_n6374 ;
  assign new_n6376 = ~new_n6373 & ~new_n6375 ;
  assign new_n6377 = ~new_n6372 & new_n6376 ;
  assign new_n6378 = new_n2506 & ~new_n6377 ;
  assign new_n6379 = lo0208 & new_n2490 ;
  assign new_n6380 = lo0207 & new_n3310 ;
  assign new_n6381 = ~new_n2492 & ~new_n6380 ;
  assign new_n6382 = ~new_n6379 & new_n6381 ;
  assign new_n6383 = ~lo0250 & ~new_n6382 ;
  assign new_n6384 = lo0250 & new_n6382 ;
  assign new_n6385 = ~new_n6383 & ~new_n6384 ;
  assign new_n6386 = lo0206 & ~new_n6385 ;
  assign new_n6387 = ~lo0206 & new_n6383 ;
  assign new_n6388 = lo0209 & lo0250 ;
  assign new_n6389 = ~new_n6382 & new_n6388 ;
  assign new_n6390 = ~new_n6387 & ~new_n6389 ;
  assign new_n6391 = ~new_n6386 & new_n6390 ;
  assign new_n6392 = new_n2522 & ~new_n6391 ;
  assign new_n6393 = ~new_n2521 & ~new_n6392 ;
  assign new_n6394 = ~new_n6378 & new_n6393 ;
  assign new_n6395 = ~lo0251 & ~new_n6394 ;
  assign new_n6396 = lo0251 & new_n6394 ;
  assign new_n6397 = ~new_n6395 & ~new_n6396 ;
  assign new_n6398 = ~new_n6364 & ~new_n6397 ;
  assign new_n6399 = new_n6364 & new_n6395 ;
  assign new_n6400 = lo0215 & new_n2490 ;
  assign new_n6401 = lo0214 & new_n3310 ;
  assign new_n6402 = ~new_n2492 & ~new_n6401 ;
  assign new_n6403 = ~new_n6400 & new_n6402 ;
  assign new_n6404 = ~lo0250 & ~new_n6403 ;
  assign new_n6405 = lo0250 & new_n6403 ;
  assign new_n6406 = ~new_n6404 & ~new_n6405 ;
  assign new_n6407 = lo0213 & ~new_n6406 ;
  assign new_n6408 = ~lo0213 & new_n6404 ;
  assign new_n6409 = lo0216 & lo0250 ;
  assign new_n6410 = ~new_n6403 & new_n6409 ;
  assign new_n6411 = ~new_n6408 & ~new_n6410 ;
  assign new_n6412 = ~new_n6407 & new_n6411 ;
  assign new_n6413 = lo0251 & ~new_n6412 ;
  assign new_n6414 = ~new_n6394 & new_n6413 ;
  assign new_n6415 = ~new_n6399 & ~new_n6414 ;
  assign new_n6416 = ~new_n6398 & new_n6415 ;
  assign new_n6417 = new_n2489 & ~new_n6416 ;
  assign new_n6418 = lo0219 & new_n2565 ;
  assign new_n6419 = new_n2569 & new_n6418 ;
  assign new_n6420 = lo0218 & ~new_n2565 ;
  assign new_n6421 = new_n2569 & new_n6420 ;
  assign new_n6422 = ~new_n2572 & ~new_n6421 ;
  assign new_n6423 = ~new_n6419 & new_n6422 ;
  assign new_n6424 = new_n2569 & ~new_n6423 ;
  assign new_n6425 = ~new_n2569 & new_n6423 ;
  assign new_n6426 = ~new_n6424 & ~new_n6425 ;
  assign new_n6427 = lo0217 & ~new_n6426 ;
  assign new_n6428 = ~lo0217 & new_n6424 ;
  assign new_n6429 = lo0220 & ~new_n2569 ;
  assign new_n6430 = ~new_n6423 & new_n6429 ;
  assign new_n6431 = ~new_n6428 & ~new_n6430 ;
  assign new_n6432 = ~new_n6427 & new_n6431 ;
  assign new_n6433 = lo0090 & ~new_n6432 ;
  assign new_n6434 = ~new_n2483 & new_n6433 ;
  assign new_n6435 = lo0224 & new_n2594 ;
  assign new_n6436 = lo0221 & ~new_n5746 ;
  assign new_n6437 = lo0223 & new_n5461 ;
  assign new_n6438 = ~new_n6436 & ~new_n6437 ;
  assign new_n6439 = ~new_n6435 & new_n6438 ;
  assign new_n6440 = ~lo0105 & new_n2592 ;
  assign new_n6441 = ~new_n6439 & new_n6440 ;
  assign new_n6442 = ~lo0107 & lo0223 ;
  assign new_n6443 = lo0108 & new_n6442 ;
  assign new_n6444 = lo0105 & lo0224 ;
  assign new_n6445 = new_n2592 & new_n6444 ;
  assign new_n6446 = lo0107 & lo0221 ;
  assign new_n6447 = ~new_n6445 & ~new_n6446 ;
  assign new_n6448 = ~new_n6443 & new_n6447 ;
  assign new_n6449 = ~new_n6441 & new_n6448 ;
  assign new_n6450 = ~lo0106 & ~new_n6449 ;
  assign new_n6451 = new_n2591 & new_n6450 ;
  assign new_n6452 = lo0226 & new_n2601 ;
  assign new_n6453 = lo0321 & new_n2605 ;
  assign new_n6454 = ~new_n6452 & ~new_n6453 ;
  assign new_n6455 = lo1295 & new_n2610 ;
  assign new_n6456 = lo0225 & new_n2613 ;
  assign new_n6457 = ~new_n6455 & ~new_n6456 ;
  assign new_n6458 = new_n6454 & new_n6457 ;
  assign new_n6459 = ~new_n6451 & new_n6458 ;
  assign new_n6460 = ~new_n6434 & new_n6459 ;
  assign new_n6461 = ~new_n6417 & new_n6460 ;
  assign new_n6462 = new_n4180 & ~new_n6461 ;
  assign new_n6463 = ~new_n3819 & ~new_n6462 ;
  assign new_n6464 = ~new_n6351 & new_n6463 ;
  assign new_n6465 = new_n3736 & ~new_n6464 ;
  assign new_n6466 = ~new_n3736 & new_n6464 ;
  assign new_n6467 = ~new_n6465 & ~new_n6466 ;
  assign new_n6468 = ~new_n4630 & ~new_n6467 ;
  assign new_n6469 = new_n4630 & new_n6465 ;
  assign new_n6470 = ~new_n3736 & ~new_n4179 ;
  assign new_n6471 = ~new_n6464 & new_n6470 ;
  assign new_n6472 = ~new_n6469 & ~new_n6471 ;
  assign new_n6473 = ~new_n6468 & new_n6472 ;
  assign new_n6474 = new_n5673 & new_n6473 ;
  assign new_n6475 = ~new_n5782 & ~new_n6473 ;
  assign new_n6476 = ~new_n3908 & new_n5784 ;
  assign new_n6477 = ~new_n6475 & ~new_n6476 ;
  assign new_n6478 = ~new_n6474 & new_n6477 ;
  assign new_n6479 = ~new_n5672 & ~new_n6478 ;
  assign new_n6480 = new_n5672 & new_n6478 ;
  assign new_n6481 = ~new_n6479 & ~new_n6480 ;
  assign new_n6482 = ~new_n3549 & ~new_n6481 ;
  assign new_n6483 = new_n3549 & new_n6479 ;
  assign new_n6484 = ~new_n3464 & new_n5672 ;
  assign new_n6485 = ~new_n6478 & new_n6484 ;
  assign new_n6486 = ~new_n6483 & ~new_n6485 ;
  assign new_n6487 = ~new_n6482 & new_n6486 ;
  assign new_n6488 = new_n3102 & ~new_n6487 ;
  assign new_n6489 = ~new_n3102 & ~new_n4268 ;
  assign new_n6490 = ~new_n6488 & ~new_n6489 ;
  assign new_n6491 = lo0232 & new_n3186 ;
  assign new_n6492 = lo0231 & new_n3559 ;
  assign new_n6493 = ~new_n3201 & ~new_n6492 ;
  assign new_n6494 = ~new_n6491 & new_n6493 ;
  assign new_n6495 = ~lo0065 & ~new_n6494 ;
  assign new_n6496 = lo0065 & new_n6494 ;
  assign new_n6497 = ~new_n6495 & ~new_n6496 ;
  assign new_n6498 = lo0230 & ~new_n6497 ;
  assign new_n6499 = ~lo0230 & new_n6495 ;
  assign new_n6500 = lo0065 & lo0233 ;
  assign new_n6501 = ~new_n6494 & new_n6500 ;
  assign new_n6502 = ~new_n6499 & ~new_n6501 ;
  assign new_n6503 = ~new_n6498 & new_n6502 ;
  assign new_n6504 = lo0227 & new_n3186 ;
  assign new_n6505 = lo0239 & new_n3202 ;
  assign new_n6506 = ~new_n3201 & ~new_n6505 ;
  assign new_n6507 = ~new_n6504 & new_n6506 ;
  assign new_n6508 = ~lo0063 & ~new_n6507 ;
  assign new_n6509 = lo0063 & new_n6507 ;
  assign new_n6510 = ~new_n6508 & ~new_n6509 ;
  assign new_n6511 = lo0238 & ~new_n6510 ;
  assign new_n6512 = ~lo0238 & new_n6508 ;
  assign new_n6513 = lo0063 & lo0240 ;
  assign new_n6514 = ~new_n6507 & new_n6513 ;
  assign new_n6515 = ~new_n6512 & ~new_n6514 ;
  assign new_n6516 = ~new_n6511 & new_n6515 ;
  assign new_n6517 = new_n3170 & ~new_n6516 ;
  assign new_n6518 = lo0236 & new_n3186 ;
  assign new_n6519 = lo0235 & new_n3202 ;
  assign new_n6520 = ~new_n3201 & ~new_n6519 ;
  assign new_n6521 = ~new_n6518 & new_n6520 ;
  assign new_n6522 = ~lo0063 & ~new_n6521 ;
  assign new_n6523 = lo0063 & new_n6521 ;
  assign new_n6524 = ~new_n6522 & ~new_n6523 ;
  assign new_n6525 = lo0234 & ~new_n6524 ;
  assign new_n6526 = ~lo0234 & new_n6522 ;
  assign new_n6527 = lo0063 & lo0237 ;
  assign new_n6528 = ~new_n6521 & new_n6527 ;
  assign new_n6529 = ~new_n6526 & ~new_n6528 ;
  assign new_n6530 = ~new_n6525 & new_n6529 ;
  assign new_n6531 = new_n3204 & ~new_n6530 ;
  assign new_n6532 = ~new_n3172 & ~new_n6531 ;
  assign new_n6533 = ~new_n6517 & new_n6532 ;
  assign new_n6534 = ~lo0061 & ~new_n6533 ;
  assign new_n6535 = lo0061 & new_n6533 ;
  assign new_n6536 = ~new_n6534 & ~new_n6535 ;
  assign new_n6537 = ~new_n6503 & ~new_n6536 ;
  assign new_n6538 = new_n6503 & new_n6534 ;
  assign new_n6539 = lo0243 & new_n3186 ;
  assign new_n6540 = lo0242 & new_n3559 ;
  assign new_n6541 = ~new_n3201 & ~new_n6540 ;
  assign new_n6542 = ~new_n6539 & new_n6541 ;
  assign new_n6543 = ~lo0065 & ~new_n6542 ;
  assign new_n6544 = lo0065 & new_n6542 ;
  assign new_n6545 = ~new_n6543 & ~new_n6544 ;
  assign new_n6546 = lo0241 & ~new_n6545 ;
  assign new_n6547 = ~lo0241 & new_n6543 ;
  assign new_n6548 = lo0065 & lo0244 ;
  assign new_n6549 = ~new_n6542 & new_n6548 ;
  assign new_n6550 = ~new_n6547 & ~new_n6549 ;
  assign new_n6551 = ~new_n6546 & new_n6550 ;
  assign new_n6552 = lo0061 & ~new_n6551 ;
  assign new_n6553 = ~new_n6533 & new_n6552 ;
  assign new_n6554 = ~new_n6538 & ~new_n6553 ;
  assign new_n6555 = ~new_n6537 & new_n6554 ;
  assign new_n6556 = new_n3169 & ~new_n6555 ;
  assign new_n6557 = ~new_n3160 & new_n4257 ;
  assign new_n6558 = lo1299 & new_n3267 ;
  assign new_n6559 = lo1301 & new_n3246 ;
  assign new_n6560 = lo0246 & new_n3258 ;
  assign new_n6561 = ~new_n6559 & ~new_n6560 ;
  assign new_n6562 = ~new_n6558 & new_n6561 ;
  assign new_n6563 = lo1300 & new_n3254 ;
  assign new_n6564 = lo1302 & new_n3270 ;
  assign new_n6565 = lo0245 & new_n3274 ;
  assign new_n6566 = ~new_n6564 & ~new_n6565 ;
  assign new_n6567 = ~new_n6563 & new_n6566 ;
  assign new_n6568 = ~new_n3265 & new_n6567 ;
  assign new_n6569 = new_n6562 & new_n6568 ;
  assign new_n6570 = ~new_n6557 & new_n6569 ;
  assign new_n6571 = ~new_n6556 & new_n6570 ;
  assign new_n6572 = new_n3141 & ~new_n6571 ;
  assign new_n6573 = new_n3140 & ~new_n6572 ;
  assign new_n6574 = ~new_n3121 & ~new_n6573 ;
  assign new_n6575 = new_n3121 & new_n6573 ;
  assign new_n6576 = ~new_n6574 & ~new_n6575 ;
  assign new_n6577 = lo0227 & ~new_n6576 ;
  assign new_n6578 = ~lo0227 & new_n6574 ;
  assign new_n6579 = new_n3121 & new_n4257 ;
  assign new_n6580 = ~new_n6573 & new_n6579 ;
  assign new_n6581 = ~new_n6578 & ~new_n6580 ;
  assign new_n6582 = ~new_n6577 & new_n6581 ;
  assign new_n6583 = ~new_n3112 & new_n6582 ;
  assign new_n6584 = new_n3112 & ~new_n6582 ;
  assign new_n6585 = ~new_n6583 & ~new_n6584 ;
  assign new_n6586 = lo0562 & new_n2506 ;
  assign new_n6587 = lo0561 & new_n2831 ;
  assign new_n6588 = ~new_n2521 & ~new_n6587 ;
  assign new_n6589 = ~new_n6586 & new_n6588 ;
  assign new_n6590 = ~lo0252 & ~new_n6589 ;
  assign new_n6591 = lo0252 & new_n6589 ;
  assign new_n6592 = ~new_n6590 & ~new_n6591 ;
  assign new_n6593 = lo0560 & ~new_n6592 ;
  assign new_n6594 = ~lo0560 & new_n6590 ;
  assign new_n6595 = lo0252 & lo0563 ;
  assign new_n6596 = ~new_n6589 & new_n6595 ;
  assign new_n6597 = ~new_n6594 & ~new_n6596 ;
  assign new_n6598 = ~new_n6593 & new_n6597 ;
  assign new_n6599 = lo0570 & new_n2506 ;
  assign new_n6600 = lo0569 & new_n2831 ;
  assign new_n6601 = ~new_n2521 & ~new_n6600 ;
  assign new_n6602 = ~new_n6599 & new_n6601 ;
  assign new_n6603 = ~lo0252 & ~new_n6602 ;
  assign new_n6604 = lo0252 & new_n6602 ;
  assign new_n6605 = ~new_n6603 & ~new_n6604 ;
  assign new_n6606 = lo0568 & ~new_n6605 ;
  assign new_n6607 = ~lo0568 & new_n6603 ;
  assign new_n6608 = lo0252 & lo0571 ;
  assign new_n6609 = ~new_n6602 & new_n6608 ;
  assign new_n6610 = ~new_n6607 & ~new_n6609 ;
  assign new_n6611 = ~new_n6606 & new_n6610 ;
  assign new_n6612 = new_n2490 & ~new_n6611 ;
  assign new_n6613 = lo0566 & new_n2506 ;
  assign new_n6614 = lo0565 & new_n2522 ;
  assign new_n6615 = ~new_n2521 & ~new_n6614 ;
  assign new_n6616 = ~new_n6613 & new_n6615 ;
  assign new_n6617 = ~lo0251 & ~new_n6616 ;
  assign new_n6618 = lo0251 & new_n6616 ;
  assign new_n6619 = ~new_n6617 & ~new_n6618 ;
  assign new_n6620 = lo0564 & ~new_n6619 ;
  assign new_n6621 = ~lo0564 & new_n6617 ;
  assign new_n6622 = lo0251 & lo0567 ;
  assign new_n6623 = ~new_n6616 & new_n6622 ;
  assign new_n6624 = ~new_n6621 & ~new_n6623 ;
  assign new_n6625 = ~new_n6620 & new_n6624 ;
  assign new_n6626 = new_n2493 & ~new_n6625 ;
  assign new_n6627 = ~new_n2492 & ~new_n6626 ;
  assign new_n6628 = ~new_n6612 & new_n6627 ;
  assign new_n6629 = ~lo0249 & ~new_n6628 ;
  assign new_n6630 = lo0249 & new_n6628 ;
  assign new_n6631 = ~new_n6629 & ~new_n6630 ;
  assign new_n6632 = ~new_n6598 & ~new_n6631 ;
  assign new_n6633 = new_n6598 & new_n6629 ;
  assign new_n6634 = lo0574 & new_n2506 ;
  assign new_n6635 = lo0573 & new_n2522 ;
  assign new_n6636 = ~new_n2521 & ~new_n6635 ;
  assign new_n6637 = ~new_n6634 & new_n6636 ;
  assign new_n6638 = ~lo0251 & ~new_n6637 ;
  assign new_n6639 = lo0251 & new_n6637 ;
  assign new_n6640 = ~new_n6638 & ~new_n6639 ;
  assign new_n6641 = lo0572 & ~new_n6640 ;
  assign new_n6642 = ~lo0572 & new_n6638 ;
  assign new_n6643 = lo0251 & lo0575 ;
  assign new_n6644 = ~new_n6637 & new_n6643 ;
  assign new_n6645 = ~new_n6642 & ~new_n6644 ;
  assign new_n6646 = ~new_n6641 & new_n6645 ;
  assign new_n6647 = lo0249 & ~new_n6646 ;
  assign new_n6648 = ~new_n6628 & new_n6647 ;
  assign new_n6649 = ~new_n6633 & ~new_n6648 ;
  assign new_n6650 = ~new_n6632 & new_n6649 ;
  assign new_n6651 = new_n2489 & ~new_n6650 ;
  assign new_n6652 = lo0577 & new_n2565 ;
  assign new_n6653 = new_n2569 & new_n6652 ;
  assign new_n6654 = lo0576 & new_n2565 ;
  assign new_n6655 = ~new_n2569 & new_n6654 ;
  assign new_n6656 = ~new_n2572 & ~new_n6655 ;
  assign new_n6657 = ~new_n6653 & new_n6656 ;
  assign new_n6658 = new_n2565 & ~new_n6657 ;
  assign new_n6659 = ~new_n2565 & new_n6657 ;
  assign new_n6660 = ~new_n6658 & ~new_n6659 ;
  assign new_n6661 = lo0317 & ~new_n6660 ;
  assign new_n6662 = ~lo0317 & new_n6658 ;
  assign new_n6663 = lo0578 & ~new_n2565 ;
  assign new_n6664 = ~new_n6657 & new_n6663 ;
  assign new_n6665 = ~new_n6662 & ~new_n6664 ;
  assign new_n6666 = ~new_n6661 & new_n6665 ;
  assign new_n6667 = lo0090 & ~new_n6666 ;
  assign new_n6668 = ~new_n2483 & new_n6667 ;
  assign new_n6669 = new_n2592 & ~new_n5748 ;
  assign new_n6670 = ~lo0106 & ~new_n6669 ;
  assign new_n6671 = lo0221 & ~new_n6670 ;
  assign new_n6672 = ~lo0105 & ~lo0108 ;
  assign new_n6673 = ~new_n5746 & new_n6672 ;
  assign new_n6674 = ~lo0107 & ~new_n6673 ;
  assign new_n6675 = lo0223 & ~new_n6674 ;
  assign new_n6676 = lo0579 & new_n6674 ;
  assign new_n6677 = ~new_n6675 & ~new_n6676 ;
  assign new_n6678 = new_n6670 & ~new_n6677 ;
  assign new_n6679 = ~new_n6671 & ~new_n6678 ;
  assign new_n6680 = new_n2591 & ~new_n6679 ;
  assign new_n6681 = lo0580 & new_n2601 ;
  assign new_n6682 = lo0581 & new_n2605 ;
  assign new_n6683 = ~new_n6681 & ~new_n6682 ;
  assign new_n6684 = lo1333 & new_n2610 ;
  assign new_n6685 = lo0582 & new_n2613 ;
  assign new_n6686 = ~new_n6684 & ~new_n6685 ;
  assign new_n6687 = new_n6683 & new_n6686 ;
  assign new_n6688 = ~new_n6680 & new_n6687 ;
  assign new_n6689 = ~new_n6668 & new_n6688 ;
  assign new_n6690 = ~new_n6651 & new_n6689 ;
  assign new_n6691 = new_n3737 & ~new_n5276 ;
  assign new_n6692 = ~new_n3819 & ~new_n6691 ;
  assign new_n6693 = new_n3820 & ~new_n4992 ;
  assign new_n6694 = new_n6692 & ~new_n6693 ;
  assign new_n6695 = ~new_n3735 & ~new_n6694 ;
  assign new_n6696 = new_n3735 & new_n6694 ;
  assign new_n6697 = ~new_n6695 & ~new_n6696 ;
  assign new_n6698 = ~new_n6690 & ~new_n6697 ;
  assign new_n6699 = new_n6690 & new_n6695 ;
  assign new_n6700 = new_n3735 & ~new_n4461 ;
  assign new_n6701 = ~new_n6694 & new_n6700 ;
  assign new_n6702 = ~new_n6699 & ~new_n6701 ;
  assign new_n6703 = ~new_n6698 & new_n6702 ;
  assign new_n6704 = new_n5673 & new_n6703 ;
  assign new_n6705 = ~new_n5782 & ~new_n6703 ;
  assign new_n6706 = ~new_n4268 & new_n5784 ;
  assign new_n6707 = ~new_n6705 & ~new_n6706 ;
  assign new_n6708 = ~new_n6704 & new_n6707 ;
  assign new_n6709 = ~new_n5672 & ~new_n6708 ;
  assign new_n6710 = new_n5672 & new_n6708 ;
  assign new_n6711 = ~new_n6709 & ~new_n6710 ;
  assign new_n6712 = ~new_n3908 & ~new_n6711 ;
  assign new_n6713 = new_n3908 & new_n6709 ;
  assign new_n6714 = ~new_n3817 & new_n5672 ;
  assign new_n6715 = ~new_n6708 & new_n6714 ;
  assign new_n6716 = ~new_n6713 & ~new_n6715 ;
  assign new_n6717 = ~new_n6712 & new_n6716 ;
  assign new_n6718 = new_n3102 & ~new_n6717 ;
  assign new_n6719 = ~new_n3102 & ~new_n4630 ;
  assign new_n6720 = ~new_n6718 & ~new_n6719 ;
  assign new_n6721 = lo0303 & new_n3170 ;
  assign new_n6722 = lo0302 & new_n3173 ;
  assign new_n6723 = ~new_n3172 & ~new_n6722 ;
  assign new_n6724 = ~new_n6721 & new_n6723 ;
  assign new_n6725 = ~lo0059 & ~new_n6724 ;
  assign new_n6726 = lo0059 & new_n6724 ;
  assign new_n6727 = ~new_n6725 & ~new_n6726 ;
  assign new_n6728 = lo0301 & ~new_n6727 ;
  assign new_n6729 = ~lo0301 & new_n6725 ;
  assign new_n6730 = lo0059 & lo0304 ;
  assign new_n6731 = ~new_n6724 & new_n6730 ;
  assign new_n6732 = ~new_n6729 & ~new_n6731 ;
  assign new_n6733 = ~new_n6728 & new_n6732 ;
  assign new_n6734 = lo0311 & new_n3170 ;
  assign new_n6735 = lo0310 & new_n3173 ;
  assign new_n6736 = ~new_n3172 & ~new_n6735 ;
  assign new_n6737 = ~new_n6734 & new_n6736 ;
  assign new_n6738 = ~lo0059 & ~new_n6737 ;
  assign new_n6739 = lo0059 & new_n6737 ;
  assign new_n6740 = ~new_n6738 & ~new_n6739 ;
  assign new_n6741 = lo0309 & ~new_n6740 ;
  assign new_n6742 = ~lo0309 & new_n6738 ;
  assign new_n6743 = lo0059 & lo0312 ;
  assign new_n6744 = ~new_n6737 & new_n6743 ;
  assign new_n6745 = ~new_n6742 & ~new_n6744 ;
  assign new_n6746 = ~new_n6741 & new_n6745 ;
  assign new_n6747 = new_n3186 & ~new_n6746 ;
  assign new_n6748 = lo0307 & new_n3170 ;
  assign new_n6749 = lo0306 & new_n3204 ;
  assign new_n6750 = ~new_n3172 & ~new_n6749 ;
  assign new_n6751 = ~new_n6748 & new_n6750 ;
  assign new_n6752 = ~lo0061 & ~new_n6751 ;
  assign new_n6753 = lo0061 & new_n6751 ;
  assign new_n6754 = ~new_n6752 & ~new_n6753 ;
  assign new_n6755 = lo0305 & ~new_n6754 ;
  assign new_n6756 = ~lo0305 & new_n6752 ;
  assign new_n6757 = lo0061 & lo0308 ;
  assign new_n6758 = ~new_n6751 & new_n6757 ;
  assign new_n6759 = ~new_n6756 & ~new_n6758 ;
  assign new_n6760 = ~new_n6755 & new_n6759 ;
  assign new_n6761 = new_n3202 & ~new_n6760 ;
  assign new_n6762 = ~new_n3201 & ~new_n6761 ;
  assign new_n6763 = ~new_n6747 & new_n6762 ;
  assign new_n6764 = ~lo0063 & ~new_n6763 ;
  assign new_n6765 = lo0063 & new_n6763 ;
  assign new_n6766 = ~new_n6764 & ~new_n6765 ;
  assign new_n6767 = ~new_n6733 & ~new_n6766 ;
  assign new_n6768 = new_n6733 & new_n6764 ;
  assign new_n6769 = lo0315 & new_n3170 ;
  assign new_n6770 = lo0314 & new_n3204 ;
  assign new_n6771 = ~new_n3172 & ~new_n6770 ;
  assign new_n6772 = ~new_n6769 & new_n6771 ;
  assign new_n6773 = ~lo0061 & ~new_n6772 ;
  assign new_n6774 = lo0061 & new_n6772 ;
  assign new_n6775 = ~new_n6773 & ~new_n6774 ;
  assign new_n6776 = lo0313 & ~new_n6775 ;
  assign new_n6777 = ~lo0313 & new_n6773 ;
  assign new_n6778 = lo0061 & lo0316 ;
  assign new_n6779 = ~new_n6772 & new_n6778 ;
  assign new_n6780 = ~new_n6777 & ~new_n6779 ;
  assign new_n6781 = ~new_n6776 & new_n6780 ;
  assign new_n6782 = lo0063 & ~new_n6781 ;
  assign new_n6783 = ~new_n6763 & new_n6782 ;
  assign new_n6784 = ~new_n6768 & ~new_n6783 ;
  assign new_n6785 = ~new_n6767 & new_n6784 ;
  assign new_n6786 = new_n3169 & ~new_n6785 ;
  assign new_n6787 = ~new_n3160 & new_n4619 ;
  assign new_n6788 = lo1378 & new_n3246 ;
  assign new_n6789 = lo1305 & new_n3254 ;
  assign new_n6790 = lo0319 & new_n3258 ;
  assign new_n6791 = ~new_n6789 & ~new_n6790 ;
  assign new_n6792 = ~new_n6788 & new_n6791 ;
  assign new_n6793 = lo1377 & new_n3267 ;
  assign new_n6794 = lo1379 & new_n3270 ;
  assign new_n6795 = lo0318 & new_n3274 ;
  assign new_n6796 = ~new_n6794 & ~new_n6795 ;
  assign new_n6797 = ~new_n6793 & new_n6796 ;
  assign new_n6798 = ~new_n3265 & new_n6797 ;
  assign new_n6799 = new_n6792 & new_n6798 ;
  assign new_n6800 = ~new_n6787 & new_n6799 ;
  assign new_n6801 = ~new_n6786 & new_n6800 ;
  assign new_n6802 = new_n3141 & ~new_n6801 ;
  assign new_n6803 = new_n3140 & ~new_n6802 ;
  assign new_n6804 = ~new_n3121 & ~new_n6803 ;
  assign new_n6805 = new_n3121 & new_n6803 ;
  assign new_n6806 = ~new_n6804 & ~new_n6805 ;
  assign new_n6807 = lo0311 & ~new_n6806 ;
  assign new_n6808 = ~lo0311 & new_n6804 ;
  assign new_n6809 = new_n3121 & new_n4619 ;
  assign new_n6810 = ~new_n6803 & new_n6809 ;
  assign new_n6811 = ~new_n6808 & ~new_n6810 ;
  assign new_n6812 = ~new_n6807 & new_n6811 ;
  assign new_n6813 = ~new_n3112 & new_n6812 ;
  assign new_n6814 = new_n3112 & ~new_n6812 ;
  assign new_n6815 = ~new_n6813 & ~new_n6814 ;
  assign new_n6816 = new_n3737 & ~new_n5560 ;
  assign new_n6817 = ~new_n3819 & ~new_n6816 ;
  assign new_n6818 = lo0624 & new_n2490 ;
  assign new_n6819 = lo0623 & new_n2493 ;
  assign new_n6820 = ~new_n2492 & ~new_n6819 ;
  assign new_n6821 = ~new_n6818 & new_n6820 ;
  assign new_n6822 = ~lo0249 & ~new_n6821 ;
  assign new_n6823 = lo0249 & new_n6821 ;
  assign new_n6824 = ~new_n6822 & ~new_n6823 ;
  assign new_n6825 = lo0622 & ~new_n6824 ;
  assign new_n6826 = ~lo0622 & new_n6822 ;
  assign new_n6827 = lo0249 & lo0625 ;
  assign new_n6828 = ~new_n6821 & new_n6827 ;
  assign new_n6829 = ~new_n6826 & ~new_n6828 ;
  assign new_n6830 = ~new_n6825 & new_n6829 ;
  assign new_n6831 = lo0632 & new_n2490 ;
  assign new_n6832 = lo0631 & new_n3310 ;
  assign new_n6833 = ~new_n2492 & ~new_n6832 ;
  assign new_n6834 = ~new_n6831 & new_n6833 ;
  assign new_n6835 = ~lo0250 & ~new_n6834 ;
  assign new_n6836 = lo0250 & new_n6834 ;
  assign new_n6837 = ~new_n6835 & ~new_n6836 ;
  assign new_n6838 = lo0630 & ~new_n6837 ;
  assign new_n6839 = ~lo0630 & new_n6835 ;
  assign new_n6840 = lo0250 & lo0633 ;
  assign new_n6841 = ~new_n6834 & new_n6840 ;
  assign new_n6842 = ~new_n6839 & ~new_n6841 ;
  assign new_n6843 = ~new_n6838 & new_n6842 ;
  assign new_n6844 = new_n2506 & ~new_n6843 ;
  assign new_n6845 = lo0628 & new_n2490 ;
  assign new_n6846 = lo0627 & new_n3310 ;
  assign new_n6847 = ~new_n2492 & ~new_n6846 ;
  assign new_n6848 = ~new_n6845 & new_n6847 ;
  assign new_n6849 = ~lo0250 & ~new_n6848 ;
  assign new_n6850 = lo0250 & new_n6848 ;
  assign new_n6851 = ~new_n6849 & ~new_n6850 ;
  assign new_n6852 = lo0626 & ~new_n6851 ;
  assign new_n6853 = ~lo0626 & new_n6849 ;
  assign new_n6854 = lo0250 & lo0629 ;
  assign new_n6855 = ~new_n6848 & new_n6854 ;
  assign new_n6856 = ~new_n6853 & ~new_n6855 ;
  assign new_n6857 = ~new_n6852 & new_n6856 ;
  assign new_n6858 = new_n2831 & ~new_n6857 ;
  assign new_n6859 = ~new_n2521 & ~new_n6858 ;
  assign new_n6860 = ~new_n6844 & new_n6859 ;
  assign new_n6861 = ~lo0252 & ~new_n6860 ;
  assign new_n6862 = lo0252 & new_n6860 ;
  assign new_n6863 = ~new_n6861 & ~new_n6862 ;
  assign new_n6864 = ~new_n6830 & ~new_n6863 ;
  assign new_n6865 = new_n6830 & new_n6861 ;
  assign new_n6866 = lo0636 & new_n2490 ;
  assign new_n6867 = lo0635 & new_n2493 ;
  assign new_n6868 = ~new_n2492 & ~new_n6867 ;
  assign new_n6869 = ~new_n6866 & new_n6868 ;
  assign new_n6870 = ~lo0249 & ~new_n6869 ;
  assign new_n6871 = lo0249 & new_n6869 ;
  assign new_n6872 = ~new_n6870 & ~new_n6871 ;
  assign new_n6873 = lo0634 & ~new_n6872 ;
  assign new_n6874 = ~lo0634 & new_n6870 ;
  assign new_n6875 = lo0249 & lo0637 ;
  assign new_n6876 = ~new_n6869 & new_n6875 ;
  assign new_n6877 = ~new_n6874 & ~new_n6876 ;
  assign new_n6878 = ~new_n6873 & new_n6877 ;
  assign new_n6879 = lo0252 & ~new_n6878 ;
  assign new_n6880 = ~new_n6860 & new_n6879 ;
  assign new_n6881 = ~new_n6865 & ~new_n6880 ;
  assign new_n6882 = ~new_n6864 & new_n6881 ;
  assign new_n6883 = new_n2489 & ~new_n6882 ;
  assign new_n6884 = lo0639 & new_n2565 ;
  assign new_n6885 = new_n2569 & new_n6884 ;
  assign new_n6886 = lo0338 & ~new_n2565 ;
  assign new_n6887 = new_n2569 & new_n6886 ;
  assign new_n6888 = ~new_n2572 & ~new_n6887 ;
  assign new_n6889 = ~new_n6885 & new_n6888 ;
  assign new_n6890 = new_n2569 & ~new_n6889 ;
  assign new_n6891 = ~new_n2569 & new_n6889 ;
  assign new_n6892 = ~new_n6890 & ~new_n6891 ;
  assign new_n6893 = lo0638 & ~new_n6892 ;
  assign new_n6894 = ~lo0638 & new_n6890 ;
  assign new_n6895 = lo0640 & ~new_n2569 ;
  assign new_n6896 = ~new_n6889 & new_n6895 ;
  assign new_n6897 = ~new_n6894 & ~new_n6896 ;
  assign new_n6898 = ~new_n6893 & new_n6897 ;
  assign new_n6899 = lo0090 & ~new_n6898 ;
  assign new_n6900 = ~new_n2483 & new_n6899 ;
  assign new_n6901 = lo0223 & ~new_n6670 ;
  assign new_n6902 = lo0579 & ~new_n6674 ;
  assign new_n6903 = lo0641 & new_n6674 ;
  assign new_n6904 = ~new_n6902 & ~new_n6903 ;
  assign new_n6905 = new_n6670 & ~new_n6904 ;
  assign new_n6906 = ~new_n6901 & ~new_n6905 ;
  assign new_n6907 = new_n2591 & ~new_n6906 ;
  assign new_n6908 = lo0642 & new_n2601 ;
  assign new_n6909 = lo0643 & new_n2605 ;
  assign new_n6910 = ~new_n6908 & ~new_n6909 ;
  assign new_n6911 = lo1348 & new_n2610 ;
  assign new_n6912 = lo0644 & new_n2613 ;
  assign new_n6913 = ~new_n6911 & ~new_n6912 ;
  assign new_n6914 = new_n6910 & new_n6913 ;
  assign new_n6915 = ~new_n6907 & new_n6914 ;
  assign new_n6916 = ~new_n6900 & new_n6915 ;
  assign new_n6917 = ~new_n6883 & new_n6916 ;
  assign new_n6918 = new_n4180 & ~new_n6917 ;
  assign new_n6919 = new_n6817 & ~new_n6918 ;
  assign new_n6920 = new_n3736 & ~new_n6919 ;
  assign new_n6921 = ~new_n3736 & new_n6919 ;
  assign new_n6922 = ~new_n6920 & ~new_n6921 ;
  assign new_n6923 = ~new_n5276 & ~new_n6922 ;
  assign new_n6924 = new_n5276 & new_n6920 ;
  assign new_n6925 = ~new_n3736 & ~new_n4904 ;
  assign new_n6926 = ~new_n6919 & new_n6925 ;
  assign new_n6927 = ~new_n6924 & ~new_n6926 ;
  assign new_n6928 = ~new_n6923 & new_n6927 ;
  assign new_n6929 = new_n5673 & new_n6928 ;
  assign new_n6930 = ~new_n5782 & ~new_n6928 ;
  assign new_n6931 = ~new_n4630 & new_n5784 ;
  assign new_n6932 = ~new_n6930 & ~new_n6931 ;
  assign new_n6933 = ~new_n6929 & new_n6932 ;
  assign new_n6934 = ~new_n5672 & ~new_n6933 ;
  assign new_n6935 = new_n5672 & new_n6933 ;
  assign new_n6936 = ~new_n6934 & ~new_n6935 ;
  assign new_n6937 = ~new_n4268 & ~new_n6936 ;
  assign new_n6938 = new_n4268 & new_n6934 ;
  assign new_n6939 = ~new_n4097 & new_n5672 ;
  assign new_n6940 = ~new_n6933 & new_n6939 ;
  assign new_n6941 = ~new_n6938 & ~new_n6940 ;
  assign new_n6942 = ~new_n6937 & new_n6941 ;
  assign new_n6943 = new_n3102 & ~new_n6942 ;
  assign new_n6944 = ~new_n3102 & ~new_n4992 ;
  assign new_n6945 = ~new_n6943 & ~new_n6944 ;
  assign new_n6946 = lo0324 & new_n3186 ;
  assign new_n6947 = lo0323 & new_n3559 ;
  assign new_n6948 = ~new_n3201 & ~new_n6947 ;
  assign new_n6949 = ~new_n6946 & new_n6948 ;
  assign new_n6950 = ~lo0065 & ~new_n6949 ;
  assign new_n6951 = lo0065 & new_n6949 ;
  assign new_n6952 = ~new_n6950 & ~new_n6951 ;
  assign new_n6953 = lo0322 & ~new_n6952 ;
  assign new_n6954 = ~lo0322 & new_n6950 ;
  assign new_n6955 = lo0065 & lo0325 ;
  assign new_n6956 = ~new_n6949 & new_n6955 ;
  assign new_n6957 = ~new_n6954 & ~new_n6956 ;
  assign new_n6958 = ~new_n6953 & new_n6957 ;
  assign new_n6959 = lo0332 & new_n3186 ;
  assign new_n6960 = lo0331 & new_n3559 ;
  assign new_n6961 = ~new_n3201 & ~new_n6960 ;
  assign new_n6962 = ~new_n6959 & new_n6961 ;
  assign new_n6963 = ~lo0065 & ~new_n6962 ;
  assign new_n6964 = lo0065 & new_n6962 ;
  assign new_n6965 = ~new_n6963 & ~new_n6964 ;
  assign new_n6966 = lo0330 & ~new_n6965 ;
  assign new_n6967 = ~lo0330 & new_n6963 ;
  assign new_n6968 = lo0065 & lo0333 ;
  assign new_n6969 = ~new_n6962 & new_n6968 ;
  assign new_n6970 = ~new_n6967 & ~new_n6969 ;
  assign new_n6971 = ~new_n6966 & new_n6970 ;
  assign new_n6972 = new_n3170 & ~new_n6971 ;
  assign new_n6973 = lo0328 & new_n3186 ;
  assign new_n6974 = lo0327 & new_n3202 ;
  assign new_n6975 = ~new_n3201 & ~new_n6974 ;
  assign new_n6976 = ~new_n6973 & new_n6975 ;
  assign new_n6977 = ~lo0063 & ~new_n6976 ;
  assign new_n6978 = lo0063 & new_n6976 ;
  assign new_n6979 = ~new_n6977 & ~new_n6978 ;
  assign new_n6980 = lo0326 & ~new_n6979 ;
  assign new_n6981 = ~lo0326 & new_n6977 ;
  assign new_n6982 = lo0063 & lo0329 ;
  assign new_n6983 = ~new_n6976 & new_n6982 ;
  assign new_n6984 = ~new_n6981 & ~new_n6983 ;
  assign new_n6985 = ~new_n6980 & new_n6984 ;
  assign new_n6986 = new_n3173 & ~new_n6985 ;
  assign new_n6987 = ~new_n3172 & ~new_n6986 ;
  assign new_n6988 = ~new_n6972 & new_n6987 ;
  assign new_n6989 = ~lo0059 & ~new_n6988 ;
  assign new_n6990 = lo0059 & new_n6988 ;
  assign new_n6991 = ~new_n6989 & ~new_n6990 ;
  assign new_n6992 = ~new_n6958 & ~new_n6991 ;
  assign new_n6993 = new_n6958 & new_n6989 ;
  assign new_n6994 = lo0336 & new_n3186 ;
  assign new_n6995 = lo0335 & new_n3202 ;
  assign new_n6996 = ~new_n3201 & ~new_n6995 ;
  assign new_n6997 = ~new_n6994 & new_n6996 ;
  assign new_n6998 = ~lo0063 & ~new_n6997 ;
  assign new_n6999 = lo0063 & new_n6997 ;
  assign new_n7000 = ~new_n6998 & ~new_n6999 ;
  assign new_n7001 = lo0334 & ~new_n7000 ;
  assign new_n7002 = ~lo0334 & new_n6998 ;
  assign new_n7003 = lo0063 & lo0337 ;
  assign new_n7004 = ~new_n6997 & new_n7003 ;
  assign new_n7005 = ~new_n7002 & ~new_n7004 ;
  assign new_n7006 = ~new_n7001 & new_n7005 ;
  assign new_n7007 = lo0059 & ~new_n7006 ;
  assign new_n7008 = ~new_n6988 & new_n7007 ;
  assign new_n7009 = ~new_n6993 & ~new_n7008 ;
  assign new_n7010 = ~new_n6992 & new_n7009 ;
  assign new_n7011 = new_n3169 & ~new_n7010 ;
  assign new_n7012 = ~new_n3160 & new_n4981 ;
  assign new_n7013 = lo1372 & new_n3246 ;
  assign new_n7014 = lo1306 & new_n3254 ;
  assign new_n7015 = lo0340 & new_n3258 ;
  assign new_n7016 = ~new_n7014 & ~new_n7015 ;
  assign new_n7017 = ~new_n7013 & new_n7016 ;
  assign new_n7018 = lo1371 & new_n3267 ;
  assign new_n7019 = lo1373 & new_n3270 ;
  assign new_n7020 = lo0339 & new_n3274 ;
  assign new_n7021 = ~new_n7019 & ~new_n7020 ;
  assign new_n7022 = ~new_n7018 & new_n7021 ;
  assign new_n7023 = ~new_n3265 & new_n7022 ;
  assign new_n7024 = new_n7017 & new_n7023 ;
  assign new_n7025 = ~new_n7012 & new_n7024 ;
  assign new_n7026 = ~new_n7011 & new_n7025 ;
  assign new_n7027 = new_n3141 & ~new_n7026 ;
  assign new_n7028 = new_n3140 & ~new_n7027 ;
  assign new_n7029 = ~new_n3121 & ~new_n7028 ;
  assign new_n7030 = new_n3121 & new_n7028 ;
  assign new_n7031 = ~new_n7029 & ~new_n7030 ;
  assign new_n7032 = lo0332 & ~new_n7031 ;
  assign new_n7033 = ~lo0332 & new_n7029 ;
  assign new_n7034 = new_n3121 & new_n4981 ;
  assign new_n7035 = ~new_n7028 & new_n7034 ;
  assign new_n7036 = ~new_n7033 & ~new_n7035 ;
  assign new_n7037 = ~new_n7032 & new_n7036 ;
  assign new_n7038 = ~new_n3112 & new_n7037 ;
  assign new_n7039 = new_n3112 & ~new_n7037 ;
  assign new_n7040 = ~new_n7038 & ~new_n7039 ;
  assign new_n7041 = lo0786 & new_n2506 ;
  assign new_n7042 = lo0785 & new_n2831 ;
  assign new_n7043 = ~new_n2521 & ~new_n7042 ;
  assign new_n7044 = ~new_n7041 & new_n7043 ;
  assign new_n7045 = ~lo0252 & ~new_n7044 ;
  assign new_n7046 = lo0252 & new_n7044 ;
  assign new_n7047 = ~new_n7045 & ~new_n7046 ;
  assign new_n7048 = lo0784 & ~new_n7047 ;
  assign new_n7049 = ~lo0784 & new_n7045 ;
  assign new_n7050 = lo0252 & lo0787 ;
  assign new_n7051 = ~new_n7044 & new_n7050 ;
  assign new_n7052 = ~new_n7049 & ~new_n7051 ;
  assign new_n7053 = ~new_n7048 & new_n7052 ;
  assign new_n7054 = lo0794 & new_n2506 ;
  assign new_n7055 = lo0793 & new_n2522 ;
  assign new_n7056 = ~new_n2521 & ~new_n7055 ;
  assign new_n7057 = ~new_n7054 & new_n7056 ;
  assign new_n7058 = ~lo0251 & ~new_n7057 ;
  assign new_n7059 = lo0251 & new_n7057 ;
  assign new_n7060 = ~new_n7058 & ~new_n7059 ;
  assign new_n7061 = lo0792 & ~new_n7060 ;
  assign new_n7062 = ~lo0792 & new_n7058 ;
  assign new_n7063 = lo0251 & lo0795 ;
  assign new_n7064 = ~new_n7057 & new_n7063 ;
  assign new_n7065 = ~new_n7062 & ~new_n7064 ;
  assign new_n7066 = ~new_n7061 & new_n7065 ;
  assign new_n7067 = new_n2490 & ~new_n7066 ;
  assign new_n7068 = lo0790 & new_n2506 ;
  assign new_n7069 = lo0789 & new_n2522 ;
  assign new_n7070 = ~new_n2521 & ~new_n7069 ;
  assign new_n7071 = ~new_n7068 & new_n7070 ;
  assign new_n7072 = ~lo0251 & ~new_n7071 ;
  assign new_n7073 = lo0251 & new_n7071 ;
  assign new_n7074 = ~new_n7072 & ~new_n7073 ;
  assign new_n7075 = lo0788 & ~new_n7074 ;
  assign new_n7076 = ~lo0788 & new_n7072 ;
  assign new_n7077 = lo0251 & lo0791 ;
  assign new_n7078 = ~new_n7071 & new_n7077 ;
  assign new_n7079 = ~new_n7076 & ~new_n7078 ;
  assign new_n7080 = ~new_n7075 & new_n7079 ;
  assign new_n7081 = new_n3310 & ~new_n7080 ;
  assign new_n7082 = ~new_n2492 & ~new_n7081 ;
  assign new_n7083 = ~new_n7067 & new_n7082 ;
  assign new_n7084 = ~lo0250 & ~new_n7083 ;
  assign new_n7085 = lo0250 & new_n7083 ;
  assign new_n7086 = ~new_n7084 & ~new_n7085 ;
  assign new_n7087 = ~new_n7053 & ~new_n7086 ;
  assign new_n7088 = new_n7053 & new_n7084 ;
  assign new_n7089 = lo0798 & new_n2506 ;
  assign new_n7090 = lo0797 & new_n2831 ;
  assign new_n7091 = ~new_n2521 & ~new_n7090 ;
  assign new_n7092 = ~new_n7089 & new_n7091 ;
  assign new_n7093 = ~lo0252 & ~new_n7092 ;
  assign new_n7094 = lo0252 & new_n7092 ;
  assign new_n7095 = ~new_n7093 & ~new_n7094 ;
  assign new_n7096 = lo0796 & ~new_n7095 ;
  assign new_n7097 = ~lo0796 & new_n7093 ;
  assign new_n7098 = lo0252 & lo0799 ;
  assign new_n7099 = ~new_n7092 & new_n7098 ;
  assign new_n7100 = ~new_n7097 & ~new_n7099 ;
  assign new_n7101 = ~new_n7096 & new_n7100 ;
  assign new_n7102 = lo0250 & ~new_n7101 ;
  assign new_n7103 = ~new_n7083 & new_n7102 ;
  assign new_n7104 = ~new_n7088 & ~new_n7103 ;
  assign new_n7105 = ~new_n7087 & new_n7104 ;
  assign new_n7106 = new_n2489 & ~new_n7105 ;
  assign new_n7107 = lo0801 & new_n2565 ;
  assign new_n7108 = new_n2569 & new_n7107 ;
  assign new_n7109 = lo0800 & new_n2565 ;
  assign new_n7110 = ~new_n2569 & new_n7109 ;
  assign new_n7111 = ~new_n2572 & ~new_n7110 ;
  assign new_n7112 = ~new_n7108 & new_n7111 ;
  assign new_n7113 = new_n2565 & ~new_n7112 ;
  assign new_n7114 = ~new_n2565 & new_n7112 ;
  assign new_n7115 = ~new_n7113 & ~new_n7114 ;
  assign new_n7116 = lo0780 & ~new_n7115 ;
  assign new_n7117 = ~lo0780 & new_n7113 ;
  assign new_n7118 = lo0802 & ~new_n2565 ;
  assign new_n7119 = ~new_n7112 & new_n7118 ;
  assign new_n7120 = ~new_n7117 & ~new_n7119 ;
  assign new_n7121 = ~new_n7116 & new_n7120 ;
  assign new_n7122 = lo0090 & ~new_n7121 ;
  assign new_n7123 = ~new_n2483 & new_n7122 ;
  assign new_n7124 = ~lo0106 & lo0641 ;
  assign new_n7125 = ~new_n6674 & new_n7124 ;
  assign new_n7126 = lo0579 & ~new_n2597 ;
  assign new_n7127 = ~new_n7125 & ~new_n7126 ;
  assign new_n7128 = new_n2591 & ~new_n7127 ;
  assign new_n7129 = lo0803 & new_n2601 ;
  assign new_n7130 = lo0804 & new_n2605 ;
  assign new_n7131 = ~new_n7129 & ~new_n7130 ;
  assign new_n7132 = lo1380 & new_n2610 ;
  assign new_n7133 = lo0805 & new_n2613 ;
  assign new_n7134 = ~new_n7132 & ~new_n7133 ;
  assign new_n7135 = new_n7131 & new_n7134 ;
  assign new_n7136 = ~new_n7128 & new_n7135 ;
  assign new_n7137 = ~new_n7123 & new_n7136 ;
  assign new_n7138 = ~new_n7106 & new_n7137 ;
  assign new_n7139 = new_n3820 & ~new_n5560 ;
  assign new_n7140 = ~new_n2910 & new_n3737 ;
  assign new_n7141 = ~new_n3819 & ~new_n7140 ;
  assign new_n7142 = ~new_n7139 & new_n7141 ;
  assign new_n7143 = ~new_n3735 & ~new_n7142 ;
  assign new_n7144 = new_n3735 & new_n7142 ;
  assign new_n7145 = ~new_n7143 & ~new_n7144 ;
  assign new_n7146 = ~new_n7138 & ~new_n7145 ;
  assign new_n7147 = new_n7138 & new_n7143 ;
  assign new_n7148 = new_n3735 & ~new_n5187 ;
  assign new_n7149 = ~new_n7142 & new_n7148 ;
  assign new_n7150 = ~new_n7147 & ~new_n7149 ;
  assign new_n7151 = ~new_n7146 & new_n7150 ;
  assign new_n7152 = new_n5673 & new_n7151 ;
  assign new_n7153 = ~new_n5782 & ~new_n7151 ;
  assign new_n7154 = ~new_n4992 & new_n5784 ;
  assign new_n7155 = ~new_n7153 & ~new_n7154 ;
  assign new_n7156 = ~new_n7152 & new_n7155 ;
  assign new_n7157 = ~new_n5672 & ~new_n7156 ;
  assign new_n7158 = new_n5672 & new_n7156 ;
  assign new_n7159 = ~new_n7157 & ~new_n7158 ;
  assign new_n7160 = ~new_n4630 & ~new_n7159 ;
  assign new_n7161 = new_n4630 & new_n7157 ;
  assign new_n7162 = ~new_n4541 & new_n5672 ;
  assign new_n7163 = ~new_n7156 & new_n7162 ;
  assign new_n7164 = ~new_n7161 & ~new_n7163 ;
  assign new_n7165 = ~new_n7160 & new_n7164 ;
  assign new_n7166 = new_n3102 & ~new_n7165 ;
  assign new_n7167 = ~new_n3102 & ~new_n5276 ;
  assign new_n7168 = ~new_n7166 & ~new_n7167 ;
  assign new_n7169 = lo0766 & new_n3170 ;
  assign new_n7170 = lo0765 & new_n3173 ;
  assign new_n7171 = ~new_n3172 & ~new_n7170 ;
  assign new_n7172 = ~new_n7169 & new_n7171 ;
  assign new_n7173 = ~lo0059 & ~new_n7172 ;
  assign new_n7174 = lo0059 & new_n7172 ;
  assign new_n7175 = ~new_n7173 & ~new_n7174 ;
  assign new_n7176 = lo0764 & ~new_n7175 ;
  assign new_n7177 = ~lo0764 & new_n7173 ;
  assign new_n7178 = lo0059 & lo0767 ;
  assign new_n7179 = ~new_n7172 & new_n7178 ;
  assign new_n7180 = ~new_n7177 & ~new_n7179 ;
  assign new_n7181 = ~new_n7176 & new_n7180 ;
  assign new_n7182 = lo0774 & new_n3170 ;
  assign new_n7183 = lo0773 & new_n3204 ;
  assign new_n7184 = ~new_n3172 & ~new_n7183 ;
  assign new_n7185 = ~new_n7182 & new_n7184 ;
  assign new_n7186 = ~lo0061 & ~new_n7185 ;
  assign new_n7187 = lo0061 & new_n7185 ;
  assign new_n7188 = ~new_n7186 & ~new_n7187 ;
  assign new_n7189 = lo0772 & ~new_n7188 ;
  assign new_n7190 = ~lo0772 & new_n7186 ;
  assign new_n7191 = lo0061 & lo0775 ;
  assign new_n7192 = ~new_n7185 & new_n7191 ;
  assign new_n7193 = ~new_n7190 & ~new_n7192 ;
  assign new_n7194 = ~new_n7189 & new_n7193 ;
  assign new_n7195 = new_n3186 & ~new_n7194 ;
  assign new_n7196 = lo0770 & new_n3170 ;
  assign new_n7197 = lo0769 & new_n3204 ;
  assign new_n7198 = ~new_n3172 & ~new_n7197 ;
  assign new_n7199 = ~new_n7196 & new_n7198 ;
  assign new_n7200 = ~lo0061 & ~new_n7199 ;
  assign new_n7201 = lo0061 & new_n7199 ;
  assign new_n7202 = ~new_n7200 & ~new_n7201 ;
  assign new_n7203 = lo0768 & ~new_n7202 ;
  assign new_n7204 = ~lo0768 & new_n7200 ;
  assign new_n7205 = lo0061 & lo0771 ;
  assign new_n7206 = ~new_n7199 & new_n7205 ;
  assign new_n7207 = ~new_n7204 & ~new_n7206 ;
  assign new_n7208 = ~new_n7203 & new_n7207 ;
  assign new_n7209 = new_n3559 & ~new_n7208 ;
  assign new_n7210 = ~new_n3201 & ~new_n7209 ;
  assign new_n7211 = ~new_n7195 & new_n7210 ;
  assign new_n7212 = ~lo0065 & ~new_n7211 ;
  assign new_n7213 = lo0065 & new_n7211 ;
  assign new_n7214 = ~new_n7212 & ~new_n7213 ;
  assign new_n7215 = ~new_n7181 & ~new_n7214 ;
  assign new_n7216 = new_n7181 & new_n7212 ;
  assign new_n7217 = lo0778 & new_n3170 ;
  assign new_n7218 = lo0777 & new_n3173 ;
  assign new_n7219 = ~new_n3172 & ~new_n7218 ;
  assign new_n7220 = ~new_n7217 & new_n7219 ;
  assign new_n7221 = ~lo0059 & ~new_n7220 ;
  assign new_n7222 = lo0059 & new_n7220 ;
  assign new_n7223 = ~new_n7221 & ~new_n7222 ;
  assign new_n7224 = lo0776 & ~new_n7223 ;
  assign new_n7225 = ~lo0776 & new_n7221 ;
  assign new_n7226 = lo0059 & lo0779 ;
  assign new_n7227 = ~new_n7220 & new_n7226 ;
  assign new_n7228 = ~new_n7225 & ~new_n7227 ;
  assign new_n7229 = ~new_n7224 & new_n7228 ;
  assign new_n7230 = lo0065 & ~new_n7229 ;
  assign new_n7231 = ~new_n7211 & new_n7230 ;
  assign new_n7232 = ~new_n7216 & ~new_n7231 ;
  assign new_n7233 = ~new_n7215 & new_n7232 ;
  assign new_n7234 = new_n3169 & ~new_n7233 ;
  assign new_n7235 = ~new_n3160 & new_n5265 ;
  assign new_n7236 = lo1390 & new_n3246 ;
  assign new_n7237 = lo1367 & new_n3254 ;
  assign new_n7238 = lo0782 & new_n3258 ;
  assign new_n7239 = ~new_n7237 & ~new_n7238 ;
  assign new_n7240 = ~new_n7236 & new_n7239 ;
  assign new_n7241 = lo1389 & new_n3267 ;
  assign new_n7242 = lo1391 & new_n3270 ;
  assign new_n7243 = lo0781 & new_n3274 ;
  assign new_n7244 = ~new_n7242 & ~new_n7243 ;
  assign new_n7245 = ~new_n7241 & new_n7244 ;
  assign new_n7246 = ~new_n3265 & new_n7245 ;
  assign new_n7247 = new_n7240 & new_n7246 ;
  assign new_n7248 = ~new_n7235 & new_n7247 ;
  assign new_n7249 = ~new_n7234 & new_n7248 ;
  assign new_n7250 = new_n3141 & ~new_n7249 ;
  assign new_n7251 = new_n3140 & ~new_n7250 ;
  assign new_n7252 = ~new_n3121 & ~new_n7251 ;
  assign new_n7253 = new_n3121 & new_n7251 ;
  assign new_n7254 = ~new_n7252 & ~new_n7253 ;
  assign new_n7255 = lo0774 & ~new_n7254 ;
  assign new_n7256 = ~lo0774 & new_n7252 ;
  assign new_n7257 = new_n3121 & new_n5265 ;
  assign new_n7258 = ~new_n7251 & new_n7257 ;
  assign new_n7259 = ~new_n7256 & ~new_n7258 ;
  assign new_n7260 = ~new_n7255 & new_n7259 ;
  assign new_n7261 = ~new_n3112 & new_n7260 ;
  assign new_n7262 = new_n3112 & ~new_n7260 ;
  assign new_n7263 = ~new_n7261 & ~new_n7262 ;
  assign new_n7264 = ~new_n3383 & new_n3737 ;
  assign new_n7265 = ~new_n3819 & ~new_n7264 ;
  assign new_n7266 = ~new_n2619 & new_n4180 ;
  assign new_n7267 = new_n7265 & ~new_n7266 ;
  assign new_n7268 = new_n3736 & ~new_n7267 ;
  assign new_n7269 = ~new_n3736 & new_n7267 ;
  assign new_n7270 = ~new_n7268 & ~new_n7269 ;
  assign new_n7271 = ~new_n2910 & ~new_n7270 ;
  assign new_n7272 = new_n2910 & new_n7268 ;
  assign new_n7273 = ~new_n3736 & ~new_n5472 ;
  assign new_n7274 = ~new_n7267 & new_n7273 ;
  assign new_n7275 = ~new_n7272 & ~new_n7274 ;
  assign new_n7276 = ~new_n7271 & new_n7275 ;
  assign new_n7277 = new_n5673 & new_n7276 ;
  assign new_n7278 = ~new_n5782 & ~new_n7276 ;
  assign new_n7279 = ~new_n5276 & new_n5784 ;
  assign new_n7280 = ~new_n7278 & ~new_n7279 ;
  assign new_n7281 = ~new_n7277 & new_n7280 ;
  assign new_n7282 = ~new_n5672 & ~new_n7281 ;
  assign new_n7283 = new_n5672 & new_n7281 ;
  assign new_n7284 = ~new_n7282 & ~new_n7283 ;
  assign new_n7285 = ~new_n4992 & ~new_n7284 ;
  assign new_n7286 = new_n4992 & new_n7282 ;
  assign new_n7287 = ~new_n4818 & new_n5672 ;
  assign new_n7288 = ~new_n7281 & new_n7287 ;
  assign new_n7289 = ~new_n7286 & ~new_n7288 ;
  assign new_n7290 = ~new_n7285 & new_n7289 ;
  assign new_n7291 = new_n3102 & ~new_n7290 ;
  assign new_n7292 = ~new_n3102 & ~new_n5560 ;
  assign new_n7293 = ~new_n7291 & ~new_n7292 ;
  assign new_n7294 = lo0541 & new_n3186 ;
  assign new_n7295 = lo0540 & new_n3559 ;
  assign new_n7296 = ~new_n3201 & ~new_n7295 ;
  assign new_n7297 = ~new_n7294 & new_n7296 ;
  assign new_n7298 = ~lo0065 & ~new_n7297 ;
  assign new_n7299 = lo0065 & new_n7297 ;
  assign new_n7300 = ~new_n7298 & ~new_n7299 ;
  assign new_n7301 = lo0539 & ~new_n7300 ;
  assign new_n7302 = ~lo0539 & new_n7298 ;
  assign new_n7303 = lo0065 & lo0542 ;
  assign new_n7304 = ~new_n7297 & new_n7303 ;
  assign new_n7305 = ~new_n7302 & ~new_n7304 ;
  assign new_n7306 = ~new_n7301 & new_n7305 ;
  assign new_n7307 = lo0549 & new_n3186 ;
  assign new_n7308 = lo0548 & new_n3202 ;
  assign new_n7309 = ~new_n3201 & ~new_n7308 ;
  assign new_n7310 = ~new_n7307 & new_n7309 ;
  assign new_n7311 = ~lo0063 & ~new_n7310 ;
  assign new_n7312 = lo0063 & new_n7310 ;
  assign new_n7313 = ~new_n7311 & ~new_n7312 ;
  assign new_n7314 = lo0547 & ~new_n7313 ;
  assign new_n7315 = ~lo0547 & new_n7311 ;
  assign new_n7316 = lo0063 & lo0550 ;
  assign new_n7317 = ~new_n7310 & new_n7316 ;
  assign new_n7318 = ~new_n7315 & ~new_n7317 ;
  assign new_n7319 = ~new_n7314 & new_n7318 ;
  assign new_n7320 = new_n3170 & ~new_n7319 ;
  assign new_n7321 = lo0545 & new_n3186 ;
  assign new_n7322 = lo0544 & new_n3202 ;
  assign new_n7323 = ~new_n3201 & ~new_n7322 ;
  assign new_n7324 = ~new_n7321 & new_n7323 ;
  assign new_n7325 = ~lo0063 & ~new_n7324 ;
  assign new_n7326 = lo0063 & new_n7324 ;
  assign new_n7327 = ~new_n7325 & ~new_n7326 ;
  assign new_n7328 = lo0543 & ~new_n7327 ;
  assign new_n7329 = ~lo0543 & new_n7325 ;
  assign new_n7330 = lo0063 & lo0546 ;
  assign new_n7331 = ~new_n7324 & new_n7330 ;
  assign new_n7332 = ~new_n7329 & ~new_n7331 ;
  assign new_n7333 = ~new_n7328 & new_n7332 ;
  assign new_n7334 = new_n3204 & ~new_n7333 ;
  assign new_n7335 = ~new_n3172 & ~new_n7334 ;
  assign new_n7336 = ~new_n7320 & new_n7335 ;
  assign new_n7337 = ~lo0061 & ~new_n7336 ;
  assign new_n7338 = lo0061 & new_n7336 ;
  assign new_n7339 = ~new_n7337 & ~new_n7338 ;
  assign new_n7340 = ~new_n7306 & ~new_n7339 ;
  assign new_n7341 = new_n7306 & new_n7337 ;
  assign new_n7342 = lo0553 & new_n3186 ;
  assign new_n7343 = lo0552 & new_n3559 ;
  assign new_n7344 = ~new_n3201 & ~new_n7343 ;
  assign new_n7345 = ~new_n7342 & new_n7344 ;
  assign new_n7346 = ~lo0065 & ~new_n7345 ;
  assign new_n7347 = lo0065 & new_n7345 ;
  assign new_n7348 = ~new_n7346 & ~new_n7347 ;
  assign new_n7349 = lo0551 & ~new_n7348 ;
  assign new_n7350 = ~lo0551 & new_n7346 ;
  assign new_n7351 = lo0065 & lo0554 ;
  assign new_n7352 = ~new_n7345 & new_n7351 ;
  assign new_n7353 = ~new_n7350 & ~new_n7352 ;
  assign new_n7354 = ~new_n7349 & new_n7353 ;
  assign new_n7355 = lo0061 & ~new_n7354 ;
  assign new_n7356 = ~new_n7336 & new_n7355 ;
  assign new_n7357 = ~new_n7341 & ~new_n7356 ;
  assign new_n7358 = ~new_n7340 & new_n7357 ;
  assign new_n7359 = new_n3169 & ~new_n7358 ;
  assign new_n7360 = ~new_n3160 & new_n5549 ;
  assign new_n7361 = lo1365 & new_n3246 ;
  assign new_n7362 = lo1329 & new_n3254 ;
  assign new_n7363 = lo0557 & new_n3258 ;
  assign new_n7364 = ~new_n7362 & ~new_n7363 ;
  assign new_n7365 = ~new_n7361 & new_n7364 ;
  assign new_n7366 = lo1364 & new_n3267 ;
  assign new_n7367 = lo1366 & new_n3270 ;
  assign new_n7368 = lo0556 & new_n3274 ;
  assign new_n7369 = ~new_n7367 & ~new_n7368 ;
  assign new_n7370 = ~new_n7366 & new_n7369 ;
  assign new_n7371 = ~new_n3265 & new_n7370 ;
  assign new_n7372 = new_n7365 & new_n7371 ;
  assign new_n7373 = ~new_n7360 & new_n7372 ;
  assign new_n7374 = ~new_n7359 & new_n7373 ;
  assign new_n7375 = new_n3141 & ~new_n7374 ;
  assign new_n7376 = new_n3140 & ~new_n7375 ;
  assign new_n7377 = ~new_n3121 & ~new_n7376 ;
  assign new_n7378 = new_n3121 & new_n7376 ;
  assign new_n7379 = ~new_n7377 & ~new_n7378 ;
  assign new_n7380 = lo0549 & ~new_n7379 ;
  assign new_n7381 = ~lo0549 & new_n7377 ;
  assign new_n7382 = new_n3121 & new_n5549 ;
  assign new_n7383 = ~new_n7376 & new_n7382 ;
  assign new_n7384 = ~new_n7381 & ~new_n7383 ;
  assign new_n7385 = ~new_n7380 & new_n7384 ;
  assign new_n7386 = ~new_n3112 & new_n7385 ;
  assign new_n7387 = new_n3112 & ~new_n7385 ;
  assign new_n7388 = ~new_n7386 & ~new_n7387 ;
  assign new_n7389 = lo0300 & new_n2825 ;
  assign new_n7390 = ~lo0298 & ~new_n7389 ;
  assign new_n7391 = lo0299 & new_n7390 ;
  assign new_n7392 = new_n2825 & ~new_n7391 ;
  assign new_n7393 = new_n6692 & ~new_n7139 ;
  assign new_n7394 = ~new_n3735 & ~new_n7393 ;
  assign new_n7395 = new_n3735 & new_n7393 ;
  assign new_n7396 = ~new_n7394 & ~new_n7395 ;
  assign new_n7397 = ~new_n2739 & ~new_n7396 ;
  assign new_n7398 = new_n2739 & new_n7394 ;
  assign new_n7399 = ~new_n2824 & new_n3735 ;
  assign new_n7400 = ~new_n7393 & new_n7399 ;
  assign new_n7401 = ~new_n7398 & ~new_n7400 ;
  assign new_n7402 = ~new_n7397 & new_n7401 ;
  assign new_n7403 = ~new_n2825 & ~new_n7390 ;
  assign new_n7404 = ~new_n7402 & new_n7403 ;
  assign new_n7405 = new_n2825 & ~new_n7390 ;
  assign new_n7406 = ~new_n2825 & new_n7390 ;
  assign new_n7407 = ~new_n7405 & ~new_n7406 ;
  assign new_n7408 = ~new_n3383 & ~new_n7407 ;
  assign new_n7409 = new_n3383 & new_n7405 ;
  assign new_n7410 = ~new_n7408 & ~new_n7409 ;
  assign new_n7411 = ~new_n7404 & new_n7410 ;
  assign new_n7412 = ~new_n7392 & ~new_n7411 ;
  assign new_n7413 = new_n7392 & new_n7411 ;
  assign new_n7414 = ~new_n7412 & ~new_n7413 ;
  assign new_n7415 = ~new_n3734 & ~new_n7414 ;
  assign new_n7416 = new_n3734 & new_n7412 ;
  assign new_n7417 = ~new_n5766 & new_n7392 ;
  assign new_n7418 = ~new_n7411 & new_n7417 ;
  assign new_n7419 = ~new_n7416 & ~new_n7418 ;
  assign new_n7420 = ~new_n7415 & new_n7419 ;
  assign new_n7421 = new_n3102 & ~new_n7420 ;
  assign new_n7422 = ~new_n2910 & ~new_n3102 ;
  assign new_n7423 = ~new_n7421 & ~new_n7422 ;
  assign new_n7424 = ~lo0065 & lo0404 ;
  assign new_n7425 = ~lo0063 & new_n7424 ;
  assign new_n7426 = ~lo0065 & lo0403 ;
  assign new_n7427 = lo0063 & new_n7426 ;
  assign new_n7428 = ~new_n3201 & ~new_n7427 ;
  assign new_n7429 = ~new_n7425 & new_n7428 ;
  assign new_n7430 = ~lo0065 & ~new_n7429 ;
  assign new_n7431 = lo0065 & new_n7429 ;
  assign new_n7432 = ~new_n7430 & ~new_n7431 ;
  assign new_n7433 = lo0402 & ~new_n7432 ;
  assign new_n7434 = ~lo0402 & new_n7430 ;
  assign new_n7435 = lo0065 & lo0405 ;
  assign new_n7436 = ~new_n7429 & new_n7435 ;
  assign new_n7437 = ~new_n7434 & ~new_n7436 ;
  assign new_n7438 = ~new_n7433 & new_n7437 ;
  assign new_n7439 = ~lo0065 & lo0401 ;
  assign new_n7440 = ~lo0063 & new_n7439 ;
  assign new_n7441 = ~lo0065 & lo0411 ;
  assign new_n7442 = lo0063 & new_n7441 ;
  assign new_n7443 = ~new_n3201 & ~new_n7442 ;
  assign new_n7444 = ~new_n7440 & new_n7443 ;
  assign new_n7445 = ~lo0065 & ~new_n7444 ;
  assign new_n7446 = lo0065 & new_n7444 ;
  assign new_n7447 = ~new_n7445 & ~new_n7446 ;
  assign new_n7448 = lo0410 & ~new_n7447 ;
  assign new_n7449 = ~lo0410 & new_n7445 ;
  assign new_n7450 = lo0065 & lo0412 ;
  assign new_n7451 = ~new_n7444 & new_n7450 ;
  assign new_n7452 = ~new_n7449 & ~new_n7451 ;
  assign new_n7453 = ~new_n7448 & new_n7452 ;
  assign new_n7454 = new_n3170 & ~new_n7453 ;
  assign new_n7455 = ~lo0063 & lo0408 ;
  assign new_n7456 = ~lo0065 & new_n7455 ;
  assign new_n7457 = ~lo0063 & lo0407 ;
  assign new_n7458 = lo0065 & new_n7457 ;
  assign new_n7459 = ~new_n3201 & ~new_n7458 ;
  assign new_n7460 = ~new_n7456 & new_n7459 ;
  assign new_n7461 = ~lo0063 & ~new_n7460 ;
  assign new_n7462 = lo0063 & new_n7460 ;
  assign new_n7463 = ~new_n7461 & ~new_n7462 ;
  assign new_n7464 = lo0406 & ~new_n7463 ;
  assign new_n7465 = ~lo0406 & new_n7461 ;
  assign new_n7466 = lo0063 & lo0409 ;
  assign new_n7467 = ~new_n7460 & new_n7466 ;
  assign new_n7468 = ~new_n7465 & ~new_n7467 ;
  assign new_n7469 = ~new_n7464 & new_n7468 ;
  assign new_n7470 = new_n3173 & ~new_n7469 ;
  assign new_n7471 = ~new_n3172 & ~new_n7470 ;
  assign new_n7472 = ~new_n7454 & new_n7471 ;
  assign new_n7473 = ~lo0059 & ~new_n7472 ;
  assign new_n7474 = lo0059 & new_n7472 ;
  assign new_n7475 = ~new_n7473 & ~new_n7474 ;
  assign new_n7476 = ~new_n7438 & ~new_n7475 ;
  assign new_n7477 = new_n7438 & new_n7473 ;
  assign new_n7478 = ~lo0063 & lo0415 ;
  assign new_n7479 = ~lo0065 & new_n7478 ;
  assign new_n7480 = ~lo0063 & lo0414 ;
  assign new_n7481 = lo0065 & new_n7480 ;
  assign new_n7482 = ~new_n3201 & ~new_n7481 ;
  assign new_n7483 = ~new_n7479 & new_n7482 ;
  assign new_n7484 = ~lo0063 & ~new_n7483 ;
  assign new_n7485 = lo0063 & new_n7483 ;
  assign new_n7486 = ~new_n7484 & ~new_n7485 ;
  assign new_n7487 = lo0413 & ~new_n7486 ;
  assign new_n7488 = ~lo0413 & new_n7484 ;
  assign new_n7489 = lo0063 & lo0416 ;
  assign new_n7490 = ~new_n7483 & new_n7489 ;
  assign new_n7491 = ~new_n7488 & ~new_n7490 ;
  assign new_n7492 = ~new_n7487 & new_n7491 ;
  assign new_n7493 = lo0059 & ~new_n7492 ;
  assign new_n7494 = ~new_n7472 & new_n7493 ;
  assign new_n7495 = ~new_n7477 & ~new_n7494 ;
  assign new_n7496 = ~new_n7476 & new_n7495 ;
  assign new_n7497 = new_n3169 & ~new_n7496 ;
  assign new_n7498 = new_n2899 & ~new_n3160 ;
  assign new_n7499 = lo1315 & new_n3246 ;
  assign new_n7500 = lo1314 & new_n3254 ;
  assign new_n7501 = lo0418 & new_n3258 ;
  assign new_n7502 = ~new_n7500 & ~new_n7501 ;
  assign new_n7503 = ~new_n7499 & new_n7502 ;
  assign new_n7504 = lo1313 & new_n3267 ;
  assign new_n7505 = lo1316 & new_n3270 ;
  assign new_n7506 = lo0417 & new_n3274 ;
  assign new_n7507 = ~new_n7505 & ~new_n7506 ;
  assign new_n7508 = ~new_n7504 & new_n7507 ;
  assign new_n7509 = ~new_n3265 & new_n7508 ;
  assign new_n7510 = new_n7503 & new_n7509 ;
  assign new_n7511 = ~new_n7498 & new_n7510 ;
  assign new_n7512 = ~new_n7497 & new_n7511 ;
  assign new_n7513 = new_n3141 & ~new_n7512 ;
  assign new_n7514 = new_n3140 & ~new_n7513 ;
  assign new_n7515 = ~new_n3121 & ~new_n7514 ;
  assign new_n7516 = new_n3121 & new_n7514 ;
  assign new_n7517 = ~new_n7515 & ~new_n7516 ;
  assign new_n7518 = lo0401 & ~new_n7517 ;
  assign new_n7519 = ~lo0401 & new_n7515 ;
  assign new_n7520 = new_n2899 & new_n3121 ;
  assign new_n7521 = ~new_n7514 & new_n7520 ;
  assign new_n7522 = ~new_n7519 & ~new_n7521 ;
  assign new_n7523 = ~new_n7518 & new_n7522 ;
  assign new_n7524 = ~new_n3112 & new_n7523 ;
  assign new_n7525 = new_n3112 & ~new_n7523 ;
  assign new_n7526 = ~new_n7524 & ~new_n7525 ;
  assign new_n7527 = ~new_n3092 & new_n4180 ;
  assign new_n7528 = new_n6817 & ~new_n7527 ;
  assign new_n7529 = new_n3736 & ~new_n7528 ;
  assign new_n7530 = ~new_n3736 & new_n7528 ;
  assign new_n7531 = ~new_n7529 & ~new_n7530 ;
  assign new_n7532 = ~new_n2910 & ~new_n7531 ;
  assign new_n7533 = new_n2910 & new_n7529 ;
  assign new_n7534 = ~new_n3549 & ~new_n3736 ;
  assign new_n7535 = ~new_n7528 & new_n7534 ;
  assign new_n7536 = ~new_n7533 & ~new_n7535 ;
  assign new_n7537 = ~new_n7532 & new_n7536 ;
  assign new_n7538 = new_n7403 & ~new_n7537 ;
  assign new_n7539 = ~new_n3734 & ~new_n7407 ;
  assign new_n7540 = new_n3734 & new_n7405 ;
  assign new_n7541 = ~new_n7539 & ~new_n7540 ;
  assign new_n7542 = ~new_n7538 & new_n7541 ;
  assign new_n7543 = ~new_n7392 & ~new_n7542 ;
  assign new_n7544 = new_n7392 & new_n7542 ;
  assign new_n7545 = ~new_n7543 & ~new_n7544 ;
  assign new_n7546 = ~new_n4179 & ~new_n7545 ;
  assign new_n7547 = new_n4179 & new_n7543 ;
  assign new_n7548 = ~new_n5996 & new_n7392 ;
  assign new_n7549 = ~new_n7542 & new_n7548 ;
  assign new_n7550 = ~new_n7547 & ~new_n7549 ;
  assign new_n7551 = ~new_n7546 & new_n7550 ;
  assign new_n7552 = new_n3102 & ~new_n7551 ;
  assign new_n7553 = ~new_n3102 & ~new_n3383 ;
  assign new_n7554 = ~new_n7552 & ~new_n7553 ;
  assign new_n7555 = lo0421 & new_n3170 ;
  assign new_n7556 = lo0420 & new_n3173 ;
  assign new_n7557 = ~new_n3172 & ~new_n7556 ;
  assign new_n7558 = ~new_n7555 & new_n7557 ;
  assign new_n7559 = ~lo0059 & ~new_n7558 ;
  assign new_n7560 = lo0059 & new_n7558 ;
  assign new_n7561 = ~new_n7559 & ~new_n7560 ;
  assign new_n7562 = lo0419 & ~new_n7561 ;
  assign new_n7563 = ~lo0419 & new_n7559 ;
  assign new_n7564 = lo0059 & lo0422 ;
  assign new_n7565 = ~new_n7558 & new_n7564 ;
  assign new_n7566 = ~new_n7563 & ~new_n7565 ;
  assign new_n7567 = ~new_n7562 & new_n7566 ;
  assign new_n7568 = lo0429 & new_n3170 ;
  assign new_n7569 = ~lo0061 & lo0428 ;
  assign new_n7570 = lo0059 & new_n7569 ;
  assign new_n7571 = ~new_n3172 & ~new_n7570 ;
  assign new_n7572 = ~new_n7568 & new_n7571 ;
  assign new_n7573 = ~lo0061 & ~new_n7572 ;
  assign new_n7574 = lo0061 & new_n7572 ;
  assign new_n7575 = ~new_n7573 & ~new_n7574 ;
  assign new_n7576 = lo0427 & ~new_n7575 ;
  assign new_n7577 = ~lo0427 & new_n7573 ;
  assign new_n7578 = lo0061 & lo0430 ;
  assign new_n7579 = ~new_n7572 & new_n7578 ;
  assign new_n7580 = ~new_n7577 & ~new_n7579 ;
  assign new_n7581 = ~new_n7576 & new_n7580 ;
  assign new_n7582 = new_n3186 & ~new_n7581 ;
  assign new_n7583 = lo0425 & new_n3170 ;
  assign new_n7584 = ~lo0061 & lo0424 ;
  assign new_n7585 = lo0059 & new_n7584 ;
  assign new_n7586 = ~new_n3172 & ~new_n7585 ;
  assign new_n7587 = ~new_n7583 & new_n7586 ;
  assign new_n7588 = ~lo0061 & ~new_n7587 ;
  assign new_n7589 = lo0061 & new_n7587 ;
  assign new_n7590 = ~new_n7588 & ~new_n7589 ;
  assign new_n7591 = lo0423 & ~new_n7590 ;
  assign new_n7592 = ~lo0423 & new_n7588 ;
  assign new_n7593 = lo0061 & lo0426 ;
  assign new_n7594 = ~new_n7587 & new_n7593 ;
  assign new_n7595 = ~new_n7592 & ~new_n7594 ;
  assign new_n7596 = ~new_n7591 & new_n7595 ;
  assign new_n7597 = new_n3559 & ~new_n7596 ;
  assign new_n7598 = ~new_n3201 & ~new_n7597 ;
  assign new_n7599 = ~new_n7582 & new_n7598 ;
  assign new_n7600 = ~lo0065 & ~new_n7599 ;
  assign new_n7601 = lo0065 & new_n7599 ;
  assign new_n7602 = ~new_n7600 & ~new_n7601 ;
  assign new_n7603 = ~new_n7567 & ~new_n7602 ;
  assign new_n7604 = new_n7567 & new_n7600 ;
  assign new_n7605 = lo0433 & new_n3170 ;
  assign new_n7606 = lo0432 & new_n3173 ;
  assign new_n7607 = ~new_n3172 & ~new_n7606 ;
  assign new_n7608 = ~new_n7605 & new_n7607 ;
  assign new_n7609 = ~lo0059 & ~new_n7608 ;
  assign new_n7610 = lo0059 & new_n7608 ;
  assign new_n7611 = ~new_n7609 & ~new_n7610 ;
  assign new_n7612 = lo0431 & ~new_n7611 ;
  assign new_n7613 = ~lo0431 & new_n7609 ;
  assign new_n7614 = lo0059 & lo0434 ;
  assign new_n7615 = ~new_n7608 & new_n7614 ;
  assign new_n7616 = ~new_n7613 & ~new_n7615 ;
  assign new_n7617 = ~new_n7612 & new_n7616 ;
  assign new_n7618 = lo0065 & ~new_n7617 ;
  assign new_n7619 = ~new_n7599 & new_n7618 ;
  assign new_n7620 = ~new_n7604 & ~new_n7619 ;
  assign new_n7621 = ~new_n7603 & new_n7620 ;
  assign new_n7622 = new_n3169 & ~new_n7621 ;
  assign new_n7623 = ~new_n3160 & ~new_n3372 ;
  assign new_n7624 = lo1326 & new_n3246 ;
  assign new_n7625 = lo1317 & new_n3254 ;
  assign new_n7626 = lo0438 & new_n3258 ;
  assign new_n7627 = ~new_n7625 & ~new_n7626 ;
  assign new_n7628 = ~new_n7624 & new_n7627 ;
  assign new_n7629 = lo1325 & new_n3267 ;
  assign new_n7630 = lo1327 & new_n3270 ;
  assign new_n7631 = lo0437 & new_n3274 ;
  assign new_n7632 = ~new_n7630 & ~new_n7631 ;
  assign new_n7633 = ~new_n7629 & new_n7632 ;
  assign new_n7634 = ~new_n3265 & new_n7633 ;
  assign new_n7635 = new_n7628 & new_n7634 ;
  assign new_n7636 = ~new_n7623 & new_n7635 ;
  assign new_n7637 = ~new_n7622 & new_n7636 ;
  assign new_n7638 = new_n3141 & ~new_n7637 ;
  assign new_n7639 = new_n3140 & ~new_n7638 ;
  assign new_n7640 = ~new_n3121 & ~new_n7639 ;
  assign new_n7641 = new_n3121 & new_n7639 ;
  assign new_n7642 = ~new_n7640 & ~new_n7641 ;
  assign new_n7643 = lo0429 & ~new_n7642 ;
  assign new_n7644 = ~lo0429 & new_n7640 ;
  assign new_n7645 = new_n3121 & ~new_n3372 ;
  assign new_n7646 = ~new_n7639 & new_n7645 ;
  assign new_n7647 = ~new_n7644 & ~new_n7646 ;
  assign new_n7648 = ~new_n7643 & new_n7647 ;
  assign new_n7649 = ~new_n3112 & new_n7648 ;
  assign new_n7650 = new_n3112 & ~new_n7648 ;
  assign new_n7651 = ~new_n7649 & ~new_n7650 ;
  assign new_n7652 = ~new_n3383 & new_n3820 ;
  assign new_n7653 = new_n7141 & ~new_n7652 ;
  assign new_n7654 = ~new_n3735 & ~new_n7653 ;
  assign new_n7655 = new_n3735 & new_n7653 ;
  assign new_n7656 = ~new_n7654 & ~new_n7655 ;
  assign new_n7657 = ~new_n3001 & ~new_n7656 ;
  assign new_n7658 = new_n3001 & new_n7654 ;
  assign new_n7659 = new_n3909 & ~new_n7653 ;
  assign new_n7660 = ~new_n7658 & ~new_n7659 ;
  assign new_n7661 = ~new_n7657 & new_n7660 ;
  assign new_n7662 = new_n7403 & ~new_n7661 ;
  assign new_n7663 = ~new_n4179 & ~new_n7407 ;
  assign new_n7664 = new_n4179 & new_n7405 ;
  assign new_n7665 = ~new_n7663 & ~new_n7664 ;
  assign new_n7666 = ~new_n7662 & new_n7665 ;
  assign new_n7667 = ~new_n7392 & ~new_n7666 ;
  assign new_n7668 = new_n7392 & new_n7666 ;
  assign new_n7669 = ~new_n7667 & ~new_n7668 ;
  assign new_n7670 = ~new_n4461 & ~new_n7669 ;
  assign new_n7671 = new_n4461 & new_n7667 ;
  assign new_n7672 = ~new_n6225 & new_n7392 ;
  assign new_n7673 = ~new_n7666 & new_n7672 ;
  assign new_n7674 = ~new_n7671 & ~new_n7673 ;
  assign new_n7675 = ~new_n7670 & new_n7674 ;
  assign new_n7676 = new_n3102 & ~new_n7675 ;
  assign new_n7677 = ~new_n3102 & ~new_n3734 ;
  assign new_n7678 = ~new_n7676 & ~new_n7677 ;
  assign new_n7679 = lo0520 & new_n3186 ;
  assign new_n7680 = lo0519 & new_n3559 ;
  assign new_n7681 = ~new_n3201 & ~new_n7680 ;
  assign new_n7682 = ~new_n7679 & new_n7681 ;
  assign new_n7683 = ~lo0065 & ~new_n7682 ;
  assign new_n7684 = lo0065 & new_n7682 ;
  assign new_n7685 = ~new_n7683 & ~new_n7684 ;
  assign new_n7686 = lo0518 & ~new_n7685 ;
  assign new_n7687 = ~lo0518 & new_n7683 ;
  assign new_n7688 = lo0065 & lo0521 ;
  assign new_n7689 = ~new_n7682 & new_n7688 ;
  assign new_n7690 = ~new_n7687 & ~new_n7689 ;
  assign new_n7691 = ~new_n7686 & new_n7690 ;
  assign new_n7692 = lo0528 & new_n3186 ;
  assign new_n7693 = ~lo0063 & lo0527 ;
  assign new_n7694 = lo0065 & new_n7693 ;
  assign new_n7695 = ~new_n3201 & ~new_n7694 ;
  assign new_n7696 = ~new_n7692 & new_n7695 ;
  assign new_n7697 = ~lo0063 & ~new_n7696 ;
  assign new_n7698 = lo0063 & new_n7696 ;
  assign new_n7699 = ~new_n7697 & ~new_n7698 ;
  assign new_n7700 = lo0526 & ~new_n7699 ;
  assign new_n7701 = ~lo0526 & new_n7697 ;
  assign new_n7702 = lo0063 & lo0529 ;
  assign new_n7703 = ~new_n7696 & new_n7702 ;
  assign new_n7704 = ~new_n7701 & ~new_n7703 ;
  assign new_n7705 = ~new_n7700 & new_n7704 ;
  assign new_n7706 = new_n3170 & ~new_n7705 ;
  assign new_n7707 = lo0524 & new_n3186 ;
  assign new_n7708 = ~lo0063 & lo0523 ;
  assign new_n7709 = lo0065 & new_n7708 ;
  assign new_n7710 = ~new_n3201 & ~new_n7709 ;
  assign new_n7711 = ~new_n7707 & new_n7710 ;
  assign new_n7712 = ~lo0063 & ~new_n7711 ;
  assign new_n7713 = lo0063 & new_n7711 ;
  assign new_n7714 = ~new_n7712 & ~new_n7713 ;
  assign new_n7715 = lo0522 & ~new_n7714 ;
  assign new_n7716 = ~lo0522 & new_n7712 ;
  assign new_n7717 = lo0063 & lo0525 ;
  assign new_n7718 = ~new_n7711 & new_n7717 ;
  assign new_n7719 = ~new_n7716 & ~new_n7718 ;
  assign new_n7720 = ~new_n7715 & new_n7719 ;
  assign new_n7721 = new_n3204 & ~new_n7720 ;
  assign new_n7722 = ~new_n3172 & ~new_n7721 ;
  assign new_n7723 = ~new_n7706 & new_n7722 ;
  assign new_n7724 = ~lo0061 & ~new_n7723 ;
  assign new_n7725 = lo0061 & new_n7723 ;
  assign new_n7726 = ~new_n7724 & ~new_n7725 ;
  assign new_n7727 = ~new_n7691 & ~new_n7726 ;
  assign new_n7728 = new_n7691 & new_n7724 ;
  assign new_n7729 = lo0532 & new_n3186 ;
  assign new_n7730 = lo0531 & new_n3559 ;
  assign new_n7731 = ~new_n3201 & ~new_n7730 ;
  assign new_n7732 = ~new_n7729 & new_n7731 ;
  assign new_n7733 = ~lo0065 & ~new_n7732 ;
  assign new_n7734 = lo0065 & new_n7732 ;
  assign new_n7735 = ~new_n7733 & ~new_n7734 ;
  assign new_n7736 = lo0530 & ~new_n7735 ;
  assign new_n7737 = ~lo0530 & new_n7733 ;
  assign new_n7738 = lo0065 & lo0533 ;
  assign new_n7739 = ~new_n7732 & new_n7738 ;
  assign new_n7740 = ~new_n7737 & ~new_n7739 ;
  assign new_n7741 = ~new_n7736 & new_n7740 ;
  assign new_n7742 = lo0061 & ~new_n7741 ;
  assign new_n7743 = ~new_n7723 & new_n7742 ;
  assign new_n7744 = ~new_n7728 & ~new_n7743 ;
  assign new_n7745 = ~new_n7727 & new_n7744 ;
  assign new_n7746 = new_n3169 & ~new_n7745 ;
  assign new_n7747 = ~new_n3160 & ~new_n3723 ;
  assign new_n7748 = lo1339 & new_n3246 ;
  assign new_n7749 = lo1328 & new_n3254 ;
  assign new_n7750 = lo0536 & new_n3258 ;
  assign new_n7751 = ~new_n7749 & ~new_n7750 ;
  assign new_n7752 = ~new_n7748 & new_n7751 ;
  assign new_n7753 = lo1338 & new_n3267 ;
  assign new_n7754 = lo1340 & new_n3270 ;
  assign new_n7755 = lo0535 & new_n3274 ;
  assign new_n7756 = ~new_n7754 & ~new_n7755 ;
  assign new_n7757 = ~new_n7753 & new_n7756 ;
  assign new_n7758 = ~new_n3265 & new_n7757 ;
  assign new_n7759 = new_n7752 & new_n7758 ;
  assign new_n7760 = ~new_n7747 & new_n7759 ;
  assign new_n7761 = ~new_n7746 & new_n7760 ;
  assign new_n7762 = new_n3141 & ~new_n7761 ;
  assign new_n7763 = new_n3140 & ~new_n7762 ;
  assign new_n7764 = ~new_n3121 & ~new_n7763 ;
  assign new_n7765 = new_n3121 & new_n7763 ;
  assign new_n7766 = ~new_n7764 & ~new_n7765 ;
  assign new_n7767 = lo0528 & ~new_n7766 ;
  assign new_n7768 = ~lo0528 & new_n7764 ;
  assign new_n7769 = new_n3121 & ~new_n3723 ;
  assign new_n7770 = ~new_n7763 & new_n7769 ;
  assign new_n7771 = ~new_n7768 & ~new_n7770 ;
  assign new_n7772 = ~new_n7767 & new_n7771 ;
  assign new_n7773 = ~new_n3112 & new_n7772 ;
  assign new_n7774 = new_n3112 & ~new_n7772 ;
  assign new_n7775 = ~new_n7773 & ~new_n7774 ;
  assign new_n7776 = ~new_n3464 & new_n4180 ;
  assign new_n7777 = new_n7265 & ~new_n7776 ;
  assign new_n7778 = new_n3736 & ~new_n7777 ;
  assign new_n7779 = ~new_n3736 & new_n7777 ;
  assign new_n7780 = ~new_n7778 & ~new_n7779 ;
  assign new_n7781 = ~new_n3734 & ~new_n7780 ;
  assign new_n7782 = new_n3734 & new_n7778 ;
  assign new_n7783 = new_n4269 & ~new_n7777 ;
  assign new_n7784 = ~new_n7782 & ~new_n7783 ;
  assign new_n7785 = ~new_n7781 & new_n7784 ;
  assign new_n7786 = new_n7403 & ~new_n7785 ;
  assign new_n7787 = ~new_n4461 & ~new_n7407 ;
  assign new_n7788 = new_n4461 & new_n7405 ;
  assign new_n7789 = ~new_n7787 & ~new_n7788 ;
  assign new_n7790 = ~new_n7786 & new_n7789 ;
  assign new_n7791 = ~new_n7392 & ~new_n7790 ;
  assign new_n7792 = new_n7392 & new_n7790 ;
  assign new_n7793 = ~new_n7791 & ~new_n7792 ;
  assign new_n7794 = ~new_n4904 & ~new_n7793 ;
  assign new_n7795 = new_n4904 & new_n7791 ;
  assign new_n7796 = ~new_n6461 & new_n7392 ;
  assign new_n7797 = ~new_n7790 & new_n7796 ;
  assign new_n7798 = ~new_n7795 & ~new_n7797 ;
  assign new_n7799 = ~new_n7794 & new_n7798 ;
  assign new_n7800 = new_n3102 & ~new_n7799 ;
  assign new_n7801 = ~new_n3102 & ~new_n4179 ;
  assign new_n7802 = ~new_n7800 & ~new_n7801 ;
  assign new_n7803 = lo0344 & new_n3170 ;
  assign new_n7804 = lo0343 & new_n3173 ;
  assign new_n7805 = ~new_n3172 & ~new_n7804 ;
  assign new_n7806 = ~new_n7803 & new_n7805 ;
  assign new_n7807 = ~lo0059 & ~new_n7806 ;
  assign new_n7808 = lo0059 & new_n7806 ;
  assign new_n7809 = ~new_n7807 & ~new_n7808 ;
  assign new_n7810 = lo0342 & ~new_n7809 ;
  assign new_n7811 = ~lo0342 & new_n7807 ;
  assign new_n7812 = lo0059 & lo0345 ;
  assign new_n7813 = ~new_n7806 & new_n7812 ;
  assign new_n7814 = ~new_n7811 & ~new_n7813 ;
  assign new_n7815 = ~new_n7810 & new_n7814 ;
  assign new_n7816 = lo1307 & new_n3170 ;
  assign new_n7817 = lo0351 & new_n3173 ;
  assign new_n7818 = ~new_n3172 & ~new_n7817 ;
  assign new_n7819 = ~new_n7816 & new_n7818 ;
  assign new_n7820 = ~lo0059 & ~new_n7819 ;
  assign new_n7821 = lo0059 & new_n7819 ;
  assign new_n7822 = ~new_n7820 & ~new_n7821 ;
  assign new_n7823 = lo0350 & ~new_n7822 ;
  assign new_n7824 = ~lo0350 & new_n7820 ;
  assign new_n7825 = lo0059 & lo0352 ;
  assign new_n7826 = ~new_n7819 & new_n7825 ;
  assign new_n7827 = ~new_n7824 & ~new_n7826 ;
  assign new_n7828 = ~new_n7823 & new_n7827 ;
  assign new_n7829 = new_n3186 & ~new_n7828 ;
  assign new_n7830 = lo0348 & new_n3170 ;
  assign new_n7831 = lo0347 & new_n3204 ;
  assign new_n7832 = ~new_n3172 & ~new_n7831 ;
  assign new_n7833 = ~new_n7830 & new_n7832 ;
  assign new_n7834 = ~lo0061 & ~new_n7833 ;
  assign new_n7835 = lo0061 & new_n7833 ;
  assign new_n7836 = ~new_n7834 & ~new_n7835 ;
  assign new_n7837 = lo0346 & ~new_n7836 ;
  assign new_n7838 = ~lo0346 & new_n7834 ;
  assign new_n7839 = lo0061 & lo0349 ;
  assign new_n7840 = ~new_n7833 & new_n7839 ;
  assign new_n7841 = ~new_n7838 & ~new_n7840 ;
  assign new_n7842 = ~new_n7837 & new_n7841 ;
  assign new_n7843 = new_n3202 & ~new_n7842 ;
  assign new_n7844 = ~new_n3201 & ~new_n7843 ;
  assign new_n7845 = ~new_n7829 & new_n7844 ;
  assign new_n7846 = ~lo0063 & ~new_n7845 ;
  assign new_n7847 = lo0063 & new_n7845 ;
  assign new_n7848 = ~new_n7846 & ~new_n7847 ;
  assign new_n7849 = ~new_n7815 & ~new_n7848 ;
  assign new_n7850 = new_n7815 & new_n7846 ;
  assign new_n7851 = lo0355 & new_n3170 ;
  assign new_n7852 = lo0354 & new_n3204 ;
  assign new_n7853 = ~new_n3172 & ~new_n7852 ;
  assign new_n7854 = ~new_n7851 & new_n7853 ;
  assign new_n7855 = ~lo0061 & ~new_n7854 ;
  assign new_n7856 = lo0061 & new_n7854 ;
  assign new_n7857 = ~new_n7855 & ~new_n7856 ;
  assign new_n7858 = lo0353 & ~new_n7857 ;
  assign new_n7859 = ~lo0353 & new_n7855 ;
  assign new_n7860 = lo0061 & lo0356 ;
  assign new_n7861 = ~new_n7854 & new_n7860 ;
  assign new_n7862 = ~new_n7859 & ~new_n7861 ;
  assign new_n7863 = ~new_n7858 & new_n7862 ;
  assign new_n7864 = lo0063 & ~new_n7863 ;
  assign new_n7865 = ~new_n7845 & new_n7864 ;
  assign new_n7866 = ~new_n7850 & ~new_n7865 ;
  assign new_n7867 = ~new_n7849 & new_n7866 ;
  assign new_n7868 = new_n3169 & ~new_n7867 ;
  assign new_n7869 = ~new_n3160 & ~new_n4168 ;
  assign new_n7870 = lo1346 & new_n3246 ;
  assign new_n7871 = lo0360 & new_n3254 ;
  assign new_n7872 = lo0358 & new_n3258 ;
  assign new_n7873 = ~new_n7871 & ~new_n7872 ;
  assign new_n7874 = ~new_n7870 & new_n7873 ;
  assign new_n7875 = lo1345 & new_n3267 ;
  assign new_n7876 = lo1347 & new_n3270 ;
  assign new_n7877 = lo0357 & new_n3274 ;
  assign new_n7878 = ~new_n7876 & ~new_n7877 ;
  assign new_n7879 = ~new_n7875 & new_n7878 ;
  assign new_n7880 = ~new_n3265 & new_n7879 ;
  assign new_n7881 = new_n7874 & new_n7880 ;
  assign new_n7882 = ~new_n7869 & new_n7881 ;
  assign new_n7883 = ~new_n7868 & new_n7882 ;
  assign new_n7884 = new_n3141 & ~new_n7883 ;
  assign new_n7885 = new_n3140 & ~new_n7884 ;
  assign new_n7886 = ~new_n3121 & ~new_n7885 ;
  assign new_n7887 = new_n3121 & new_n7885 ;
  assign new_n7888 = ~new_n7886 & ~new_n7887 ;
  assign new_n7889 = lo1307 & ~new_n7888 ;
  assign new_n7890 = ~lo1307 & new_n7886 ;
  assign new_n7891 = new_n3121 & ~new_n4168 ;
  assign new_n7892 = ~new_n7885 & new_n7891 ;
  assign new_n7893 = ~new_n7890 & ~new_n7892 ;
  assign new_n7894 = ~new_n7889 & new_n7893 ;
  assign new_n7895 = ~new_n3112 & new_n7894 ;
  assign new_n7896 = new_n3112 & ~new_n7894 ;
  assign new_n7897 = ~new_n7895 & ~new_n7896 ;
  assign new_n7898 = ~new_n3734 & new_n3737 ;
  assign new_n7899 = new_n3820 & ~new_n4179 ;
  assign new_n7900 = ~new_n3819 & ~new_n7899 ;
  assign new_n7901 = ~new_n7898 & new_n7900 ;
  assign new_n7902 = ~new_n3735 & ~new_n7901 ;
  assign new_n7903 = new_n3735 & new_n7901 ;
  assign new_n7904 = ~new_n7902 & ~new_n7903 ;
  assign new_n7905 = ~new_n3817 & ~new_n7904 ;
  assign new_n7906 = new_n3817 & new_n7902 ;
  assign new_n7907 = new_n4631 & ~new_n7901 ;
  assign new_n7908 = ~new_n7906 & ~new_n7907 ;
  assign new_n7909 = ~new_n7905 & new_n7908 ;
  assign new_n7910 = new_n7403 & ~new_n7909 ;
  assign new_n7911 = ~new_n4904 & ~new_n7407 ;
  assign new_n7912 = new_n4904 & new_n7405 ;
  assign new_n7913 = ~new_n7911 & ~new_n7912 ;
  assign new_n7914 = ~new_n7910 & new_n7913 ;
  assign new_n7915 = ~new_n7392 & ~new_n7914 ;
  assign new_n7916 = new_n7392 & new_n7914 ;
  assign new_n7917 = ~new_n7915 & ~new_n7916 ;
  assign new_n7918 = ~new_n5187 & ~new_n7917 ;
  assign new_n7919 = new_n5187 & new_n7915 ;
  assign new_n7920 = ~new_n6690 & new_n7392 ;
  assign new_n7921 = ~new_n7914 & new_n7920 ;
  assign new_n7922 = ~new_n7919 & ~new_n7921 ;
  assign new_n7923 = ~new_n7918 & new_n7922 ;
  assign new_n7924 = new_n3102 & ~new_n7923 ;
  assign new_n7925 = ~new_n3102 & ~new_n4461 ;
  assign new_n7926 = ~new_n7924 & ~new_n7925 ;
  assign new_n7927 = lo0705 & new_n3186 ;
  assign new_n7928 = lo0704 & new_n3559 ;
  assign new_n7929 = ~new_n3201 & ~new_n7928 ;
  assign new_n7930 = ~new_n7927 & new_n7929 ;
  assign new_n7931 = ~lo0065 & ~new_n7930 ;
  assign new_n7932 = lo0065 & new_n7930 ;
  assign new_n7933 = ~new_n7931 & ~new_n7932 ;
  assign new_n7934 = lo0703 & ~new_n7933 ;
  assign new_n7935 = ~lo0703 & new_n7931 ;
  assign new_n7936 = lo0065 & lo0706 ;
  assign new_n7937 = ~new_n7930 & new_n7936 ;
  assign new_n7938 = ~new_n7935 & ~new_n7937 ;
  assign new_n7939 = ~new_n7934 & new_n7938 ;
  assign new_n7940 = lo0713 & new_n3186 ;
  assign new_n7941 = lo0712 & new_n3559 ;
  assign new_n7942 = ~new_n3201 & ~new_n7941 ;
  assign new_n7943 = ~new_n7940 & new_n7942 ;
  assign new_n7944 = ~lo0065 & ~new_n7943 ;
  assign new_n7945 = lo0065 & new_n7943 ;
  assign new_n7946 = ~new_n7944 & ~new_n7945 ;
  assign new_n7947 = lo0711 & ~new_n7946 ;
  assign new_n7948 = ~lo0711 & new_n7944 ;
  assign new_n7949 = lo0065 & lo0714 ;
  assign new_n7950 = ~new_n7943 & new_n7949 ;
  assign new_n7951 = ~new_n7948 & ~new_n7950 ;
  assign new_n7952 = ~new_n7947 & new_n7951 ;
  assign new_n7953 = new_n3170 & ~new_n7952 ;
  assign new_n7954 = lo0709 & new_n3186 ;
  assign new_n7955 = lo0708 & new_n3202 ;
  assign new_n7956 = ~new_n3201 & ~new_n7955 ;
  assign new_n7957 = ~new_n7954 & new_n7956 ;
  assign new_n7958 = ~lo0063 & ~new_n7957 ;
  assign new_n7959 = lo0063 & new_n7957 ;
  assign new_n7960 = ~new_n7958 & ~new_n7959 ;
  assign new_n7961 = lo0707 & ~new_n7960 ;
  assign new_n7962 = ~lo0707 & new_n7958 ;
  assign new_n7963 = lo0063 & lo0710 ;
  assign new_n7964 = ~new_n7957 & new_n7963 ;
  assign new_n7965 = ~new_n7962 & ~new_n7964 ;
  assign new_n7966 = ~new_n7961 & new_n7965 ;
  assign new_n7967 = new_n3173 & ~new_n7966 ;
  assign new_n7968 = ~new_n3172 & ~new_n7967 ;
  assign new_n7969 = ~new_n7953 & new_n7968 ;
  assign new_n7970 = ~lo0059 & ~new_n7969 ;
  assign new_n7971 = lo0059 & new_n7969 ;
  assign new_n7972 = ~new_n7970 & ~new_n7971 ;
  assign new_n7973 = ~new_n7939 & ~new_n7972 ;
  assign new_n7974 = new_n7939 & new_n7970 ;
  assign new_n7975 = lo0717 & new_n3186 ;
  assign new_n7976 = lo0716 & new_n3202 ;
  assign new_n7977 = ~new_n3201 & ~new_n7976 ;
  assign new_n7978 = ~new_n7975 & new_n7977 ;
  assign new_n7979 = ~lo0063 & ~new_n7978 ;
  assign new_n7980 = lo0063 & new_n7978 ;
  assign new_n7981 = ~new_n7979 & ~new_n7980 ;
  assign new_n7982 = lo0715 & ~new_n7981 ;
  assign new_n7983 = ~lo0715 & new_n7979 ;
  assign new_n7984 = lo0063 & lo0718 ;
  assign new_n7985 = ~new_n7978 & new_n7984 ;
  assign new_n7986 = ~new_n7983 & ~new_n7985 ;
  assign new_n7987 = ~new_n7982 & new_n7986 ;
  assign new_n7988 = lo0059 & ~new_n7987 ;
  assign new_n7989 = ~new_n7969 & new_n7988 ;
  assign new_n7990 = ~new_n7974 & ~new_n7989 ;
  assign new_n7991 = ~new_n7973 & new_n7990 ;
  assign new_n7992 = new_n3169 & ~new_n7991 ;
  assign new_n7993 = ~new_n3160 & ~new_n4446 ;
  assign new_n7994 = lo1398 & new_n3267 ;
  assign new_n7995 = lo1397 & new_n3246 ;
  assign new_n7996 = lo0722 & new_n3258 ;
  assign new_n7997 = ~new_n7995 & ~new_n7996 ;
  assign new_n7998 = ~new_n7994 & new_n7997 ;
  assign new_n7999 = new_n3264 & new_n4450 ;
  assign new_n8000 = lo1352 & new_n3254 ;
  assign new_n8001 = lo1396 & new_n3270 ;
  assign new_n8002 = lo0720 & new_n3274 ;
  assign new_n8003 = ~new_n8001 & ~new_n8002 ;
  assign new_n8004 = ~new_n8000 & new_n8003 ;
  assign new_n8005 = ~new_n7999 & new_n8004 ;
  assign new_n8006 = new_n7998 & new_n8005 ;
  assign new_n8007 = ~new_n7993 & new_n8006 ;
  assign new_n8008 = ~new_n7992 & new_n8007 ;
  assign new_n8009 = new_n3100 & new_n3114 ;
  assign new_n8010 = new_n3125 & new_n8009 ;
  assign new_n8011 = lo0197 & new_n3109 ;
  assign new_n8012 = ~lo0196 & ~new_n8011 ;
  assign new_n8013 = ~lo0198 & lo0199 ;
  assign new_n8014 = lo0200 & new_n8013 ;
  assign new_n8015 = ~new_n3099 & ~new_n8014 ;
  assign new_n8016 = ~new_n8012 & new_n8015 ;
  assign new_n8017 = ~new_n8010 & new_n8016 ;
  assign new_n8018 = ~lo0197 & new_n3100 ;
  assign new_n8019 = ~new_n8009 & new_n8018 ;
  assign new_n8020 = new_n8017 & new_n8019 ;
  assign new_n8021 = new_n4450 & new_n8020 ;
  assign new_n8022 = new_n8009 & ~new_n8017 ;
  assign new_n8023 = lo0713 & new_n8009 ;
  assign new_n8024 = new_n8017 & new_n8023 ;
  assign new_n8025 = ~new_n8022 & ~new_n8024 ;
  assign new_n8026 = ~new_n8021 & new_n8025 ;
  assign new_n8027 = new_n8017 & ~new_n8026 ;
  assign new_n8028 = new_n8008 & new_n8027 ;
  assign new_n8029 = ~new_n8017 & new_n8026 ;
  assign new_n8030 = ~new_n8027 & ~new_n8029 ;
  assign new_n8031 = ~new_n8008 & ~new_n8030 ;
  assign new_n8032 = ~new_n8017 & ~new_n8026 ;
  assign new_n8033 = ~new_n4446 & new_n8032 ;
  assign new_n8034 = ~new_n8031 & ~new_n8033 ;
  assign new_n8035 = ~new_n8028 & new_n8034 ;
  assign new_n8036 = ~new_n3112 & new_n8035 ;
  assign new_n8037 = new_n3112 & ~new_n8035 ;
  assign new_n8038 = ~new_n8036 & ~new_n8037 ;
  assign new_n8039 = new_n3737 & ~new_n4179 ;
  assign new_n8040 = ~new_n4097 & new_n4180 ;
  assign new_n8041 = ~new_n3819 & ~new_n8040 ;
  assign new_n8042 = ~new_n8039 & new_n8041 ;
  assign new_n8043 = new_n3736 & ~new_n8042 ;
  assign new_n8044 = ~new_n3736 & new_n8042 ;
  assign new_n8045 = ~new_n8043 & ~new_n8044 ;
  assign new_n8046 = ~new_n4461 & ~new_n8045 ;
  assign new_n8047 = new_n4461 & new_n8043 ;
  assign new_n8048 = new_n4993 & ~new_n8042 ;
  assign new_n8049 = ~new_n8047 & ~new_n8048 ;
  assign new_n8050 = ~new_n8046 & new_n8049 ;
  assign new_n8051 = new_n7403 & ~new_n8050 ;
  assign new_n8052 = ~new_n5187 & ~new_n7407 ;
  assign new_n8053 = new_n5187 & new_n7405 ;
  assign new_n8054 = ~new_n8052 & ~new_n8053 ;
  assign new_n8055 = ~new_n8051 & new_n8054 ;
  assign new_n8056 = ~new_n7392 & ~new_n8055 ;
  assign new_n8057 = new_n7392 & new_n8055 ;
  assign new_n8058 = ~new_n8056 & ~new_n8057 ;
  assign new_n8059 = ~new_n5472 & ~new_n8058 ;
  assign new_n8060 = new_n5472 & new_n8056 ;
  assign new_n8061 = ~new_n6917 & new_n7392 ;
  assign new_n8062 = ~new_n8055 & new_n8061 ;
  assign new_n8063 = ~new_n8060 & ~new_n8062 ;
  assign new_n8064 = ~new_n8059 & new_n8063 ;
  assign new_n8065 = new_n3102 & ~new_n8064 ;
  assign new_n8066 = ~new_n3102 & ~new_n4904 ;
  assign new_n8067 = ~new_n8065 & ~new_n8066 ;
  assign new_n8068 = lo0685 & new_n3170 ;
  assign new_n8069 = lo0684 & new_n3173 ;
  assign new_n8070 = ~new_n3172 & ~new_n8069 ;
  assign new_n8071 = ~new_n8068 & new_n8070 ;
  assign new_n8072 = ~lo0059 & ~new_n8071 ;
  assign new_n8073 = lo0059 & new_n8071 ;
  assign new_n8074 = ~new_n8072 & ~new_n8073 ;
  assign new_n8075 = lo0683 & ~new_n8074 ;
  assign new_n8076 = ~lo0683 & new_n8072 ;
  assign new_n8077 = lo0059 & lo0686 ;
  assign new_n8078 = ~new_n8071 & new_n8077 ;
  assign new_n8079 = ~new_n8076 & ~new_n8078 ;
  assign new_n8080 = ~new_n8075 & new_n8079 ;
  assign new_n8081 = lo1351 & new_n3170 ;
  assign new_n8082 = lo0692 & new_n3204 ;
  assign new_n8083 = ~new_n3172 & ~new_n8082 ;
  assign new_n8084 = ~new_n8081 & new_n8083 ;
  assign new_n8085 = ~lo0061 & ~new_n8084 ;
  assign new_n8086 = lo0061 & new_n8084 ;
  assign new_n8087 = ~new_n8085 & ~new_n8086 ;
  assign new_n8088 = lo0691 & ~new_n8087 ;
  assign new_n8089 = ~lo0691 & new_n8085 ;
  assign new_n8090 = lo0061 & lo0693 ;
  assign new_n8091 = ~new_n8084 & new_n8090 ;
  assign new_n8092 = ~new_n8089 & ~new_n8091 ;
  assign new_n8093 = ~new_n8088 & new_n8092 ;
  assign new_n8094 = new_n3186 & ~new_n8093 ;
  assign new_n8095 = lo0689 & new_n3170 ;
  assign new_n8096 = lo0688 & new_n3204 ;
  assign new_n8097 = ~new_n3172 & ~new_n8096 ;
  assign new_n8098 = ~new_n8095 & new_n8097 ;
  assign new_n8099 = ~lo0061 & ~new_n8098 ;
  assign new_n8100 = lo0061 & new_n8098 ;
  assign new_n8101 = ~new_n8099 & ~new_n8100 ;
  assign new_n8102 = lo0687 & ~new_n8101 ;
  assign new_n8103 = ~lo0687 & new_n8099 ;
  assign new_n8104 = lo0061 & lo0690 ;
  assign new_n8105 = ~new_n8098 & new_n8104 ;
  assign new_n8106 = ~new_n8103 & ~new_n8105 ;
  assign new_n8107 = ~new_n8102 & new_n8106 ;
  assign new_n8108 = new_n3559 & ~new_n8107 ;
  assign new_n8109 = ~new_n3201 & ~new_n8108 ;
  assign new_n8110 = ~new_n8094 & new_n8109 ;
  assign new_n8111 = ~lo0065 & ~new_n8110 ;
  assign new_n8112 = lo0065 & new_n8110 ;
  assign new_n8113 = ~new_n8111 & ~new_n8112 ;
  assign new_n8114 = ~new_n8080 & ~new_n8113 ;
  assign new_n8115 = new_n8080 & new_n8111 ;
  assign new_n8116 = lo0696 & new_n3170 ;
  assign new_n8117 = lo0695 & new_n3173 ;
  assign new_n8118 = ~new_n3172 & ~new_n8117 ;
  assign new_n8119 = ~new_n8116 & new_n8118 ;
  assign new_n8120 = ~lo0059 & ~new_n8119 ;
  assign new_n8121 = lo0059 & new_n8119 ;
  assign new_n8122 = ~new_n8120 & ~new_n8121 ;
  assign new_n8123 = lo0694 & ~new_n8122 ;
  assign new_n8124 = ~lo0694 & new_n8120 ;
  assign new_n8125 = lo0059 & lo0697 ;
  assign new_n8126 = ~new_n8119 & new_n8125 ;
  assign new_n8127 = ~new_n8124 & ~new_n8126 ;
  assign new_n8128 = ~new_n8123 & new_n8127 ;
  assign new_n8129 = lo0065 & ~new_n8128 ;
  assign new_n8130 = ~new_n8110 & new_n8129 ;
  assign new_n8131 = ~new_n8115 & ~new_n8130 ;
  assign new_n8132 = ~new_n8114 & new_n8131 ;
  assign new_n8133 = new_n3169 & ~new_n8132 ;
  assign new_n8134 = ~new_n3160 & ~new_n4889 ;
  assign new_n8135 = lo1413 & new_n3267 ;
  assign new_n8136 = lo1412 & new_n3246 ;
  assign new_n8137 = lo0702 & new_n3258 ;
  assign new_n8138 = ~new_n8136 & ~new_n8137 ;
  assign new_n8139 = ~new_n8135 & new_n8138 ;
  assign new_n8140 = new_n3264 & new_n4893 ;
  assign new_n8141 = lo0700 & new_n3254 ;
  assign new_n8142 = lo1411 & new_n3270 ;
  assign new_n8143 = lo0699 & new_n3274 ;
  assign new_n8144 = ~new_n8142 & ~new_n8143 ;
  assign new_n8145 = ~new_n8141 & new_n8144 ;
  assign new_n8146 = ~new_n8140 & new_n8145 ;
  assign new_n8147 = new_n8139 & new_n8146 ;
  assign new_n8148 = ~new_n8134 & new_n8147 ;
  assign new_n8149 = ~new_n8133 & new_n8148 ;
  assign new_n8150 = ~new_n8009 & ~new_n8017 ;
  assign new_n8151 = ~new_n8149 & new_n8150 ;
  assign new_n8152 = new_n4893 & new_n8020 ;
  assign new_n8153 = ~new_n8022 & ~new_n8152 ;
  assign new_n8154 = ~new_n8151 & new_n8153 ;
  assign new_n8155 = ~new_n8009 & ~new_n8154 ;
  assign new_n8156 = new_n8009 & new_n8154 ;
  assign new_n8157 = ~new_n8155 & ~new_n8156 ;
  assign new_n8158 = lo1351 & ~new_n8157 ;
  assign new_n8159 = ~lo1351 & new_n8155 ;
  assign new_n8160 = ~new_n4889 & new_n8009 ;
  assign new_n8161 = ~new_n8154 & new_n8160 ;
  assign new_n8162 = ~new_n8159 & ~new_n8161 ;
  assign new_n8163 = ~new_n8158 & new_n8162 ;
  assign new_n8164 = ~new_n3112 & new_n8163 ;
  assign new_n8165 = new_n3112 & ~new_n8163 ;
  assign new_n8166 = ~new_n8164 & ~new_n8165 ;
  assign new_n8167 = new_n3737 & ~new_n4461 ;
  assign new_n8168 = new_n3820 & ~new_n4904 ;
  assign new_n8169 = ~new_n3819 & ~new_n8168 ;
  assign new_n8170 = ~new_n8167 & new_n8169 ;
  assign new_n8171 = ~new_n3735 & ~new_n8170 ;
  assign new_n8172 = new_n3735 & new_n8170 ;
  assign new_n8173 = ~new_n8171 & ~new_n8172 ;
  assign new_n8174 = ~new_n4541 & ~new_n8173 ;
  assign new_n8175 = new_n4541 & new_n8171 ;
  assign new_n8176 = new_n5277 & ~new_n8170 ;
  assign new_n8177 = ~new_n8175 & ~new_n8176 ;
  assign new_n8178 = ~new_n8174 & new_n8177 ;
  assign new_n8179 = new_n7403 & ~new_n8178 ;
  assign new_n8180 = ~new_n5472 & ~new_n7407 ;
  assign new_n8181 = new_n5472 & new_n7405 ;
  assign new_n8182 = ~new_n8180 & ~new_n8181 ;
  assign new_n8183 = ~new_n8179 & new_n8182 ;
  assign new_n8184 = ~new_n7392 & ~new_n8183 ;
  assign new_n8185 = new_n7392 & new_n8183 ;
  assign new_n8186 = ~new_n8184 & ~new_n8185 ;
  assign new_n8187 = ~new_n5766 & ~new_n8186 ;
  assign new_n8188 = new_n5766 & new_n8184 ;
  assign new_n8189 = ~new_n7138 & new_n7392 ;
  assign new_n8190 = ~new_n8183 & new_n8189 ;
  assign new_n8191 = ~new_n8188 & ~new_n8190 ;
  assign new_n8192 = ~new_n8187 & new_n8191 ;
  assign new_n8193 = new_n3102 & ~new_n8192 ;
  assign new_n8194 = ~new_n3102 & ~new_n5187 ;
  assign new_n8195 = ~new_n8193 & ~new_n8194 ;
  assign new_n8196 = lo0808 & new_n3186 ;
  assign new_n8197 = lo0807 & new_n3559 ;
  assign new_n8198 = ~new_n3201 & ~new_n8197 ;
  assign new_n8199 = ~new_n8196 & new_n8198 ;
  assign new_n8200 = ~lo0065 & ~new_n8199 ;
  assign new_n8201 = lo0065 & new_n8199 ;
  assign new_n8202 = ~new_n8200 & ~new_n8201 ;
  assign new_n8203 = lo0806 & ~new_n8202 ;
  assign new_n8204 = ~lo0806 & new_n8200 ;
  assign new_n8205 = lo0065 & lo0809 ;
  assign new_n8206 = ~new_n8199 & new_n8205 ;
  assign new_n8207 = ~new_n8204 & ~new_n8206 ;
  assign new_n8208 = ~new_n8203 & new_n8207 ;
  assign new_n8209 = lo0816 & new_n3186 ;
  assign new_n8210 = lo0815 & new_n3202 ;
  assign new_n8211 = ~new_n3201 & ~new_n8210 ;
  assign new_n8212 = ~new_n8209 & new_n8211 ;
  assign new_n8213 = ~lo0063 & ~new_n8212 ;
  assign new_n8214 = lo0063 & new_n8212 ;
  assign new_n8215 = ~new_n8213 & ~new_n8214 ;
  assign new_n8216 = lo0814 & ~new_n8215 ;
  assign new_n8217 = ~lo0814 & new_n8213 ;
  assign new_n8218 = lo0063 & lo0817 ;
  assign new_n8219 = ~new_n8212 & new_n8218 ;
  assign new_n8220 = ~new_n8217 & ~new_n8219 ;
  assign new_n8221 = ~new_n8216 & new_n8220 ;
  assign new_n8222 = new_n3170 & ~new_n8221 ;
  assign new_n8223 = lo0812 & new_n3186 ;
  assign new_n8224 = lo0811 & new_n3202 ;
  assign new_n8225 = ~new_n3201 & ~new_n8224 ;
  assign new_n8226 = ~new_n8223 & new_n8225 ;
  assign new_n8227 = ~lo0063 & ~new_n8226 ;
  assign new_n8228 = lo0063 & new_n8226 ;
  assign new_n8229 = ~new_n8227 & ~new_n8228 ;
  assign new_n8230 = lo0810 & ~new_n8229 ;
  assign new_n8231 = ~lo0810 & new_n8227 ;
  assign new_n8232 = lo0063 & lo0813 ;
  assign new_n8233 = ~new_n8226 & new_n8232 ;
  assign new_n8234 = ~new_n8231 & ~new_n8233 ;
  assign new_n8235 = ~new_n8230 & new_n8234 ;
  assign new_n8236 = new_n3204 & ~new_n8235 ;
  assign new_n8237 = ~new_n3172 & ~new_n8236 ;
  assign new_n8238 = ~new_n8222 & new_n8237 ;
  assign new_n8239 = ~lo0061 & ~new_n8238 ;
  assign new_n8240 = lo0061 & new_n8238 ;
  assign new_n8241 = ~new_n8239 & ~new_n8240 ;
  assign new_n8242 = ~new_n8208 & ~new_n8241 ;
  assign new_n8243 = new_n8208 & new_n8239 ;
  assign new_n8244 = lo0820 & new_n3186 ;
  assign new_n8245 = lo0819 & new_n3559 ;
  assign new_n8246 = ~new_n3201 & ~new_n8245 ;
  assign new_n8247 = ~new_n8244 & new_n8246 ;
  assign new_n8248 = ~lo0065 & ~new_n8247 ;
  assign new_n8249 = lo0065 & new_n8247 ;
  assign new_n8250 = ~new_n8248 & ~new_n8249 ;
  assign new_n8251 = lo0818 & ~new_n8250 ;
  assign new_n8252 = ~lo0818 & new_n8248 ;
  assign new_n8253 = lo0065 & lo0821 ;
  assign new_n8254 = ~new_n8247 & new_n8253 ;
  assign new_n8255 = ~new_n8252 & ~new_n8254 ;
  assign new_n8256 = ~new_n8251 & new_n8255 ;
  assign new_n8257 = lo0061 & ~new_n8256 ;
  assign new_n8258 = ~new_n8238 & new_n8257 ;
  assign new_n8259 = ~new_n8243 & ~new_n8258 ;
  assign new_n8260 = ~new_n8242 & new_n8259 ;
  assign new_n8261 = new_n3169 & ~new_n8260 ;
  assign new_n8262 = ~new_n3160 & ~new_n5170 ;
  assign new_n8263 = lo0070 & ~lo0071 ;
  assign new_n8264 = new_n3256 & new_n8263 ;
  assign new_n8265 = lo0826 & new_n8264 ;
  assign new_n8266 = lo0824 & new_n3258 ;
  assign new_n8267 = lo1387 & new_n3267 ;
  assign new_n8268 = ~new_n8266 & ~new_n8267 ;
  assign new_n8269 = ~new_n8265 & new_n8268 ;
  assign new_n8270 = lo1388 & new_n3246 ;
  assign new_n8271 = lo1386 & new_n3270 ;
  assign new_n8272 = lo0825 & new_n3274 ;
  assign new_n8273 = ~new_n8271 & ~new_n8272 ;
  assign new_n8274 = ~new_n8270 & new_n8273 ;
  assign new_n8275 = new_n3264 & new_n5176 ;
  assign new_n8276 = lo1381 & new_n3254 ;
  assign new_n8277 = ~new_n8275 & ~new_n8276 ;
  assign new_n8278 = new_n8274 & new_n8277 ;
  assign new_n8279 = new_n8269 & new_n8278 ;
  assign new_n8280 = ~new_n8262 & new_n8279 ;
  assign new_n8281 = ~new_n8261 & new_n8280 ;
  assign new_n8282 = new_n5176 & new_n8020 ;
  assign new_n8283 = lo0816 & new_n8009 ;
  assign new_n8284 = new_n8017 & new_n8283 ;
  assign new_n8285 = ~new_n8022 & ~new_n8284 ;
  assign new_n8286 = ~new_n8282 & new_n8285 ;
  assign new_n8287 = new_n8017 & ~new_n8286 ;
  assign new_n8288 = new_n8281 & new_n8287 ;
  assign new_n8289 = ~new_n8017 & new_n8286 ;
  assign new_n8290 = ~new_n8287 & ~new_n8289 ;
  assign new_n8291 = ~new_n8281 & ~new_n8290 ;
  assign new_n8292 = ~new_n8017 & ~new_n8286 ;
  assign new_n8293 = ~new_n5170 & new_n8292 ;
  assign new_n8294 = ~new_n8291 & ~new_n8293 ;
  assign new_n8295 = ~new_n8288 & new_n8294 ;
  assign new_n8296 = ~new_n3112 & new_n8295 ;
  assign new_n8297 = new_n3112 & ~new_n8295 ;
  assign new_n8298 = ~new_n8296 & ~new_n8297 ;
  assign new_n8299 = new_n3737 & ~new_n4904 ;
  assign new_n8300 = new_n4180 & ~new_n4818 ;
  assign new_n8301 = ~new_n3819 & ~new_n8300 ;
  assign new_n8302 = ~new_n8299 & new_n8301 ;
  assign new_n8303 = new_n3736 & ~new_n8302 ;
  assign new_n8304 = ~new_n3736 & new_n8302 ;
  assign new_n8305 = ~new_n8303 & ~new_n8304 ;
  assign new_n8306 = ~new_n5187 & ~new_n8305 ;
  assign new_n8307 = new_n5187 & new_n8303 ;
  assign new_n8308 = new_n5561 & ~new_n8302 ;
  assign new_n8309 = ~new_n8307 & ~new_n8308 ;
  assign new_n8310 = ~new_n8306 & new_n8309 ;
  assign new_n8311 = new_n7403 & ~new_n8310 ;
  assign new_n8312 = ~new_n5766 & ~new_n7407 ;
  assign new_n8313 = new_n5766 & new_n7405 ;
  assign new_n8314 = ~new_n8312 & ~new_n8313 ;
  assign new_n8315 = ~new_n8311 & new_n8314 ;
  assign new_n8316 = ~new_n7392 & ~new_n8315 ;
  assign new_n8317 = new_n7392 & new_n8315 ;
  assign new_n8318 = ~new_n8316 & ~new_n8317 ;
  assign new_n8319 = ~new_n5996 & ~new_n8318 ;
  assign new_n8320 = new_n5996 & new_n8316 ;
  assign new_n8321 = ~new_n2619 & new_n7392 ;
  assign new_n8322 = ~new_n8315 & new_n8321 ;
  assign new_n8323 = ~new_n8320 & ~new_n8322 ;
  assign new_n8324 = ~new_n8319 & new_n8323 ;
  assign new_n8325 = new_n3102 & ~new_n8324 ;
  assign new_n8326 = ~new_n3102 & ~new_n5472 ;
  assign new_n8327 = ~new_n8325 & ~new_n8326 ;
  assign new_n8328 = lo0076 & new_n3170 ;
  assign new_n8329 = lo0075 & new_n3173 ;
  assign new_n8330 = ~new_n3172 & ~new_n8329 ;
  assign new_n8331 = ~new_n8328 & new_n8330 ;
  assign new_n8332 = ~lo0059 & ~new_n8331 ;
  assign new_n8333 = lo0059 & new_n8331 ;
  assign new_n8334 = ~new_n8332 & ~new_n8333 ;
  assign new_n8335 = lo0074 & ~new_n8334 ;
  assign new_n8336 = ~lo0074 & new_n8332 ;
  assign new_n8337 = lo0059 & lo0077 ;
  assign new_n8338 = ~new_n8331 & new_n8337 ;
  assign new_n8339 = ~new_n8336 & ~new_n8338 ;
  assign new_n8340 = ~new_n8335 & new_n8339 ;
  assign new_n8341 = lo0084 & new_n3170 ;
  assign new_n8342 = lo0083 & new_n3173 ;
  assign new_n8343 = ~new_n3172 & ~new_n8342 ;
  assign new_n8344 = ~new_n8341 & new_n8343 ;
  assign new_n8345 = ~lo0059 & ~new_n8344 ;
  assign new_n8346 = lo0059 & new_n8344 ;
  assign new_n8347 = ~new_n8345 & ~new_n8346 ;
  assign new_n8348 = lo0082 & ~new_n8347 ;
  assign new_n8349 = ~lo0082 & new_n8345 ;
  assign new_n8350 = lo0059 & lo0085 ;
  assign new_n8351 = ~new_n8344 & new_n8350 ;
  assign new_n8352 = ~new_n8349 & ~new_n8351 ;
  assign new_n8353 = ~new_n8348 & new_n8352 ;
  assign new_n8354 = new_n3186 & ~new_n8353 ;
  assign new_n8355 = lo0080 & new_n3170 ;
  assign new_n8356 = lo0079 & new_n3204 ;
  assign new_n8357 = ~new_n3172 & ~new_n8356 ;
  assign new_n8358 = ~new_n8355 & new_n8357 ;
  assign new_n8359 = ~lo0061 & ~new_n8358 ;
  assign new_n8360 = lo0061 & new_n8358 ;
  assign new_n8361 = ~new_n8359 & ~new_n8360 ;
  assign new_n8362 = lo0078 & ~new_n8361 ;
  assign new_n8363 = ~lo0078 & new_n8359 ;
  assign new_n8364 = lo0061 & lo0081 ;
  assign new_n8365 = ~new_n8358 & new_n8364 ;
  assign new_n8366 = ~new_n8363 & ~new_n8365 ;
  assign new_n8367 = ~new_n8362 & new_n8366 ;
  assign new_n8368 = new_n3202 & ~new_n8367 ;
  assign new_n8369 = ~new_n3201 & ~new_n8368 ;
  assign new_n8370 = ~new_n8354 & new_n8369 ;
  assign new_n8371 = ~lo0063 & ~new_n8370 ;
  assign new_n8372 = lo0063 & new_n8370 ;
  assign new_n8373 = ~new_n8371 & ~new_n8372 ;
  assign new_n8374 = ~new_n8340 & ~new_n8373 ;
  assign new_n8375 = new_n8340 & new_n8371 ;
  assign new_n8376 = lo0088 & new_n3170 ;
  assign new_n8377 = lo0087 & new_n3204 ;
  assign new_n8378 = ~new_n3172 & ~new_n8377 ;
  assign new_n8379 = ~new_n8376 & new_n8378 ;
  assign new_n8380 = ~lo0061 & ~new_n8379 ;
  assign new_n8381 = lo0061 & new_n8379 ;
  assign new_n8382 = ~new_n8380 & ~new_n8381 ;
  assign new_n8383 = lo0086 & ~new_n8382 ;
  assign new_n8384 = ~lo0086 & new_n8380 ;
  assign new_n8385 = lo0061 & lo0089 ;
  assign new_n8386 = ~new_n8379 & new_n8385 ;
  assign new_n8387 = ~new_n8384 & ~new_n8386 ;
  assign new_n8388 = ~new_n8383 & new_n8387 ;
  assign new_n8389 = lo0063 & ~new_n8388 ;
  assign new_n8390 = ~new_n8370 & new_n8389 ;
  assign new_n8391 = ~new_n8375 & ~new_n8390 ;
  assign new_n8392 = ~new_n8374 & new_n8391 ;
  assign new_n8393 = new_n3169 & ~new_n8392 ;
  assign new_n8394 = ~new_n3160 & ~new_n5455 ;
  assign new_n8395 = lo1288 & new_n3254 ;
  assign new_n8396 = lo1286 & new_n3246 ;
  assign new_n8397 = lo0110 & new_n8264 ;
  assign new_n8398 = ~new_n8396 & ~new_n8397 ;
  assign new_n8399 = ~new_n8395 & new_n8398 ;
  assign new_n8400 = new_n3264 & new_n5465 ;
  assign new_n8401 = lo1287 & new_n3270 ;
  assign new_n8402 = lo0111 & new_n3274 ;
  assign new_n8403 = ~new_n8401 & ~new_n8402 ;
  assign new_n8404 = ~new_n8400 & new_n8403 ;
  assign new_n8405 = lo0109 & new_n3258 ;
  assign new_n8406 = lo1289 & new_n3267 ;
  assign new_n8407 = ~new_n8405 & ~new_n8406 ;
  assign new_n8408 = new_n8404 & new_n8407 ;
  assign new_n8409 = new_n8399 & new_n8408 ;
  assign new_n8410 = ~new_n8394 & new_n8409 ;
  assign new_n8411 = ~new_n8393 & new_n8410 ;
  assign new_n8412 = new_n8150 & ~new_n8411 ;
  assign new_n8413 = new_n5465 & new_n8019 ;
  assign new_n8414 = new_n8017 & new_n8413 ;
  assign new_n8415 = ~new_n8022 & ~new_n8414 ;
  assign new_n8416 = ~new_n8412 & new_n8415 ;
  assign new_n8417 = ~new_n8009 & ~new_n8416 ;
  assign new_n8418 = new_n8009 & new_n8416 ;
  assign new_n8419 = ~new_n8417 & ~new_n8418 ;
  assign new_n8420 = lo0084 & ~new_n8419 ;
  assign new_n8421 = ~lo0084 & new_n8417 ;
  assign new_n8422 = ~new_n5455 & new_n8009 ;
  assign new_n8423 = ~new_n8416 & new_n8422 ;
  assign new_n8424 = ~new_n8421 & ~new_n8423 ;
  assign new_n8425 = ~new_n8420 & new_n8424 ;
  assign new_n8426 = ~new_n3112 & new_n8425 ;
  assign new_n8427 = new_n3112 & ~new_n8425 ;
  assign new_n8428 = ~new_n8426 & ~new_n8427 ;
  assign new_n8429 = new_n3737 & ~new_n5187 ;
  assign new_n8430 = new_n3820 & ~new_n5472 ;
  assign new_n8431 = ~new_n3819 & ~new_n8430 ;
  assign new_n8432 = ~new_n8429 & new_n8431 ;
  assign new_n8433 = ~new_n3735 & ~new_n8432 ;
  assign new_n8434 = new_n3735 & new_n8432 ;
  assign new_n8435 = ~new_n8433 & ~new_n8434 ;
  assign new_n8436 = ~new_n2824 & ~new_n8435 ;
  assign new_n8437 = new_n2824 & new_n8433 ;
  assign new_n8438 = new_n5776 & ~new_n8432 ;
  assign new_n8439 = ~new_n8437 & ~new_n8438 ;
  assign new_n8440 = ~new_n8436 & new_n8439 ;
  assign new_n8441 = lo0298 & ~new_n8440 ;
  assign new_n8442 = new_n3914 & ~new_n6225 ;
  assign new_n8443 = ~lo0297 & ~new_n5996 ;
  assign new_n8444 = ~new_n8442 & ~new_n8443 ;
  assign new_n8445 = ~lo0298 & ~new_n8444 ;
  assign new_n8446 = ~new_n8441 & ~new_n8445 ;
  assign new_n8447 = new_n3102 & ~new_n8446 ;
  assign new_n8448 = ~new_n3102 & ~new_n5766 ;
  assign new_n8449 = ~new_n8447 & ~new_n8448 ;
  assign new_n8450 = lo0384 & new_n3186 ;
  assign new_n8451 = lo0383 & new_n3559 ;
  assign new_n8452 = ~new_n3201 & ~new_n8451 ;
  assign new_n8453 = ~new_n8450 & new_n8452 ;
  assign new_n8454 = ~lo0065 & ~new_n8453 ;
  assign new_n8455 = lo0065 & new_n8453 ;
  assign new_n8456 = ~new_n8454 & ~new_n8455 ;
  assign new_n8457 = lo0382 & ~new_n8456 ;
  assign new_n8458 = ~lo0382 & new_n8454 ;
  assign new_n8459 = lo0065 & lo0385 ;
  assign new_n8460 = ~new_n8453 & new_n8459 ;
  assign new_n8461 = ~new_n8458 & ~new_n8460 ;
  assign new_n8462 = ~new_n8457 & new_n8461 ;
  assign new_n8463 = lo0392 & new_n3186 ;
  assign new_n8464 = lo0391 & new_n3559 ;
  assign new_n8465 = ~new_n3201 & ~new_n8464 ;
  assign new_n8466 = ~new_n8463 & new_n8465 ;
  assign new_n8467 = ~lo0065 & ~new_n8466 ;
  assign new_n8468 = lo0065 & new_n8466 ;
  assign new_n8469 = ~new_n8467 & ~new_n8468 ;
  assign new_n8470 = lo0390 & ~new_n8469 ;
  assign new_n8471 = ~lo0390 & new_n8467 ;
  assign new_n8472 = lo0065 & lo0393 ;
  assign new_n8473 = ~new_n8466 & new_n8472 ;
  assign new_n8474 = ~new_n8471 & ~new_n8473 ;
  assign new_n8475 = ~new_n8470 & new_n8474 ;
  assign new_n8476 = new_n3170 & ~new_n8475 ;
  assign new_n8477 = lo0388 & new_n3186 ;
  assign new_n8478 = lo0387 & new_n3202 ;
  assign new_n8479 = ~new_n3201 & ~new_n8478 ;
  assign new_n8480 = ~new_n8477 & new_n8479 ;
  assign new_n8481 = ~lo0063 & ~new_n8480 ;
  assign new_n8482 = lo0063 & new_n8480 ;
  assign new_n8483 = ~new_n8481 & ~new_n8482 ;
  assign new_n8484 = lo0386 & ~new_n8483 ;
  assign new_n8485 = ~lo0386 & new_n8481 ;
  assign new_n8486 = lo0063 & lo0389 ;
  assign new_n8487 = ~new_n8480 & new_n8486 ;
  assign new_n8488 = ~new_n8485 & ~new_n8487 ;
  assign new_n8489 = ~new_n8484 & new_n8488 ;
  assign new_n8490 = new_n3173 & ~new_n8489 ;
  assign new_n8491 = ~new_n3172 & ~new_n8490 ;
  assign new_n8492 = ~new_n8476 & new_n8491 ;
  assign new_n8493 = ~lo0059 & ~new_n8492 ;
  assign new_n8494 = lo0059 & new_n8492 ;
  assign new_n8495 = ~new_n8493 & ~new_n8494 ;
  assign new_n8496 = ~new_n8462 & ~new_n8495 ;
  assign new_n8497 = new_n8462 & new_n8493 ;
  assign new_n8498 = lo0396 & new_n3186 ;
  assign new_n8499 = lo0395 & new_n3202 ;
  assign new_n8500 = ~new_n3201 & ~new_n8499 ;
  assign new_n8501 = ~new_n8498 & new_n8500 ;
  assign new_n8502 = ~lo0063 & ~new_n8501 ;
  assign new_n8503 = lo0063 & new_n8501 ;
  assign new_n8504 = ~new_n8502 & ~new_n8503 ;
  assign new_n8505 = lo0394 & ~new_n8504 ;
  assign new_n8506 = ~lo0394 & new_n8502 ;
  assign new_n8507 = lo0063 & lo0397 ;
  assign new_n8508 = ~new_n8501 & new_n8507 ;
  assign new_n8509 = ~new_n8506 & ~new_n8508 ;
  assign new_n8510 = ~new_n8505 & new_n8509 ;
  assign new_n8511 = lo0059 & ~new_n8510 ;
  assign new_n8512 = ~new_n8492 & new_n8511 ;
  assign new_n8513 = ~new_n8497 & ~new_n8512 ;
  assign new_n8514 = ~new_n8496 & new_n8513 ;
  assign new_n8515 = new_n3169 & ~new_n8514 ;
  assign new_n8516 = ~new_n3160 & ~new_n5743 ;
  assign new_n8517 = new_n3264 & new_n5755 ;
  assign new_n8518 = lo1311 & new_n3267 ;
  assign new_n8519 = lo1310 & new_n3270 ;
  assign new_n8520 = lo0399 & new_n3274 ;
  assign new_n8521 = ~new_n8519 & ~new_n8520 ;
  assign new_n8522 = ~new_n8518 & new_n8521 ;
  assign new_n8523 = lo0181 & new_n8264 ;
  assign new_n8524 = lo0400 & new_n3258 ;
  assign new_n8525 = ~new_n8523 & ~new_n8524 ;
  assign new_n8526 = lo1309 & new_n3254 ;
  assign new_n8527 = lo1312 & new_n3246 ;
  assign new_n8528 = ~new_n8526 & ~new_n8527 ;
  assign new_n8529 = new_n8525 & new_n8528 ;
  assign new_n8530 = new_n8522 & new_n8529 ;
  assign new_n8531 = ~new_n8517 & new_n8530 ;
  assign new_n8532 = ~new_n8516 & new_n8531 ;
  assign new_n8533 = ~new_n8515 & new_n8532 ;
  assign new_n8534 = ~lo0200 & ~new_n5755 ;
  assign new_n8535 = ~lo0197 & lo0199 ;
  assign new_n8536 = ~new_n8009 & new_n8535 ;
  assign new_n8537 = new_n8017 & new_n8536 ;
  assign new_n8538 = ~new_n8534 & new_n8537 ;
  assign new_n8539 = lo0392 & new_n8009 ;
  assign new_n8540 = new_n8017 & new_n8539 ;
  assign new_n8541 = ~new_n8022 & ~new_n8540 ;
  assign new_n8542 = ~new_n8538 & new_n8541 ;
  assign new_n8543 = new_n8017 & ~new_n8542 ;
  assign new_n8544 = new_n8533 & new_n8543 ;
  assign new_n8545 = ~new_n8017 & new_n8542 ;
  assign new_n8546 = ~new_n8543 & ~new_n8545 ;
  assign new_n8547 = ~new_n8533 & ~new_n8546 ;
  assign new_n8548 = ~new_n8017 & ~new_n8542 ;
  assign new_n8549 = ~new_n5743 & new_n8548 ;
  assign new_n8550 = ~new_n8547 & ~new_n8549 ;
  assign new_n8551 = ~new_n8544 & new_n8550 ;
  assign new_n8552 = ~new_n3112 & new_n8551 ;
  assign new_n8553 = new_n3112 & ~new_n8551 ;
  assign new_n8554 = ~new_n8552 & ~new_n8553 ;
  assign new_n8555 = new_n3737 & ~new_n5472 ;
  assign new_n8556 = ~new_n3549 & new_n4180 ;
  assign new_n8557 = ~new_n3819 & ~new_n8556 ;
  assign new_n8558 = ~new_n8555 & new_n8557 ;
  assign new_n8559 = new_n3736 & ~new_n8558 ;
  assign new_n8560 = ~new_n3736 & new_n8558 ;
  assign new_n8561 = ~new_n8559 & ~new_n8560 ;
  assign new_n8562 = ~new_n5766 & ~new_n8561 ;
  assign new_n8563 = new_n5766 & new_n8559 ;
  assign new_n8564 = new_n6005 & ~new_n8558 ;
  assign new_n8565 = ~new_n8563 & ~new_n8564 ;
  assign new_n8566 = ~new_n8562 & new_n8565 ;
  assign new_n8567 = lo0298 & ~new_n8566 ;
  assign new_n8568 = new_n3914 & ~new_n6461 ;
  assign new_n8569 = ~lo0297 & ~new_n6225 ;
  assign new_n8570 = ~new_n8568 & ~new_n8569 ;
  assign new_n8571 = ~lo0298 & ~new_n8570 ;
  assign new_n8572 = ~new_n8567 & ~new_n8571 ;
  assign new_n8573 = new_n3102 & ~new_n8572 ;
  assign new_n8574 = ~new_n3102 & ~new_n5996 ;
  assign new_n8575 = ~new_n8573 & ~new_n8574 ;
  assign new_n8576 = lo0501 & new_n3170 ;
  assign new_n8577 = lo0500 & new_n3173 ;
  assign new_n8578 = ~new_n3172 & ~new_n8577 ;
  assign new_n8579 = ~new_n8576 & new_n8578 ;
  assign new_n8580 = ~lo0059 & ~new_n8579 ;
  assign new_n8581 = lo0059 & new_n8579 ;
  assign new_n8582 = ~new_n8580 & ~new_n8581 ;
  assign new_n8583 = lo0499 & ~new_n8582 ;
  assign new_n8584 = ~lo0499 & new_n8580 ;
  assign new_n8585 = lo0059 & lo0502 ;
  assign new_n8586 = ~new_n8579 & new_n8585 ;
  assign new_n8587 = ~new_n8584 & ~new_n8586 ;
  assign new_n8588 = ~new_n8583 & new_n8587 ;
  assign new_n8589 = lo0498 & new_n3170 ;
  assign new_n8590 = lo0508 & new_n3204 ;
  assign new_n8591 = ~new_n3172 & ~new_n8590 ;
  assign new_n8592 = ~new_n8589 & new_n8591 ;
  assign new_n8593 = ~lo0061 & ~new_n8592 ;
  assign new_n8594 = lo0061 & new_n8592 ;
  assign new_n8595 = ~new_n8593 & ~new_n8594 ;
  assign new_n8596 = lo0507 & ~new_n8595 ;
  assign new_n8597 = ~lo0507 & new_n8593 ;
  assign new_n8598 = lo0061 & lo0509 ;
  assign new_n8599 = ~new_n8592 & new_n8598 ;
  assign new_n8600 = ~new_n8597 & ~new_n8599 ;
  assign new_n8601 = ~new_n8596 & new_n8600 ;
  assign new_n8602 = new_n3186 & ~new_n8601 ;
  assign new_n8603 = lo0505 & new_n3170 ;
  assign new_n8604 = lo0504 & new_n3204 ;
  assign new_n8605 = ~new_n3172 & ~new_n8604 ;
  assign new_n8606 = ~new_n8603 & new_n8605 ;
  assign new_n8607 = ~lo0061 & ~new_n8606 ;
  assign new_n8608 = lo0061 & new_n8606 ;
  assign new_n8609 = ~new_n8607 & ~new_n8608 ;
  assign new_n8610 = lo0503 & ~new_n8609 ;
  assign new_n8611 = ~lo0503 & new_n8607 ;
  assign new_n8612 = lo0061 & lo0506 ;
  assign new_n8613 = ~new_n8606 & new_n8612 ;
  assign new_n8614 = ~new_n8611 & ~new_n8613 ;
  assign new_n8615 = ~new_n8610 & new_n8614 ;
  assign new_n8616 = new_n3559 & ~new_n8615 ;
  assign new_n8617 = ~new_n3201 & ~new_n8616 ;
  assign new_n8618 = ~new_n8602 & new_n8617 ;
  assign new_n8619 = ~lo0065 & ~new_n8618 ;
  assign new_n8620 = lo0065 & new_n8618 ;
  assign new_n8621 = ~new_n8619 & ~new_n8620 ;
  assign new_n8622 = ~new_n8588 & ~new_n8621 ;
  assign new_n8623 = new_n8588 & new_n8619 ;
  assign new_n8624 = lo0512 & new_n3170 ;
  assign new_n8625 = lo0511 & new_n3173 ;
  assign new_n8626 = ~new_n3172 & ~new_n8625 ;
  assign new_n8627 = ~new_n8624 & new_n8626 ;
  assign new_n8628 = ~lo0059 & ~new_n8627 ;
  assign new_n8629 = lo0059 & new_n8627 ;
  assign new_n8630 = ~new_n8628 & ~new_n8629 ;
  assign new_n8631 = lo0510 & ~new_n8630 ;
  assign new_n8632 = ~lo0510 & new_n8628 ;
  assign new_n8633 = lo0059 & lo0513 ;
  assign new_n8634 = ~new_n8627 & new_n8633 ;
  assign new_n8635 = ~new_n8632 & ~new_n8634 ;
  assign new_n8636 = ~new_n8631 & new_n8635 ;
  assign new_n8637 = lo0065 & ~new_n8636 ;
  assign new_n8638 = ~new_n8618 & new_n8637 ;
  assign new_n8639 = ~new_n8623 & ~new_n8638 ;
  assign new_n8640 = ~new_n8622 & new_n8639 ;
  assign new_n8641 = new_n3169 & ~new_n8640 ;
  assign new_n8642 = ~new_n3160 & new_n5977 ;
  assign new_n8643 = new_n3264 & new_n5985 ;
  assign new_n8644 = lo1324 & new_n3246 ;
  assign new_n8645 = lo1321 & new_n3270 ;
  assign new_n8646 = lo0516 & new_n3274 ;
  assign new_n8647 = ~new_n8645 & ~new_n8646 ;
  assign new_n8648 = ~new_n8644 & new_n8647 ;
  assign new_n8649 = lo0515 & new_n3258 ;
  assign new_n8650 = lo1323 & new_n3267 ;
  assign new_n8651 = ~new_n8649 & ~new_n8650 ;
  assign new_n8652 = lo1322 & new_n3254 ;
  assign new_n8653 = lo0183 & new_n8264 ;
  assign new_n8654 = ~new_n8652 & ~new_n8653 ;
  assign new_n8655 = new_n8651 & new_n8654 ;
  assign new_n8656 = new_n8648 & new_n8655 ;
  assign new_n8657 = ~new_n8643 & new_n8656 ;
  assign new_n8658 = ~new_n8642 & new_n8657 ;
  assign new_n8659 = ~new_n8641 & new_n8658 ;
  assign new_n8660 = new_n8150 & ~new_n8659 ;
  assign new_n8661 = new_n5985 & new_n8020 ;
  assign new_n8662 = ~new_n8022 & ~new_n8661 ;
  assign new_n8663 = ~new_n8660 & new_n8662 ;
  assign new_n8664 = ~new_n8009 & ~new_n8663 ;
  assign new_n8665 = new_n8009 & new_n8663 ;
  assign new_n8666 = ~new_n8664 & ~new_n8665 ;
  assign new_n8667 = lo0498 & ~new_n8666 ;
  assign new_n8668 = ~lo0498 & new_n8664 ;
  assign new_n8669 = new_n5977 & new_n8009 ;
  assign new_n8670 = ~new_n8663 & new_n8669 ;
  assign new_n8671 = ~new_n8668 & ~new_n8670 ;
  assign new_n8672 = ~new_n8667 & new_n8671 ;
  assign new_n8673 = ~new_n3112 & new_n8672 ;
  assign new_n8674 = new_n3112 & ~new_n8672 ;
  assign new_n8675 = ~new_n8673 & ~new_n8674 ;
  assign new_n8676 = new_n3737 & ~new_n5766 ;
  assign new_n8677 = new_n3820 & ~new_n5996 ;
  assign new_n8678 = ~new_n3819 & ~new_n8677 ;
  assign new_n8679 = ~new_n8676 & new_n8678 ;
  assign new_n8680 = ~new_n3735 & ~new_n8679 ;
  assign new_n8681 = new_n3735 & new_n8679 ;
  assign new_n8682 = ~new_n8680 & ~new_n8681 ;
  assign new_n8683 = ~new_n3908 & ~new_n8682 ;
  assign new_n8684 = new_n3908 & new_n8680 ;
  assign new_n8685 = new_n6235 & ~new_n8679 ;
  assign new_n8686 = ~new_n8684 & ~new_n8685 ;
  assign new_n8687 = ~new_n8683 & new_n8686 ;
  assign new_n8688 = lo0298 & ~new_n8687 ;
  assign new_n8689 = new_n3914 & ~new_n6690 ;
  assign new_n8690 = ~lo0297 & ~new_n6461 ;
  assign new_n8691 = ~new_n8689 & ~new_n8690 ;
  assign new_n8692 = ~lo0298 & ~new_n8691 ;
  assign new_n8693 = ~new_n8688 & ~new_n8692 ;
  assign new_n8694 = new_n3102 & ~new_n8693 ;
  assign new_n8695 = ~new_n3102 & ~new_n6225 ;
  assign new_n8696 = ~new_n8694 & ~new_n8695 ;
  assign new_n8697 = lo0585 & new_n3186 ;
  assign new_n8698 = lo0584 & new_n3559 ;
  assign new_n8699 = ~new_n3201 & ~new_n8698 ;
  assign new_n8700 = ~new_n8697 & new_n8699 ;
  assign new_n8701 = ~lo0065 & ~new_n8700 ;
  assign new_n8702 = lo0065 & new_n8700 ;
  assign new_n8703 = ~new_n8701 & ~new_n8702 ;
  assign new_n8704 = lo0583 & ~new_n8703 ;
  assign new_n8705 = ~lo0583 & new_n8701 ;
  assign new_n8706 = lo0065 & lo0586 ;
  assign new_n8707 = ~new_n8700 & new_n8706 ;
  assign new_n8708 = ~new_n8705 & ~new_n8707 ;
  assign new_n8709 = ~new_n8704 & new_n8708 ;
  assign new_n8710 = lo0593 & new_n3186 ;
  assign new_n8711 = lo0592 & new_n3202 ;
  assign new_n8712 = ~new_n3201 & ~new_n8711 ;
  assign new_n8713 = ~new_n8710 & new_n8712 ;
  assign new_n8714 = ~lo0063 & ~new_n8713 ;
  assign new_n8715 = lo0063 & new_n8713 ;
  assign new_n8716 = ~new_n8714 & ~new_n8715 ;
  assign new_n8717 = lo0591 & ~new_n8716 ;
  assign new_n8718 = ~lo0591 & new_n8714 ;
  assign new_n8719 = lo0063 & lo0594 ;
  assign new_n8720 = ~new_n8713 & new_n8719 ;
  assign new_n8721 = ~new_n8718 & ~new_n8720 ;
  assign new_n8722 = ~new_n8717 & new_n8721 ;
  assign new_n8723 = new_n3170 & ~new_n8722 ;
  assign new_n8724 = lo0589 & new_n3186 ;
  assign new_n8725 = lo0588 & new_n3202 ;
  assign new_n8726 = ~new_n3201 & ~new_n8725 ;
  assign new_n8727 = ~new_n8724 & new_n8726 ;
  assign new_n8728 = ~lo0063 & ~new_n8727 ;
  assign new_n8729 = lo0063 & new_n8727 ;
  assign new_n8730 = ~new_n8728 & ~new_n8729 ;
  assign new_n8731 = lo0587 & ~new_n8730 ;
  assign new_n8732 = ~lo0587 & new_n8728 ;
  assign new_n8733 = lo0063 & lo0590 ;
  assign new_n8734 = ~new_n8727 & new_n8733 ;
  assign new_n8735 = ~new_n8732 & ~new_n8734 ;
  assign new_n8736 = ~new_n8731 & new_n8735 ;
  assign new_n8737 = new_n3204 & ~new_n8736 ;
  assign new_n8738 = ~new_n3172 & ~new_n8737 ;
  assign new_n8739 = ~new_n8723 & new_n8738 ;
  assign new_n8740 = ~lo0061 & ~new_n8739 ;
  assign new_n8741 = lo0061 & new_n8739 ;
  assign new_n8742 = ~new_n8740 & ~new_n8741 ;
  assign new_n8743 = ~new_n8709 & ~new_n8742 ;
  assign new_n8744 = new_n8709 & new_n8740 ;
  assign new_n8745 = lo0597 & new_n3186 ;
  assign new_n8746 = lo0596 & new_n3559 ;
  assign new_n8747 = ~new_n3201 & ~new_n8746 ;
  assign new_n8748 = ~new_n8745 & new_n8747 ;
  assign new_n8749 = ~lo0065 & ~new_n8748 ;
  assign new_n8750 = lo0065 & new_n8748 ;
  assign new_n8751 = ~new_n8749 & ~new_n8750 ;
  assign new_n8752 = lo0595 & ~new_n8751 ;
  assign new_n8753 = ~lo0595 & new_n8749 ;
  assign new_n8754 = lo0065 & lo0598 ;
  assign new_n8755 = ~new_n8748 & new_n8754 ;
  assign new_n8756 = ~new_n8753 & ~new_n8755 ;
  assign new_n8757 = ~new_n8752 & new_n8756 ;
  assign new_n8758 = lo0061 & ~new_n8757 ;
  assign new_n8759 = ~new_n8739 & new_n8758 ;
  assign new_n8760 = ~new_n8744 & ~new_n8759 ;
  assign new_n8761 = ~new_n8743 & new_n8760 ;
  assign new_n8762 = new_n3169 & ~new_n8761 ;
  assign new_n8763 = ~new_n3160 & new_n6202 ;
  assign new_n8764 = new_n3264 & new_n6214 ;
  assign new_n8765 = lo0602 & new_n3258 ;
  assign new_n8766 = lo1337 & new_n3270 ;
  assign new_n8767 = lo0600 & new_n3274 ;
  assign new_n8768 = ~new_n8766 & ~new_n8767 ;
  assign new_n8769 = ~new_n8765 & new_n8768 ;
  assign new_n8770 = lo1335 & new_n3267 ;
  assign new_n8771 = lo1336 & new_n3246 ;
  assign new_n8772 = ~new_n8770 & ~new_n8771 ;
  assign new_n8773 = lo1334 & new_n3254 ;
  assign new_n8774 = lo0185 & new_n8264 ;
  assign new_n8775 = ~new_n8773 & ~new_n8774 ;
  assign new_n8776 = new_n8772 & new_n8775 ;
  assign new_n8777 = new_n8769 & new_n8776 ;
  assign new_n8778 = ~new_n8764 & new_n8777 ;
  assign new_n8779 = ~new_n8763 & new_n8778 ;
  assign new_n8780 = ~new_n8762 & new_n8779 ;
  assign new_n8781 = new_n6214 & new_n8020 ;
  assign new_n8782 = lo0593 & new_n8009 ;
  assign new_n8783 = new_n8017 & new_n8782 ;
  assign new_n8784 = ~new_n8022 & ~new_n8783 ;
  assign new_n8785 = ~new_n8781 & new_n8784 ;
  assign new_n8786 = new_n8017 & ~new_n8785 ;
  assign new_n8787 = new_n8780 & new_n8786 ;
  assign new_n8788 = ~new_n8017 & new_n8785 ;
  assign new_n8789 = ~new_n8786 & ~new_n8788 ;
  assign new_n8790 = ~new_n8780 & ~new_n8789 ;
  assign new_n8791 = ~new_n8017 & ~new_n8785 ;
  assign new_n8792 = new_n6202 & new_n8791 ;
  assign new_n8793 = ~new_n8790 & ~new_n8792 ;
  assign new_n8794 = ~new_n8787 & new_n8793 ;
  assign new_n8795 = ~new_n3112 & new_n8794 ;
  assign new_n8796 = new_n3112 & ~new_n8794 ;
  assign new_n8797 = ~new_n8795 & ~new_n8796 ;
  assign new_n8798 = new_n3737 & ~new_n5996 ;
  assign new_n8799 = new_n4180 & ~new_n4268 ;
  assign new_n8800 = ~new_n3819 & ~new_n8799 ;
  assign new_n8801 = ~new_n8798 & new_n8800 ;
  assign new_n8802 = new_n3736 & ~new_n8801 ;
  assign new_n8803 = ~new_n3736 & new_n8801 ;
  assign new_n8804 = ~new_n8802 & ~new_n8803 ;
  assign new_n8805 = ~new_n6225 & ~new_n8804 ;
  assign new_n8806 = new_n6225 & new_n8802 ;
  assign new_n8807 = new_n6470 & ~new_n8801 ;
  assign new_n8808 = ~new_n8806 & ~new_n8807 ;
  assign new_n8809 = ~new_n8805 & new_n8808 ;
  assign new_n8810 = lo0298 & ~new_n8809 ;
  assign new_n8811 = new_n3914 & ~new_n6917 ;
  assign new_n8812 = ~lo0297 & ~new_n6690 ;
  assign new_n8813 = ~new_n8811 & ~new_n8812 ;
  assign new_n8814 = ~lo0298 & ~new_n8813 ;
  assign new_n8815 = ~new_n8810 & ~new_n8814 ;
  assign new_n8816 = new_n3102 & ~new_n8815 ;
  assign new_n8817 = ~new_n3102 & ~new_n6461 ;
  assign new_n8818 = ~new_n8816 & ~new_n8817 ;
  assign new_n8819 = lo0204 & new_n3170 ;
  assign new_n8820 = lo0203 & new_n3173 ;
  assign new_n8821 = ~new_n3172 & ~new_n8820 ;
  assign new_n8822 = ~new_n8819 & new_n8821 ;
  assign new_n8823 = ~lo0059 & ~new_n8822 ;
  assign new_n8824 = lo0059 & new_n8822 ;
  assign new_n8825 = ~new_n8823 & ~new_n8824 ;
  assign new_n8826 = lo0202 & ~new_n8825 ;
  assign new_n8827 = ~lo0202 & new_n8823 ;
  assign new_n8828 = lo0059 & lo0205 ;
  assign new_n8829 = ~new_n8822 & new_n8828 ;
  assign new_n8830 = ~new_n8827 & ~new_n8829 ;
  assign new_n8831 = ~new_n8826 & new_n8830 ;
  assign new_n8832 = lo0201 & new_n3170 ;
  assign new_n8833 = lo0211 & new_n3173 ;
  assign new_n8834 = ~new_n3172 & ~new_n8833 ;
  assign new_n8835 = ~new_n8832 & new_n8834 ;
  assign new_n8836 = ~lo0059 & ~new_n8835 ;
  assign new_n8837 = lo0059 & new_n8835 ;
  assign new_n8838 = ~new_n8836 & ~new_n8837 ;
  assign new_n8839 = lo0210 & ~new_n8838 ;
  assign new_n8840 = ~lo0210 & new_n8836 ;
  assign new_n8841 = lo0059 & lo0212 ;
  assign new_n8842 = ~new_n8835 & new_n8841 ;
  assign new_n8843 = ~new_n8840 & ~new_n8842 ;
  assign new_n8844 = ~new_n8839 & new_n8843 ;
  assign new_n8845 = new_n3186 & ~new_n8844 ;
  assign new_n8846 = lo0208 & new_n3170 ;
  assign new_n8847 = lo0207 & new_n3204 ;
  assign new_n8848 = ~new_n3172 & ~new_n8847 ;
  assign new_n8849 = ~new_n8846 & new_n8848 ;
  assign new_n8850 = ~lo0061 & ~new_n8849 ;
  assign new_n8851 = lo0061 & new_n8849 ;
  assign new_n8852 = ~new_n8850 & ~new_n8851 ;
  assign new_n8853 = lo0206 & ~new_n8852 ;
  assign new_n8854 = ~lo0206 & new_n8850 ;
  assign new_n8855 = lo0061 & lo0209 ;
  assign new_n8856 = ~new_n8849 & new_n8855 ;
  assign new_n8857 = ~new_n8854 & ~new_n8856 ;
  assign new_n8858 = ~new_n8853 & new_n8857 ;
  assign new_n8859 = new_n3202 & ~new_n8858 ;
  assign new_n8860 = ~new_n3201 & ~new_n8859 ;
  assign new_n8861 = ~new_n8845 & new_n8860 ;
  assign new_n8862 = ~lo0063 & ~new_n8861 ;
  assign new_n8863 = lo0063 & new_n8861 ;
  assign new_n8864 = ~new_n8862 & ~new_n8863 ;
  assign new_n8865 = ~new_n8831 & ~new_n8864 ;
  assign new_n8866 = new_n8831 & new_n8862 ;
  assign new_n8867 = lo0215 & new_n3170 ;
  assign new_n8868 = lo0214 & new_n3204 ;
  assign new_n8869 = ~new_n3172 & ~new_n8868 ;
  assign new_n8870 = ~new_n8867 & new_n8869 ;
  assign new_n8871 = ~lo0061 & ~new_n8870 ;
  assign new_n8872 = lo0061 & new_n8870 ;
  assign new_n8873 = ~new_n8871 & ~new_n8872 ;
  assign new_n8874 = lo0213 & ~new_n8873 ;
  assign new_n8875 = ~lo0213 & new_n8871 ;
  assign new_n8876 = lo0061 & lo0216 ;
  assign new_n8877 = ~new_n8870 & new_n8876 ;
  assign new_n8878 = ~new_n8875 & ~new_n8877 ;
  assign new_n8879 = ~new_n8874 & new_n8878 ;
  assign new_n8880 = lo0063 & ~new_n8879 ;
  assign new_n8881 = ~new_n8861 & new_n8880 ;
  assign new_n8882 = ~new_n8866 & ~new_n8881 ;
  assign new_n8883 = ~new_n8865 & new_n8882 ;
  assign new_n8884 = new_n3169 & ~new_n8883 ;
  assign new_n8885 = ~new_n3160 & new_n6433 ;
  assign new_n8886 = new_n3264 & new_n6450 ;
  assign new_n8887 = lo0225 & new_n3258 ;
  assign new_n8888 = lo1298 & new_n3270 ;
  assign new_n8889 = lo0226 & new_n3274 ;
  assign new_n8890 = ~new_n8888 & ~new_n8889 ;
  assign new_n8891 = ~new_n8887 & new_n8890 ;
  assign new_n8892 = lo1296 & new_n3267 ;
  assign new_n8893 = lo1297 & new_n3246 ;
  assign new_n8894 = ~new_n8892 & ~new_n8893 ;
  assign new_n8895 = lo1295 & new_n3254 ;
  assign new_n8896 = lo0187 & new_n8264 ;
  assign new_n8897 = ~new_n8895 & ~new_n8896 ;
  assign new_n8898 = new_n8894 & new_n8897 ;
  assign new_n8899 = new_n8891 & new_n8898 ;
  assign new_n8900 = ~new_n8886 & new_n8899 ;
  assign new_n8901 = ~new_n8885 & new_n8900 ;
  assign new_n8902 = ~new_n8884 & new_n8901 ;
  assign new_n8903 = new_n8150 & ~new_n8902 ;
  assign new_n8904 = new_n6450 & new_n8020 ;
  assign new_n8905 = ~new_n8022 & ~new_n8904 ;
  assign new_n8906 = ~new_n8903 & new_n8905 ;
  assign new_n8907 = ~new_n8009 & ~new_n8906 ;
  assign new_n8908 = new_n8009 & new_n8906 ;
  assign new_n8909 = ~new_n8907 & ~new_n8908 ;
  assign new_n8910 = lo0201 & ~new_n8909 ;
  assign new_n8911 = ~lo0201 & new_n8907 ;
  assign new_n8912 = new_n6433 & new_n8009 ;
  assign new_n8913 = ~new_n8906 & new_n8912 ;
  assign new_n8914 = ~new_n8911 & ~new_n8913 ;
  assign new_n8915 = ~new_n8910 & new_n8914 ;
  assign new_n8916 = ~new_n3112 & new_n8915 ;
  assign new_n8917 = new_n3112 & ~new_n8915 ;
  assign new_n8918 = ~new_n8916 & ~new_n8917 ;
  assign new_n8919 = new_n3737 & ~new_n6225 ;
  assign new_n8920 = new_n3820 & ~new_n6461 ;
  assign new_n8921 = ~new_n3819 & ~new_n8920 ;
  assign new_n8922 = ~new_n8919 & new_n8921 ;
  assign new_n8923 = ~new_n3735 & ~new_n8922 ;
  assign new_n8924 = new_n3735 & new_n8922 ;
  assign new_n8925 = ~new_n8923 & ~new_n8924 ;
  assign new_n8926 = ~new_n4630 & ~new_n8925 ;
  assign new_n8927 = new_n4630 & new_n8923 ;
  assign new_n8928 = new_n6700 & ~new_n8922 ;
  assign new_n8929 = ~new_n8927 & ~new_n8928 ;
  assign new_n8930 = ~new_n8926 & new_n8929 ;
  assign new_n8931 = lo0298 & ~new_n8930 ;
  assign new_n8932 = ~lo0297 & ~new_n6917 ;
  assign new_n8933 = new_n3914 & ~new_n7138 ;
  assign new_n8934 = ~new_n8932 & ~new_n8933 ;
  assign new_n8935 = ~lo0298 & ~new_n8934 ;
  assign new_n8936 = ~new_n8931 & ~new_n8935 ;
  assign new_n8937 = new_n3102 & ~new_n8936 ;
  assign new_n8938 = ~new_n3102 & ~new_n6690 ;
  assign new_n8939 = ~new_n8937 & ~new_n8938 ;
  assign new_n8940 = lo0562 & new_n3186 ;
  assign new_n8941 = lo0561 & new_n3559 ;
  assign new_n8942 = ~new_n3201 & ~new_n8941 ;
  assign new_n8943 = ~new_n8940 & new_n8942 ;
  assign new_n8944 = ~lo0065 & ~new_n8943 ;
  assign new_n8945 = lo0065 & new_n8943 ;
  assign new_n8946 = ~new_n8944 & ~new_n8945 ;
  assign new_n8947 = lo0560 & ~new_n8946 ;
  assign new_n8948 = ~lo0560 & new_n8944 ;
  assign new_n8949 = lo0065 & lo0563 ;
  assign new_n8950 = ~new_n8943 & new_n8949 ;
  assign new_n8951 = ~new_n8948 & ~new_n8950 ;
  assign new_n8952 = ~new_n8947 & new_n8951 ;
  assign new_n8953 = lo0570 & new_n3186 ;
  assign new_n8954 = lo0569 & new_n3559 ;
  assign new_n8955 = ~new_n3201 & ~new_n8954 ;
  assign new_n8956 = ~new_n8953 & new_n8955 ;
  assign new_n8957 = ~lo0065 & ~new_n8956 ;
  assign new_n8958 = lo0065 & new_n8956 ;
  assign new_n8959 = ~new_n8957 & ~new_n8958 ;
  assign new_n8960 = lo0568 & ~new_n8959 ;
  assign new_n8961 = ~lo0568 & new_n8957 ;
  assign new_n8962 = lo0065 & lo0571 ;
  assign new_n8963 = ~new_n8956 & new_n8962 ;
  assign new_n8964 = ~new_n8961 & ~new_n8963 ;
  assign new_n8965 = ~new_n8960 & new_n8964 ;
  assign new_n8966 = new_n3170 & ~new_n8965 ;
  assign new_n8967 = lo0566 & new_n3186 ;
  assign new_n8968 = lo0565 & new_n3202 ;
  assign new_n8969 = ~new_n3201 & ~new_n8968 ;
  assign new_n8970 = ~new_n8967 & new_n8969 ;
  assign new_n8971 = ~lo0063 & ~new_n8970 ;
  assign new_n8972 = lo0063 & new_n8970 ;
  assign new_n8973 = ~new_n8971 & ~new_n8972 ;
  assign new_n8974 = lo0564 & ~new_n8973 ;
  assign new_n8975 = ~lo0564 & new_n8971 ;
  assign new_n8976 = lo0063 & lo0567 ;
  assign new_n8977 = ~new_n8970 & new_n8976 ;
  assign new_n8978 = ~new_n8975 & ~new_n8977 ;
  assign new_n8979 = ~new_n8974 & new_n8978 ;
  assign new_n8980 = new_n3173 & ~new_n8979 ;
  assign new_n8981 = ~new_n3172 & ~new_n8980 ;
  assign new_n8982 = ~new_n8966 & new_n8981 ;
  assign new_n8983 = ~lo0059 & ~new_n8982 ;
  assign new_n8984 = lo0059 & new_n8982 ;
  assign new_n8985 = ~new_n8983 & ~new_n8984 ;
  assign new_n8986 = ~new_n8952 & ~new_n8985 ;
  assign new_n8987 = new_n8952 & new_n8983 ;
  assign new_n8988 = lo0574 & new_n3186 ;
  assign new_n8989 = lo0573 & new_n3202 ;
  assign new_n8990 = ~new_n3201 & ~new_n8989 ;
  assign new_n8991 = ~new_n8988 & new_n8990 ;
  assign new_n8992 = ~lo0063 & ~new_n8991 ;
  assign new_n8993 = lo0063 & new_n8991 ;
  assign new_n8994 = ~new_n8992 & ~new_n8993 ;
  assign new_n8995 = lo0572 & ~new_n8994 ;
  assign new_n8996 = ~lo0572 & new_n8992 ;
  assign new_n8997 = lo0063 & lo0575 ;
  assign new_n8998 = ~new_n8991 & new_n8997 ;
  assign new_n8999 = ~new_n8996 & ~new_n8998 ;
  assign new_n9000 = ~new_n8995 & new_n8999 ;
  assign new_n9001 = lo0059 & ~new_n9000 ;
  assign new_n9002 = ~new_n8982 & new_n9001 ;
  assign new_n9003 = ~new_n8987 & ~new_n9002 ;
  assign new_n9004 = ~new_n8986 & new_n9003 ;
  assign new_n9005 = new_n3169 & ~new_n9004 ;
  assign new_n9006 = ~new_n3160 & new_n6667 ;
  assign new_n9007 = new_n3264 & ~new_n6679 ;
  assign new_n9008 = lo1333 & new_n3254 ;
  assign new_n9009 = lo1376 & new_n3270 ;
  assign new_n9010 = lo0580 & new_n3274 ;
  assign new_n9011 = ~new_n9009 & ~new_n9010 ;
  assign new_n9012 = ~new_n9008 & new_n9011 ;
  assign new_n9013 = lo1374 & new_n3267 ;
  assign new_n9014 = lo1375 & new_n3246 ;
  assign new_n9015 = lo0582 & new_n3258 ;
  assign new_n9016 = ~new_n9014 & ~new_n9015 ;
  assign new_n9017 = ~new_n9013 & new_n9016 ;
  assign new_n9018 = new_n9012 & new_n9017 ;
  assign new_n9019 = ~new_n9007 & new_n9018 ;
  assign new_n9020 = ~new_n9006 & new_n9019 ;
  assign new_n9021 = ~new_n9005 & new_n9020 ;
  assign new_n9022 = ~new_n6679 & new_n8020 ;
  assign new_n9023 = lo0570 & new_n8009 ;
  assign new_n9024 = new_n8017 & new_n9023 ;
  assign new_n9025 = ~new_n8022 & ~new_n9024 ;
  assign new_n9026 = ~new_n9022 & new_n9025 ;
  assign new_n9027 = new_n8017 & ~new_n9026 ;
  assign new_n9028 = new_n9021 & new_n9027 ;
  assign new_n9029 = ~new_n8017 & new_n9026 ;
  assign new_n9030 = ~new_n9027 & ~new_n9029 ;
  assign new_n9031 = ~new_n9021 & ~new_n9030 ;
  assign new_n9032 = ~new_n8017 & ~new_n9026 ;
  assign new_n9033 = new_n6667 & new_n9032 ;
  assign new_n9034 = ~new_n9031 & ~new_n9033 ;
  assign new_n9035 = ~new_n9028 & new_n9034 ;
  assign new_n9036 = ~new_n3112 & new_n9035 ;
  assign new_n9037 = new_n3112 & ~new_n9035 ;
  assign new_n9038 = ~new_n9036 & ~new_n9037 ;
  assign new_n9039 = new_n3737 & ~new_n6461 ;
  assign new_n9040 = new_n4180 & ~new_n4992 ;
  assign new_n9041 = ~new_n3819 & ~new_n9040 ;
  assign new_n9042 = ~new_n9039 & new_n9041 ;
  assign new_n9043 = new_n3736 & ~new_n9042 ;
  assign new_n9044 = ~new_n3736 & new_n9042 ;
  assign new_n9045 = ~new_n9043 & ~new_n9044 ;
  assign new_n9046 = ~new_n6690 & ~new_n9045 ;
  assign new_n9047 = new_n6690 & new_n9043 ;
  assign new_n9048 = new_n6925 & ~new_n9042 ;
  assign new_n9049 = ~new_n9047 & ~new_n9048 ;
  assign new_n9050 = ~new_n9046 & new_n9049 ;
  assign new_n9051 = lo0298 & ~new_n9050 ;
  assign new_n9052 = ~new_n2619 & new_n3914 ;
  assign new_n9053 = ~lo0297 & ~new_n7138 ;
  assign new_n9054 = ~new_n9052 & ~new_n9053 ;
  assign new_n9055 = ~lo0298 & ~new_n9054 ;
  assign new_n9056 = ~new_n9051 & ~new_n9055 ;
  assign new_n9057 = new_n3102 & ~new_n9056 ;
  assign new_n9058 = ~new_n3102 & ~new_n6917 ;
  assign new_n9059 = ~new_n9057 & ~new_n9058 ;
  assign new_n9060 = lo0624 & new_n3170 ;
  assign new_n9061 = lo0623 & new_n3173 ;
  assign new_n9062 = ~new_n3172 & ~new_n9061 ;
  assign new_n9063 = ~new_n9060 & new_n9062 ;
  assign new_n9064 = ~lo0059 & ~new_n9063 ;
  assign new_n9065 = lo0059 & new_n9063 ;
  assign new_n9066 = ~new_n9064 & ~new_n9065 ;
  assign new_n9067 = lo0622 & ~new_n9066 ;
  assign new_n9068 = ~lo0622 & new_n9064 ;
  assign new_n9069 = lo0059 & lo0625 ;
  assign new_n9070 = ~new_n9063 & new_n9069 ;
  assign new_n9071 = ~new_n9068 & ~new_n9070 ;
  assign new_n9072 = ~new_n9067 & new_n9071 ;
  assign new_n9073 = lo0632 & new_n3170 ;
  assign new_n9074 = lo0631 & new_n3204 ;
  assign new_n9075 = ~new_n3172 & ~new_n9074 ;
  assign new_n9076 = ~new_n9073 & new_n9075 ;
  assign new_n9077 = ~lo0061 & ~new_n9076 ;
  assign new_n9078 = lo0061 & new_n9076 ;
  assign new_n9079 = ~new_n9077 & ~new_n9078 ;
  assign new_n9080 = lo0630 & ~new_n9079 ;
  assign new_n9081 = ~lo0630 & new_n9077 ;
  assign new_n9082 = lo0061 & lo0633 ;
  assign new_n9083 = ~new_n9076 & new_n9082 ;
  assign new_n9084 = ~new_n9081 & ~new_n9083 ;
  assign new_n9085 = ~new_n9080 & new_n9084 ;
  assign new_n9086 = new_n3186 & ~new_n9085 ;
  assign new_n9087 = lo0628 & new_n3170 ;
  assign new_n9088 = lo0627 & new_n3204 ;
  assign new_n9089 = ~new_n3172 & ~new_n9088 ;
  assign new_n9090 = ~new_n9087 & new_n9089 ;
  assign new_n9091 = ~lo0061 & ~new_n9090 ;
  assign new_n9092 = lo0061 & new_n9090 ;
  assign new_n9093 = ~new_n9091 & ~new_n9092 ;
  assign new_n9094 = lo0626 & ~new_n9093 ;
  assign new_n9095 = ~lo0626 & new_n9091 ;
  assign new_n9096 = lo0061 & lo0629 ;
  assign new_n9097 = ~new_n9090 & new_n9096 ;
  assign new_n9098 = ~new_n9095 & ~new_n9097 ;
  assign new_n9099 = ~new_n9094 & new_n9098 ;
  assign new_n9100 = new_n3559 & ~new_n9099 ;
  assign new_n9101 = ~new_n3201 & ~new_n9100 ;
  assign new_n9102 = ~new_n9086 & new_n9101 ;
  assign new_n9103 = ~lo0065 & ~new_n9102 ;
  assign new_n9104 = lo0065 & new_n9102 ;
  assign new_n9105 = ~new_n9103 & ~new_n9104 ;
  assign new_n9106 = ~new_n9072 & ~new_n9105 ;
  assign new_n9107 = new_n9072 & new_n9103 ;
  assign new_n9108 = lo0636 & new_n3170 ;
  assign new_n9109 = lo0635 & new_n3173 ;
  assign new_n9110 = ~new_n3172 & ~new_n9109 ;
  assign new_n9111 = ~new_n9108 & new_n9110 ;
  assign new_n9112 = ~lo0059 & ~new_n9111 ;
  assign new_n9113 = lo0059 & new_n9111 ;
  assign new_n9114 = ~new_n9112 & ~new_n9113 ;
  assign new_n9115 = lo0634 & ~new_n9114 ;
  assign new_n9116 = ~lo0634 & new_n9112 ;
  assign new_n9117 = lo0059 & lo0637 ;
  assign new_n9118 = ~new_n9111 & new_n9117 ;
  assign new_n9119 = ~new_n9116 & ~new_n9118 ;
  assign new_n9120 = ~new_n9115 & new_n9119 ;
  assign new_n9121 = lo0065 & ~new_n9120 ;
  assign new_n9122 = ~new_n9102 & new_n9121 ;
  assign new_n9123 = ~new_n9107 & ~new_n9122 ;
  assign new_n9124 = ~new_n9106 & new_n9123 ;
  assign new_n9125 = new_n3169 & ~new_n9124 ;
  assign new_n9126 = ~new_n3160 & new_n6899 ;
  assign new_n9127 = new_n3264 & ~new_n6906 ;
  assign new_n9128 = lo1348 & new_n3254 ;
  assign new_n9129 = lo1370 & new_n3270 ;
  assign new_n9130 = lo0642 & new_n3274 ;
  assign new_n9131 = ~new_n9129 & ~new_n9130 ;
  assign new_n9132 = ~new_n9128 & new_n9131 ;
  assign new_n9133 = lo1368 & new_n3267 ;
  assign new_n9134 = lo1369 & new_n3246 ;
  assign new_n9135 = lo0644 & new_n3258 ;
  assign new_n9136 = ~new_n9134 & ~new_n9135 ;
  assign new_n9137 = ~new_n9133 & new_n9136 ;
  assign new_n9138 = new_n9132 & new_n9137 ;
  assign new_n9139 = ~new_n9127 & new_n9138 ;
  assign new_n9140 = ~new_n9126 & new_n9139 ;
  assign new_n9141 = ~new_n9125 & new_n9140 ;
  assign new_n9142 = new_n8150 & ~new_n9141 ;
  assign new_n9143 = lo0198 & ~lo0199 ;
  assign new_n9144 = new_n3100 & ~new_n6906 ;
  assign new_n9145 = ~new_n9143 & ~new_n9144 ;
  assign new_n9146 = ~lo0197 & ~new_n8009 ;
  assign new_n9147 = new_n8017 & new_n9146 ;
  assign new_n9148 = ~new_n9145 & new_n9147 ;
  assign new_n9149 = ~new_n8022 & ~new_n9148 ;
  assign new_n9150 = ~new_n9142 & new_n9149 ;
  assign new_n9151 = ~new_n8009 & ~new_n9150 ;
  assign new_n9152 = new_n8009 & new_n9150 ;
  assign new_n9153 = ~new_n9151 & ~new_n9152 ;
  assign new_n9154 = lo0632 & ~new_n9153 ;
  assign new_n9155 = ~lo0632 & new_n9151 ;
  assign new_n9156 = new_n6899 & new_n8009 ;
  assign new_n9157 = ~new_n9150 & new_n9156 ;
  assign new_n9158 = ~new_n9155 & ~new_n9157 ;
  assign new_n9159 = ~new_n9154 & new_n9158 ;
  assign new_n9160 = ~new_n3112 & new_n9159 ;
  assign new_n9161 = new_n3112 & ~new_n9159 ;
  assign new_n9162 = ~new_n9160 & ~new_n9161 ;
  assign new_n9163 = ~new_n8013 & ~new_n9143 ;
  assign new_n9164 = ~lo0200 & new_n3099 ;
  assign new_n9165 = new_n9163 & new_n9164 ;
  assign new_n9166 = ~new_n7138 & ~new_n9165 ;
  assign new_n9167 = lo0198 & new_n9165 ;
  assign new_n9168 = new_n2827 & new_n5669 ;
  assign new_n9169 = ~new_n5187 & new_n9168 ;
  assign new_n9170 = ~lo0297 & ~lo0298 ;
  assign new_n9171 = ~new_n2619 & new_n9170 ;
  assign new_n9172 = lo0299 & ~new_n5276 ;
  assign new_n9173 = ~lo0299 & ~new_n6690 ;
  assign new_n9174 = ~new_n9172 & ~new_n9173 ;
  assign new_n9175 = lo0297 & ~new_n9174 ;
  assign new_n9176 = ~new_n8932 & ~new_n9175 ;
  assign new_n9177 = lo0298 & ~new_n9176 ;
  assign new_n9178 = ~new_n9171 & ~new_n9177 ;
  assign new_n9179 = ~lo0300 & ~new_n9178 ;
  assign new_n9180 = ~new_n9169 & ~new_n9179 ;
  assign new_n9181 = new_n9167 & ~new_n9180 ;
  assign new_n9182 = ~new_n9166 & ~new_n9181 ;
  assign new_n9183 = lo0786 & new_n3186 ;
  assign new_n9184 = lo0785 & new_n3559 ;
  assign new_n9185 = ~new_n3201 & ~new_n9184 ;
  assign new_n9186 = ~new_n9183 & new_n9185 ;
  assign new_n9187 = ~lo0065 & ~new_n9186 ;
  assign new_n9188 = lo0065 & new_n9186 ;
  assign new_n9189 = ~new_n9187 & ~new_n9188 ;
  assign new_n9190 = lo0784 & ~new_n9189 ;
  assign new_n9191 = ~lo0784 & new_n9187 ;
  assign new_n9192 = lo0065 & lo0787 ;
  assign new_n9193 = ~new_n9186 & new_n9192 ;
  assign new_n9194 = ~new_n9191 & ~new_n9193 ;
  assign new_n9195 = ~new_n9190 & new_n9194 ;
  assign new_n9196 = lo0794 & new_n3186 ;
  assign new_n9197 = lo0793 & new_n3202 ;
  assign new_n9198 = ~new_n3201 & ~new_n9197 ;
  assign new_n9199 = ~new_n9196 & new_n9198 ;
  assign new_n9200 = ~lo0063 & ~new_n9199 ;
  assign new_n9201 = lo0063 & new_n9199 ;
  assign new_n9202 = ~new_n9200 & ~new_n9201 ;
  assign new_n9203 = lo0792 & ~new_n9202 ;
  assign new_n9204 = ~lo0792 & new_n9200 ;
  assign new_n9205 = lo0063 & lo0795 ;
  assign new_n9206 = ~new_n9199 & new_n9205 ;
  assign new_n9207 = ~new_n9204 & ~new_n9206 ;
  assign new_n9208 = ~new_n9203 & new_n9207 ;
  assign new_n9209 = new_n3170 & ~new_n9208 ;
  assign new_n9210 = lo0790 & new_n3186 ;
  assign new_n9211 = lo0789 & new_n3202 ;
  assign new_n9212 = ~new_n3201 & ~new_n9211 ;
  assign new_n9213 = ~new_n9210 & new_n9212 ;
  assign new_n9214 = ~lo0063 & ~new_n9213 ;
  assign new_n9215 = lo0063 & new_n9213 ;
  assign new_n9216 = ~new_n9214 & ~new_n9215 ;
  assign new_n9217 = lo0788 & ~new_n9216 ;
  assign new_n9218 = ~lo0788 & new_n9214 ;
  assign new_n9219 = lo0063 & lo0791 ;
  assign new_n9220 = ~new_n9213 & new_n9219 ;
  assign new_n9221 = ~new_n9218 & ~new_n9220 ;
  assign new_n9222 = ~new_n9217 & new_n9221 ;
  assign new_n9223 = new_n3204 & ~new_n9222 ;
  assign new_n9224 = ~new_n3172 & ~new_n9223 ;
  assign new_n9225 = ~new_n9209 & new_n9224 ;
  assign new_n9226 = ~lo0061 & ~new_n9225 ;
  assign new_n9227 = lo0061 & new_n9225 ;
  assign new_n9228 = ~new_n9226 & ~new_n9227 ;
  assign new_n9229 = ~new_n9195 & ~new_n9228 ;
  assign new_n9230 = new_n9195 & new_n9226 ;
  assign new_n9231 = lo0798 & new_n3186 ;
  assign new_n9232 = lo0797 & new_n3559 ;
  assign new_n9233 = ~new_n3201 & ~new_n9232 ;
  assign new_n9234 = ~new_n9231 & new_n9233 ;
  assign new_n9235 = ~lo0065 & ~new_n9234 ;
  assign new_n9236 = lo0065 & new_n9234 ;
  assign new_n9237 = ~new_n9235 & ~new_n9236 ;
  assign new_n9238 = lo0796 & ~new_n9237 ;
  assign new_n9239 = ~lo0796 & new_n9235 ;
  assign new_n9240 = lo0065 & lo0799 ;
  assign new_n9241 = ~new_n9234 & new_n9240 ;
  assign new_n9242 = ~new_n9239 & ~new_n9241 ;
  assign new_n9243 = ~new_n9238 & new_n9242 ;
  assign new_n9244 = lo0061 & ~new_n9243 ;
  assign new_n9245 = ~new_n9225 & new_n9244 ;
  assign new_n9246 = ~new_n9230 & ~new_n9245 ;
  assign new_n9247 = ~new_n9229 & new_n9246 ;
  assign new_n9248 = new_n3169 & ~new_n9247 ;
  assign new_n9249 = ~new_n3160 & new_n7122 ;
  assign new_n9250 = new_n3264 & ~new_n7127 ;
  assign new_n9251 = lo1385 & new_n3246 ;
  assign new_n9252 = lo1382 & new_n3270 ;
  assign new_n9253 = lo0803 & new_n3274 ;
  assign new_n9254 = ~new_n9252 & ~new_n9253 ;
  assign new_n9255 = ~new_n9251 & new_n9254 ;
  assign new_n9256 = lo1380 & new_n3254 ;
  assign new_n9257 = lo0805 & new_n3258 ;
  assign new_n9258 = ~new_n9256 & ~new_n9257 ;
  assign new_n9259 = lo1383 & new_n3267 ;
  assign new_n9260 = lo1384 & new_n8264 ;
  assign new_n9261 = ~new_n9259 & ~new_n9260 ;
  assign new_n9262 = new_n9258 & new_n9261 ;
  assign new_n9263 = new_n9255 & new_n9262 ;
  assign new_n9264 = ~new_n9250 & new_n9263 ;
  assign new_n9265 = ~new_n9249 & new_n9264 ;
  assign new_n9266 = ~new_n9248 & new_n9265 ;
  assign new_n9267 = ~lo0198 & ~lo0199 ;
  assign new_n9268 = new_n3100 & ~new_n7127 ;
  assign new_n9269 = ~new_n9267 & ~new_n9268 ;
  assign new_n9270 = new_n9147 & ~new_n9269 ;
  assign new_n9271 = lo0794 & new_n8009 ;
  assign new_n9272 = new_n8017 & new_n9271 ;
  assign new_n9273 = ~new_n8022 & ~new_n9272 ;
  assign new_n9274 = ~new_n9270 & new_n9273 ;
  assign new_n9275 = new_n8017 & ~new_n9274 ;
  assign new_n9276 = new_n9266 & new_n9275 ;
  assign new_n9277 = ~new_n8017 & new_n9274 ;
  assign new_n9278 = ~new_n9275 & ~new_n9277 ;
  assign new_n9279 = ~new_n9266 & ~new_n9278 ;
  assign new_n9280 = ~new_n8017 & ~new_n9274 ;
  assign new_n9281 = new_n7122 & new_n9280 ;
  assign new_n9282 = ~new_n9279 & ~new_n9281 ;
  assign new_n9283 = ~new_n9276 & new_n9282 ;
  assign new_n9284 = ~new_n3112 & new_n9283 ;
  assign new_n9285 = new_n3112 & ~new_n9283 ;
  assign new_n9286 = ~new_n9284 & ~new_n9285 ;
  assign new_n9287 = ~new_n2619 & ~new_n9165 ;
  assign new_n9288 = new_n2911 & ~new_n5560 ;
  assign new_n9289 = lo0300 & ~new_n5472 ;
  assign new_n9290 = ~lo0300 & ~new_n6917 ;
  assign new_n9291 = ~new_n9289 & ~new_n9290 ;
  assign new_n9292 = ~lo0299 & ~new_n9291 ;
  assign new_n9293 = ~new_n9288 & ~new_n9292 ;
  assign new_n9294 = ~lo0846 & new_n5669 ;
  assign new_n9295 = ~new_n9293 & new_n9294 ;
  assign new_n9296 = lo0298 & ~new_n7138 ;
  assign new_n9297 = ~lo0299 & ~new_n2739 ;
  assign new_n9298 = ~new_n3094 & ~new_n9297 ;
  assign new_n9299 = ~lo0298 & lo0846 ;
  assign new_n9300 = ~new_n9298 & new_n9299 ;
  assign new_n9301 = ~new_n9296 & ~new_n9300 ;
  assign new_n9302 = new_n2915 & ~new_n9301 ;
  assign new_n9303 = ~new_n9295 & ~new_n9302 ;
  assign new_n9304 = new_n9167 & ~new_n9303 ;
  assign new_n9305 = ~new_n9287 & ~new_n9304 ;
  assign new_n9306 = lo0745 & new_n3170 ;
  assign new_n9307 = lo0744 & new_n3173 ;
  assign new_n9308 = ~new_n3172 & ~new_n9307 ;
  assign new_n9309 = ~new_n9306 & new_n9308 ;
  assign new_n9310 = ~lo0059 & ~new_n9309 ;
  assign new_n9311 = lo0059 & new_n9309 ;
  assign new_n9312 = ~new_n9310 & ~new_n9311 ;
  assign new_n9313 = lo0743 & ~new_n9312 ;
  assign new_n9314 = ~lo0743 & new_n9310 ;
  assign new_n9315 = lo0059 & lo0746 ;
  assign new_n9316 = ~new_n9309 & new_n9315 ;
  assign new_n9317 = ~new_n9314 & ~new_n9316 ;
  assign new_n9318 = ~new_n9313 & new_n9317 ;
  assign new_n9319 = lo0742 & new_n3170 ;
  assign new_n9320 = lo0752 & new_n3173 ;
  assign new_n9321 = ~new_n3172 & ~new_n9320 ;
  assign new_n9322 = ~new_n9319 & new_n9321 ;
  assign new_n9323 = ~lo0059 & ~new_n9322 ;
  assign new_n9324 = lo0059 & new_n9322 ;
  assign new_n9325 = ~new_n9323 & ~new_n9324 ;
  assign new_n9326 = lo0751 & ~new_n9325 ;
  assign new_n9327 = ~lo0751 & new_n9323 ;
  assign new_n9328 = lo0059 & lo0753 ;
  assign new_n9329 = ~new_n9322 & new_n9328 ;
  assign new_n9330 = ~new_n9327 & ~new_n9329 ;
  assign new_n9331 = ~new_n9326 & new_n9330 ;
  assign new_n9332 = new_n3186 & ~new_n9331 ;
  assign new_n9333 = lo0749 & new_n3170 ;
  assign new_n9334 = lo0748 & new_n3204 ;
  assign new_n9335 = ~new_n3172 & ~new_n9334 ;
  assign new_n9336 = ~new_n9333 & new_n9335 ;
  assign new_n9337 = ~lo0061 & ~new_n9336 ;
  assign new_n9338 = lo0061 & new_n9336 ;
  assign new_n9339 = ~new_n9337 & ~new_n9338 ;
  assign new_n9340 = lo0747 & ~new_n9339 ;
  assign new_n9341 = ~lo0747 & new_n9337 ;
  assign new_n9342 = lo0061 & lo0750 ;
  assign new_n9343 = ~new_n9336 & new_n9342 ;
  assign new_n9344 = ~new_n9341 & ~new_n9343 ;
  assign new_n9345 = ~new_n9340 & new_n9344 ;
  assign new_n9346 = new_n3202 & ~new_n9345 ;
  assign new_n9347 = ~new_n3201 & ~new_n9346 ;
  assign new_n9348 = ~new_n9332 & new_n9347 ;
  assign new_n9349 = ~lo0063 & ~new_n9348 ;
  assign new_n9350 = lo0063 & new_n9348 ;
  assign new_n9351 = ~new_n9349 & ~new_n9350 ;
  assign new_n9352 = ~new_n9318 & ~new_n9351 ;
  assign new_n9353 = new_n9318 & new_n9349 ;
  assign new_n9354 = lo0756 & new_n3170 ;
  assign new_n9355 = lo0755 & new_n3204 ;
  assign new_n9356 = ~new_n3172 & ~new_n9355 ;
  assign new_n9357 = ~new_n9354 & new_n9356 ;
  assign new_n9358 = ~lo0061 & ~new_n9357 ;
  assign new_n9359 = lo0061 & new_n9357 ;
  assign new_n9360 = ~new_n9358 & ~new_n9359 ;
  assign new_n9361 = lo0754 & ~new_n9360 ;
  assign new_n9362 = ~lo0754 & new_n9358 ;
  assign new_n9363 = lo0061 & lo0757 ;
  assign new_n9364 = ~new_n9357 & new_n9363 ;
  assign new_n9365 = ~new_n9362 & ~new_n9364 ;
  assign new_n9366 = ~new_n9361 & new_n9365 ;
  assign new_n9367 = lo0063 & ~new_n9366 ;
  assign new_n9368 = ~new_n9348 & new_n9367 ;
  assign new_n9369 = ~new_n9353 & ~new_n9368 ;
  assign new_n9370 = ~new_n9352 & new_n9369 ;
  assign new_n9371 = new_n3169 & ~new_n9370 ;
  assign new_n9372 = new_n2586 & ~new_n3160 ;
  assign new_n9373 = lo0760 & new_n8264 ;
  assign new_n9374 = lo0761 & new_n3258 ;
  assign new_n9375 = ~new_n9373 & ~new_n9374 ;
  assign new_n9376 = lo1360 & new_n3254 ;
  assign new_n9377 = lo1362 & new_n3267 ;
  assign new_n9378 = ~new_n9376 & ~new_n9377 ;
  assign new_n9379 = new_n9375 & new_n9378 ;
  assign new_n9380 = new_n2598 & new_n3264 ;
  assign new_n9381 = lo1363 & new_n3246 ;
  assign new_n9382 = lo1361 & new_n3270 ;
  assign new_n9383 = lo0759 & new_n3274 ;
  assign new_n9384 = ~new_n9382 & ~new_n9383 ;
  assign new_n9385 = ~new_n9381 & new_n9384 ;
  assign new_n9386 = ~new_n9380 & new_n9385 ;
  assign new_n9387 = new_n9379 & new_n9386 ;
  assign new_n9388 = ~new_n9372 & new_n9387 ;
  assign new_n9389 = ~new_n9371 & new_n9388 ;
  assign new_n9390 = new_n8150 & ~new_n9389 ;
  assign new_n9391 = new_n2598 & new_n3100 ;
  assign new_n9392 = ~lo0197 & ~new_n9391 ;
  assign new_n9393 = ~new_n8009 & new_n8017 ;
  assign new_n9394 = ~new_n9392 & new_n9393 ;
  assign new_n9395 = ~new_n8022 & ~new_n9394 ;
  assign new_n9396 = ~new_n9390 & new_n9395 ;
  assign new_n9397 = ~new_n8009 & ~new_n9396 ;
  assign new_n9398 = new_n8009 & new_n9396 ;
  assign new_n9399 = ~new_n9397 & ~new_n9398 ;
  assign new_n9400 = lo0742 & ~new_n9399 ;
  assign new_n9401 = ~lo0742 & new_n9397 ;
  assign new_n9402 = new_n2586 & new_n8009 ;
  assign new_n9403 = ~new_n9396 & new_n9402 ;
  assign new_n9404 = ~new_n9401 & ~new_n9403 ;
  assign new_n9405 = ~new_n9400 & new_n9404 ;
  assign new_n9406 = ~new_n3112 & new_n9405 ;
  assign new_n9407 = new_n3112 & ~new_n9405 ;
  assign new_n9408 = ~new_n9406 & ~new_n9407 ;
  assign new_n9409 = lo0760 & new_n9143 ;
  assign new_n9410 = new_n3116 & new_n9409 ;
  assign new_n9411 = ~new_n3112 & ~new_n9410 ;
  assign new_n9412 = new_n3112 & new_n9410 ;
  assign new_n9413 = ~new_n9411 & ~new_n9412 ;
  assign new_n9414 = new_n9408 & ~new_n9413 ;
  assign new_n9415 = new_n9408 & ~new_n9414 ;
  assign new_n9416 = ~new_n9305 & ~new_n9415 ;
  assign new_n9417 = ~new_n9408 & ~new_n9413 ;
  assign new_n9418 = new_n9305 & new_n9417 ;
  assign new_n9419 = ~new_n9416 & ~new_n9418 ;
  assign new_n9420 = new_n9286 & ~new_n9419 ;
  assign new_n9421 = new_n9286 & ~new_n9420 ;
  assign new_n9422 = ~new_n9182 & ~new_n9421 ;
  assign new_n9423 = ~new_n9286 & ~new_n9419 ;
  assign new_n9424 = new_n9182 & new_n9423 ;
  assign new_n9425 = ~new_n9422 & ~new_n9424 ;
  assign new_n9426 = new_n9162 & ~new_n9425 ;
  assign new_n9427 = new_n9162 & ~new_n9426 ;
  assign new_n9428 = ~new_n9059 & ~new_n9427 ;
  assign new_n9429 = ~new_n9162 & ~new_n9425 ;
  assign new_n9430 = new_n9059 & new_n9429 ;
  assign new_n9431 = ~new_n9428 & ~new_n9430 ;
  assign new_n9432 = new_n9038 & ~new_n9431 ;
  assign new_n9433 = new_n9038 & ~new_n9432 ;
  assign new_n9434 = ~new_n8939 & ~new_n9433 ;
  assign new_n9435 = ~new_n9038 & ~new_n9431 ;
  assign new_n9436 = new_n8939 & new_n9435 ;
  assign new_n9437 = ~new_n9434 & ~new_n9436 ;
  assign new_n9438 = new_n8918 & ~new_n9437 ;
  assign new_n9439 = new_n8918 & ~new_n9438 ;
  assign new_n9440 = ~new_n8818 & ~new_n9439 ;
  assign new_n9441 = ~new_n8918 & ~new_n9437 ;
  assign new_n9442 = new_n8818 & new_n9441 ;
  assign new_n9443 = ~new_n9440 & ~new_n9442 ;
  assign new_n9444 = new_n8797 & ~new_n9443 ;
  assign new_n9445 = new_n8797 & ~new_n9444 ;
  assign new_n9446 = ~new_n8696 & ~new_n9445 ;
  assign new_n9447 = ~new_n8797 & ~new_n9443 ;
  assign new_n9448 = new_n8696 & new_n9447 ;
  assign new_n9449 = ~new_n9446 & ~new_n9448 ;
  assign new_n9450 = new_n8675 & ~new_n9449 ;
  assign new_n9451 = new_n8675 & ~new_n9450 ;
  assign new_n9452 = ~new_n8575 & ~new_n9451 ;
  assign new_n9453 = ~new_n8675 & ~new_n9449 ;
  assign new_n9454 = new_n8575 & new_n9453 ;
  assign new_n9455 = ~new_n9452 & ~new_n9454 ;
  assign new_n9456 = new_n8554 & ~new_n9455 ;
  assign new_n9457 = new_n8554 & ~new_n9456 ;
  assign new_n9458 = ~new_n8449 & ~new_n9457 ;
  assign new_n9459 = ~new_n8554 & ~new_n9455 ;
  assign new_n9460 = new_n8449 & new_n9459 ;
  assign new_n9461 = ~new_n9458 & ~new_n9460 ;
  assign new_n9462 = new_n8428 & ~new_n9461 ;
  assign new_n9463 = new_n8428 & ~new_n9462 ;
  assign new_n9464 = ~new_n8327 & ~new_n9463 ;
  assign new_n9465 = ~new_n8428 & ~new_n9461 ;
  assign new_n9466 = new_n8327 & new_n9465 ;
  assign new_n9467 = ~new_n9464 & ~new_n9466 ;
  assign new_n9468 = new_n8298 & ~new_n9467 ;
  assign new_n9469 = new_n8298 & ~new_n9468 ;
  assign new_n9470 = ~new_n8195 & ~new_n9469 ;
  assign new_n9471 = ~new_n8298 & ~new_n9467 ;
  assign new_n9472 = new_n8195 & new_n9471 ;
  assign new_n9473 = ~new_n9470 & ~new_n9472 ;
  assign new_n9474 = new_n8166 & ~new_n9473 ;
  assign new_n9475 = new_n8166 & ~new_n9474 ;
  assign new_n9476 = ~new_n8067 & ~new_n9475 ;
  assign new_n9477 = ~new_n8166 & ~new_n9473 ;
  assign new_n9478 = new_n8067 & new_n9477 ;
  assign new_n9479 = ~new_n9476 & ~new_n9478 ;
  assign new_n9480 = new_n8038 & ~new_n9479 ;
  assign new_n9481 = new_n8038 & ~new_n9480 ;
  assign new_n9482 = ~new_n7926 & ~new_n9481 ;
  assign new_n9483 = ~new_n8038 & ~new_n9479 ;
  assign new_n9484 = new_n7926 & new_n9483 ;
  assign new_n9485 = ~new_n9482 & ~new_n9484 ;
  assign new_n9486 = new_n7897 & ~new_n9485 ;
  assign new_n9487 = new_n7897 & ~new_n9486 ;
  assign new_n9488 = ~new_n7802 & ~new_n9487 ;
  assign new_n9489 = ~new_n7897 & ~new_n9485 ;
  assign new_n9490 = new_n7802 & new_n9489 ;
  assign new_n9491 = ~new_n9488 & ~new_n9490 ;
  assign new_n9492 = new_n7775 & ~new_n9491 ;
  assign new_n9493 = new_n7775 & ~new_n9492 ;
  assign new_n9494 = ~new_n7678 & ~new_n9493 ;
  assign new_n9495 = ~new_n7775 & ~new_n9491 ;
  assign new_n9496 = new_n7678 & new_n9495 ;
  assign new_n9497 = ~new_n9494 & ~new_n9496 ;
  assign new_n9498 = new_n7651 & ~new_n9497 ;
  assign new_n9499 = new_n7651 & ~new_n9498 ;
  assign new_n9500 = ~new_n7554 & ~new_n9499 ;
  assign new_n9501 = ~new_n7651 & ~new_n9497 ;
  assign new_n9502 = new_n7554 & new_n9501 ;
  assign new_n9503 = ~new_n9500 & ~new_n9502 ;
  assign new_n9504 = new_n7526 & ~new_n9503 ;
  assign new_n9505 = new_n7526 & ~new_n9504 ;
  assign new_n9506 = ~new_n7423 & ~new_n9505 ;
  assign new_n9507 = ~new_n7526 & ~new_n9503 ;
  assign new_n9508 = new_n7423 & new_n9507 ;
  assign new_n9509 = ~new_n9506 & ~new_n9508 ;
  assign new_n9510 = new_n7388 & ~new_n9509 ;
  assign new_n9511 = new_n7388 & ~new_n9510 ;
  assign new_n9512 = ~new_n7293 & ~new_n9511 ;
  assign new_n9513 = ~new_n7388 & ~new_n9509 ;
  assign new_n9514 = new_n7293 & new_n9513 ;
  assign new_n9515 = ~new_n9512 & ~new_n9514 ;
  assign new_n9516 = new_n7263 & ~new_n9515 ;
  assign new_n9517 = new_n7263 & ~new_n9516 ;
  assign new_n9518 = ~new_n7168 & ~new_n9517 ;
  assign new_n9519 = ~new_n7263 & ~new_n9515 ;
  assign new_n9520 = new_n7168 & new_n9519 ;
  assign new_n9521 = ~new_n9518 & ~new_n9520 ;
  assign new_n9522 = new_n7040 & ~new_n9521 ;
  assign new_n9523 = new_n7040 & ~new_n9522 ;
  assign new_n9524 = ~new_n6945 & ~new_n9523 ;
  assign new_n9525 = ~new_n7040 & ~new_n9521 ;
  assign new_n9526 = new_n6945 & new_n9525 ;
  assign new_n9527 = ~new_n9524 & ~new_n9526 ;
  assign new_n9528 = new_n6815 & ~new_n9527 ;
  assign new_n9529 = new_n6815 & ~new_n9528 ;
  assign new_n9530 = ~new_n6720 & ~new_n9529 ;
  assign new_n9531 = ~new_n6815 & ~new_n9527 ;
  assign new_n9532 = new_n6720 & new_n9531 ;
  assign new_n9533 = ~new_n9530 & ~new_n9532 ;
  assign new_n9534 = new_n6585 & ~new_n9533 ;
  assign new_n9535 = new_n6585 & ~new_n9534 ;
  assign new_n9536 = ~new_n6490 & ~new_n9535 ;
  assign new_n9537 = ~new_n6585 & ~new_n9533 ;
  assign new_n9538 = new_n6490 & new_n9537 ;
  assign new_n9539 = ~new_n9536 & ~new_n9538 ;
  assign new_n9540 = new_n6350 & ~new_n9539 ;
  assign new_n9541 = new_n6350 & ~new_n9540 ;
  assign new_n9542 = ~new_n6255 & ~new_n9541 ;
  assign new_n9543 = ~new_n6350 & ~new_n9539 ;
  assign new_n9544 = new_n6255 & new_n9543 ;
  assign new_n9545 = ~new_n9542 & ~new_n9544 ;
  assign new_n9546 = new_n6120 & ~new_n9545 ;
  assign new_n9547 = new_n6120 & ~new_n9546 ;
  assign new_n9548 = ~new_n6025 & ~new_n9547 ;
  assign new_n9549 = ~new_n6120 & ~new_n9545 ;
  assign new_n9550 = new_n6025 & new_n9549 ;
  assign new_n9551 = ~new_n9548 & ~new_n9550 ;
  assign new_n9552 = new_n5894 & ~new_n9551 ;
  assign new_n9553 = new_n5894 & ~new_n9552 ;
  assign new_n9554 = ~new_n5799 & ~new_n9553 ;
  assign new_n9555 = ~new_n5894 & ~new_n9551 ;
  assign new_n9556 = new_n5799 & new_n9555 ;
  assign new_n9557 = ~new_n9554 & ~new_n9556 ;
  assign new_n9558 = new_n5668 & ~new_n9557 ;
  assign new_n9559 = new_n5668 & ~new_n9558 ;
  assign new_n9560 = ~new_n5573 & ~new_n9559 ;
  assign new_n9561 = ~new_n5668 & ~new_n9557 ;
  assign new_n9562 = new_n5573 & new_n9561 ;
  assign new_n9563 = ~new_n9560 & ~new_n9562 ;
  assign new_n9564 = new_n5384 & ~new_n9563 ;
  assign new_n9565 = new_n5384 & ~new_n9564 ;
  assign new_n9566 = ~new_n5289 & ~new_n9565 ;
  assign new_n9567 = ~new_n5384 & ~new_n9563 ;
  assign new_n9568 = new_n5289 & new_n9567 ;
  assign new_n9569 = ~new_n9566 & ~new_n9568 ;
  assign new_n9570 = new_n5100 & ~new_n9569 ;
  assign new_n9571 = new_n5100 & ~new_n9570 ;
  assign new_n9572 = ~new_n5005 & ~new_n9571 ;
  assign new_n9573 = ~new_n5100 & ~new_n9569 ;
  assign new_n9574 = new_n5005 & new_n9573 ;
  assign new_n9575 = ~new_n9572 & ~new_n9574 ;
  assign new_n9576 = new_n4738 & ~new_n9575 ;
  assign new_n9577 = new_n4738 & ~new_n9576 ;
  assign new_n9578 = ~new_n4643 & ~new_n9577 ;
  assign new_n9579 = ~new_n4738 & ~new_n9575 ;
  assign new_n9580 = new_n4643 & new_n9579 ;
  assign new_n9581 = ~new_n9578 & ~new_n9580 ;
  assign new_n9582 = new_n4376 & ~new_n9581 ;
  assign new_n9583 = new_n4376 & ~new_n9582 ;
  assign new_n9584 = ~new_n4281 & ~new_n9583 ;
  assign new_n9585 = ~new_n4376 & ~new_n9581 ;
  assign new_n9586 = new_n4281 & new_n9585 ;
  assign new_n9587 = ~new_n9584 & ~new_n9586 ;
  assign new_n9588 = new_n4017 & ~new_n9587 ;
  assign new_n9589 = new_n4017 & ~new_n9588 ;
  assign new_n9590 = ~new_n3922 & ~new_n9589 ;
  assign new_n9591 = ~new_n4017 & ~new_n9587 ;
  assign new_n9592 = new_n3922 & new_n9591 ;
  assign new_n9593 = ~new_n9590 & ~new_n9592 ;
  assign new_n9594 = new_n3653 & ~new_n9593 ;
  assign new_n9595 = new_n3653 & ~new_n9594 ;
  assign new_n9596 = ~new_n3557 & ~new_n9595 ;
  assign new_n9597 = ~new_n3653 & ~new_n9593 ;
  assign new_n9598 = new_n3557 & new_n9597 ;
  assign new_n9599 = ~new_n9596 & ~new_n9598 ;
  assign new_n9600 = ~new_n3295 & ~new_n9599 ;
  assign new_n9601 = new_n3295 & new_n9599 ;
  assign new_n9602 = ~new_n9600 & ~new_n9601 ;
  assign new_n9603 = ~new_n3105 & ~new_n9602 ;
  assign new_n9604 = new_n3295 & ~new_n9599 ;
  assign new_n9605 = ~new_n3295 & new_n9599 ;
  assign new_n9606 = ~new_n9604 & ~new_n9605 ;
  assign new_n9607 = new_n3105 & ~new_n9606 ;
  assign new_n9608 = ~new_n9603 & ~new_n9607 ;
  assign new_n9609 = new_n3653 & new_n9593 ;
  assign new_n9610 = ~new_n9597 & ~new_n9609 ;
  assign new_n9611 = ~new_n3557 & ~new_n9610 ;
  assign new_n9612 = ~new_n3653 & new_n9593 ;
  assign new_n9613 = ~new_n9594 & ~new_n9612 ;
  assign new_n9614 = new_n3557 & ~new_n9613 ;
  assign new_n9615 = ~new_n9611 & ~new_n9614 ;
  assign new_n9616 = new_n4017 & new_n9587 ;
  assign new_n9617 = ~new_n9591 & ~new_n9616 ;
  assign new_n9618 = ~new_n3922 & ~new_n9617 ;
  assign new_n9619 = ~new_n4017 & new_n9587 ;
  assign new_n9620 = ~new_n9588 & ~new_n9619 ;
  assign new_n9621 = new_n3922 & ~new_n9620 ;
  assign new_n9622 = ~new_n9618 & ~new_n9621 ;
  assign new_n9623 = new_n4376 & new_n9581 ;
  assign new_n9624 = ~new_n9585 & ~new_n9623 ;
  assign new_n9625 = ~new_n4281 & ~new_n9624 ;
  assign new_n9626 = ~new_n4376 & new_n9581 ;
  assign new_n9627 = ~new_n9582 & ~new_n9626 ;
  assign new_n9628 = new_n4281 & ~new_n9627 ;
  assign new_n9629 = ~new_n9625 & ~new_n9628 ;
  assign new_n9630 = new_n4738 & new_n9575 ;
  assign new_n9631 = ~new_n9579 & ~new_n9630 ;
  assign new_n9632 = ~new_n4643 & ~new_n9631 ;
  assign new_n9633 = ~new_n4738 & new_n9575 ;
  assign new_n9634 = ~new_n9576 & ~new_n9633 ;
  assign new_n9635 = new_n4643 & ~new_n9634 ;
  assign new_n9636 = ~new_n9632 & ~new_n9635 ;
  assign new_n9637 = new_n5100 & new_n9569 ;
  assign new_n9638 = ~new_n9573 & ~new_n9637 ;
  assign new_n9639 = ~new_n5005 & ~new_n9638 ;
  assign new_n9640 = ~new_n5100 & new_n9569 ;
  assign new_n9641 = ~new_n9570 & ~new_n9640 ;
  assign new_n9642 = new_n5005 & ~new_n9641 ;
  assign new_n9643 = ~new_n9639 & ~new_n9642 ;
  assign new_n9644 = new_n5384 & new_n9563 ;
  assign new_n9645 = ~new_n9567 & ~new_n9644 ;
  assign new_n9646 = ~new_n5289 & ~new_n9645 ;
  assign new_n9647 = ~new_n5384 & new_n9563 ;
  assign new_n9648 = ~new_n9564 & ~new_n9647 ;
  assign new_n9649 = new_n5289 & ~new_n9648 ;
  assign new_n9650 = ~new_n9646 & ~new_n9649 ;
  assign new_n9651 = new_n5668 & new_n9557 ;
  assign new_n9652 = ~new_n9561 & ~new_n9651 ;
  assign new_n9653 = ~new_n5573 & ~new_n9652 ;
  assign new_n9654 = ~new_n5668 & new_n9557 ;
  assign new_n9655 = ~new_n9558 & ~new_n9654 ;
  assign new_n9656 = new_n5573 & ~new_n9655 ;
  assign new_n9657 = ~new_n9653 & ~new_n9656 ;
  assign new_n9658 = new_n5894 & new_n9551 ;
  assign new_n9659 = ~new_n9555 & ~new_n9658 ;
  assign new_n9660 = ~new_n5799 & ~new_n9659 ;
  assign new_n9661 = ~new_n5894 & new_n9551 ;
  assign new_n9662 = ~new_n9552 & ~new_n9661 ;
  assign new_n9663 = new_n5799 & ~new_n9662 ;
  assign new_n9664 = ~new_n9660 & ~new_n9663 ;
  assign new_n9665 = new_n6120 & new_n9545 ;
  assign new_n9666 = ~new_n9549 & ~new_n9665 ;
  assign new_n9667 = ~new_n6025 & ~new_n9666 ;
  assign new_n9668 = ~new_n6120 & new_n9545 ;
  assign new_n9669 = ~new_n9546 & ~new_n9668 ;
  assign new_n9670 = new_n6025 & ~new_n9669 ;
  assign new_n9671 = ~new_n9667 & ~new_n9670 ;
  assign new_n9672 = new_n6350 & new_n9539 ;
  assign new_n9673 = ~new_n9543 & ~new_n9672 ;
  assign new_n9674 = ~new_n6255 & ~new_n9673 ;
  assign new_n9675 = ~new_n6350 & new_n9539 ;
  assign new_n9676 = ~new_n9540 & ~new_n9675 ;
  assign new_n9677 = new_n6255 & ~new_n9676 ;
  assign new_n9678 = ~new_n9674 & ~new_n9677 ;
  assign new_n9679 = new_n6585 & new_n9533 ;
  assign new_n9680 = ~new_n9537 & ~new_n9679 ;
  assign new_n9681 = ~new_n6490 & ~new_n9680 ;
  assign new_n9682 = ~new_n6585 & new_n9533 ;
  assign new_n9683 = ~new_n9534 & ~new_n9682 ;
  assign new_n9684 = new_n6490 & ~new_n9683 ;
  assign new_n9685 = ~new_n9681 & ~new_n9684 ;
  assign new_n9686 = new_n6815 & new_n9527 ;
  assign new_n9687 = ~new_n9531 & ~new_n9686 ;
  assign new_n9688 = ~new_n6720 & ~new_n9687 ;
  assign new_n9689 = ~new_n6815 & new_n9527 ;
  assign new_n9690 = ~new_n9528 & ~new_n9689 ;
  assign new_n9691 = new_n6720 & ~new_n9690 ;
  assign new_n9692 = ~new_n9688 & ~new_n9691 ;
  assign new_n9693 = new_n7040 & new_n9521 ;
  assign new_n9694 = ~new_n9525 & ~new_n9693 ;
  assign new_n9695 = ~new_n6945 & ~new_n9694 ;
  assign new_n9696 = ~new_n7040 & new_n9521 ;
  assign new_n9697 = ~new_n9522 & ~new_n9696 ;
  assign new_n9698 = new_n6945 & ~new_n9697 ;
  assign new_n9699 = ~new_n9695 & ~new_n9698 ;
  assign new_n9700 = new_n7263 & new_n9515 ;
  assign new_n9701 = ~new_n9519 & ~new_n9700 ;
  assign new_n9702 = ~new_n7168 & ~new_n9701 ;
  assign new_n9703 = ~new_n7263 & new_n9515 ;
  assign new_n9704 = ~new_n9516 & ~new_n9703 ;
  assign new_n9705 = new_n7168 & ~new_n9704 ;
  assign new_n9706 = ~new_n9702 & ~new_n9705 ;
  assign new_n9707 = new_n7388 & new_n9509 ;
  assign new_n9708 = ~new_n9513 & ~new_n9707 ;
  assign new_n9709 = ~new_n7293 & ~new_n9708 ;
  assign new_n9710 = ~new_n7388 & new_n9509 ;
  assign new_n9711 = ~new_n9510 & ~new_n9710 ;
  assign new_n9712 = new_n7293 & ~new_n9711 ;
  assign new_n9713 = ~new_n9709 & ~new_n9712 ;
  assign new_n9714 = new_n7526 & new_n9503 ;
  assign new_n9715 = ~new_n9507 & ~new_n9714 ;
  assign new_n9716 = ~new_n7423 & ~new_n9715 ;
  assign new_n9717 = ~new_n7526 & new_n9503 ;
  assign new_n9718 = ~new_n9504 & ~new_n9717 ;
  assign new_n9719 = new_n7423 & ~new_n9718 ;
  assign new_n9720 = ~new_n9716 & ~new_n9719 ;
  assign new_n9721 = new_n7651 & new_n9497 ;
  assign new_n9722 = ~new_n9501 & ~new_n9721 ;
  assign new_n9723 = ~new_n7554 & ~new_n9722 ;
  assign new_n9724 = ~new_n7651 & new_n9497 ;
  assign new_n9725 = ~new_n9498 & ~new_n9724 ;
  assign new_n9726 = new_n7554 & ~new_n9725 ;
  assign new_n9727 = ~new_n9723 & ~new_n9726 ;
  assign new_n9728 = new_n7775 & new_n9491 ;
  assign new_n9729 = ~new_n9495 & ~new_n9728 ;
  assign new_n9730 = ~new_n7678 & ~new_n9729 ;
  assign new_n9731 = ~new_n7775 & new_n9491 ;
  assign new_n9732 = ~new_n9492 & ~new_n9731 ;
  assign new_n9733 = new_n7678 & ~new_n9732 ;
  assign new_n9734 = ~new_n9730 & ~new_n9733 ;
  assign new_n9735 = new_n7897 & new_n9485 ;
  assign new_n9736 = ~new_n9489 & ~new_n9735 ;
  assign new_n9737 = ~new_n7802 & ~new_n9736 ;
  assign new_n9738 = ~new_n7897 & new_n9485 ;
  assign new_n9739 = ~new_n9486 & ~new_n9738 ;
  assign new_n9740 = new_n7802 & ~new_n9739 ;
  assign new_n9741 = ~new_n9737 & ~new_n9740 ;
  assign new_n9742 = new_n8038 & new_n9479 ;
  assign new_n9743 = ~new_n9483 & ~new_n9742 ;
  assign new_n9744 = ~new_n7926 & ~new_n9743 ;
  assign new_n9745 = ~new_n8038 & new_n9479 ;
  assign new_n9746 = ~new_n9480 & ~new_n9745 ;
  assign new_n9747 = new_n7926 & ~new_n9746 ;
  assign new_n9748 = ~new_n9744 & ~new_n9747 ;
  assign new_n9749 = new_n8166 & new_n9473 ;
  assign new_n9750 = ~new_n9477 & ~new_n9749 ;
  assign new_n9751 = ~new_n8067 & ~new_n9750 ;
  assign new_n9752 = ~new_n8166 & new_n9473 ;
  assign new_n9753 = ~new_n9474 & ~new_n9752 ;
  assign new_n9754 = new_n8067 & ~new_n9753 ;
  assign new_n9755 = ~new_n9751 & ~new_n9754 ;
  assign new_n9756 = new_n8298 & new_n9467 ;
  assign new_n9757 = ~new_n9471 & ~new_n9756 ;
  assign new_n9758 = ~new_n8195 & ~new_n9757 ;
  assign new_n9759 = ~new_n8298 & new_n9467 ;
  assign new_n9760 = ~new_n9468 & ~new_n9759 ;
  assign new_n9761 = new_n8195 & ~new_n9760 ;
  assign new_n9762 = ~new_n9758 & ~new_n9761 ;
  assign new_n9763 = new_n8428 & new_n9461 ;
  assign new_n9764 = ~new_n9465 & ~new_n9763 ;
  assign new_n9765 = ~new_n8327 & ~new_n9764 ;
  assign new_n9766 = ~new_n8428 & new_n9461 ;
  assign new_n9767 = ~new_n9462 & ~new_n9766 ;
  assign new_n9768 = new_n8327 & ~new_n9767 ;
  assign new_n9769 = ~new_n9765 & ~new_n9768 ;
  assign new_n9770 = new_n8554 & new_n9455 ;
  assign new_n9771 = ~new_n9459 & ~new_n9770 ;
  assign new_n9772 = ~new_n8449 & ~new_n9771 ;
  assign new_n9773 = ~new_n8554 & new_n9455 ;
  assign new_n9774 = ~new_n9456 & ~new_n9773 ;
  assign new_n9775 = new_n8449 & ~new_n9774 ;
  assign new_n9776 = ~new_n9772 & ~new_n9775 ;
  assign new_n9777 = new_n8675 & new_n9449 ;
  assign new_n9778 = ~new_n9453 & ~new_n9777 ;
  assign new_n9779 = ~new_n8575 & ~new_n9778 ;
  assign new_n9780 = ~new_n8675 & new_n9449 ;
  assign new_n9781 = ~new_n9450 & ~new_n9780 ;
  assign new_n9782 = new_n8575 & ~new_n9781 ;
  assign new_n9783 = ~new_n9779 & ~new_n9782 ;
  assign new_n9784 = new_n8797 & new_n9443 ;
  assign new_n9785 = ~new_n9447 & ~new_n9784 ;
  assign new_n9786 = ~new_n8696 & ~new_n9785 ;
  assign new_n9787 = ~new_n8797 & new_n9443 ;
  assign new_n9788 = ~new_n9444 & ~new_n9787 ;
  assign new_n9789 = new_n8696 & ~new_n9788 ;
  assign new_n9790 = ~new_n9786 & ~new_n9789 ;
  assign new_n9791 = new_n8918 & new_n9437 ;
  assign new_n9792 = ~new_n9441 & ~new_n9791 ;
  assign new_n9793 = ~new_n8818 & ~new_n9792 ;
  assign new_n9794 = ~new_n8918 & new_n9437 ;
  assign new_n9795 = ~new_n9438 & ~new_n9794 ;
  assign new_n9796 = new_n8818 & ~new_n9795 ;
  assign new_n9797 = ~new_n9793 & ~new_n9796 ;
  assign new_n9798 = new_n9038 & new_n9431 ;
  assign new_n9799 = ~new_n9435 & ~new_n9798 ;
  assign new_n9800 = ~new_n8939 & ~new_n9799 ;
  assign new_n9801 = ~new_n9038 & new_n9431 ;
  assign new_n9802 = ~new_n9432 & ~new_n9801 ;
  assign new_n9803 = new_n8939 & ~new_n9802 ;
  assign new_n9804 = ~new_n9800 & ~new_n9803 ;
  assign new_n9805 = new_n9162 & new_n9425 ;
  assign new_n9806 = ~new_n9429 & ~new_n9805 ;
  assign new_n9807 = ~new_n9059 & ~new_n9806 ;
  assign new_n9808 = ~new_n9162 & new_n9425 ;
  assign new_n9809 = ~new_n9426 & ~new_n9808 ;
  assign new_n9810 = new_n9059 & ~new_n9809 ;
  assign new_n9811 = ~new_n9807 & ~new_n9810 ;
  assign new_n9812 = new_n9286 & new_n9419 ;
  assign new_n9813 = ~new_n9423 & ~new_n9812 ;
  assign new_n9814 = ~new_n9182 & ~new_n9813 ;
  assign new_n9815 = ~new_n9286 & new_n9419 ;
  assign new_n9816 = ~new_n9420 & ~new_n9815 ;
  assign new_n9817 = new_n9182 & ~new_n9816 ;
  assign new_n9818 = ~new_n9814 & ~new_n9817 ;
  assign new_n9819 = new_n9408 & new_n9413 ;
  assign new_n9820 = ~new_n9417 & ~new_n9819 ;
  assign new_n9821 = ~new_n9305 & ~new_n9820 ;
  assign new_n9822 = ~new_n9408 & new_n9413 ;
  assign new_n9823 = ~new_n9414 & ~new_n9822 ;
  assign new_n9824 = new_n9305 & ~new_n9823 ;
  assign new_n9825 = ~new_n9821 & ~new_n9824 ;
  assign new_n9826 = new_n9303 & ~new_n9825 ;
  assign new_n9827 = new_n9818 & new_n9826 ;
  assign new_n9828 = new_n9818 & ~new_n9827 ;
  assign new_n9829 = new_n9180 & ~new_n9828 ;
  assign new_n9830 = ~new_n9180 & new_n9826 ;
  assign new_n9831 = ~new_n9818 & new_n9830 ;
  assign new_n9832 = ~new_n9829 & ~new_n9831 ;
  assign new_n9833 = new_n9811 & ~new_n9832 ;
  assign new_n9834 = new_n9811 & ~new_n9833 ;
  assign new_n9835 = new_n9056 & ~new_n9834 ;
  assign new_n9836 = ~new_n9056 & ~new_n9832 ;
  assign new_n9837 = ~new_n9811 & new_n9836 ;
  assign new_n9838 = ~new_n9835 & ~new_n9837 ;
  assign new_n9839 = new_n9804 & ~new_n9838 ;
  assign new_n9840 = new_n9804 & ~new_n9839 ;
  assign new_n9841 = new_n8936 & ~new_n9840 ;
  assign new_n9842 = ~new_n8936 & ~new_n9838 ;
  assign new_n9843 = ~new_n9804 & new_n9842 ;
  assign new_n9844 = ~new_n9841 & ~new_n9843 ;
  assign new_n9845 = new_n9797 & ~new_n9844 ;
  assign new_n9846 = new_n9797 & ~new_n9845 ;
  assign new_n9847 = new_n8815 & ~new_n9846 ;
  assign new_n9848 = ~new_n8815 & ~new_n9844 ;
  assign new_n9849 = ~new_n9797 & new_n9848 ;
  assign new_n9850 = ~new_n9847 & ~new_n9849 ;
  assign new_n9851 = new_n9790 & ~new_n9850 ;
  assign new_n9852 = new_n9790 & ~new_n9851 ;
  assign new_n9853 = new_n8693 & ~new_n9852 ;
  assign new_n9854 = ~new_n8693 & ~new_n9850 ;
  assign new_n9855 = ~new_n9790 & new_n9854 ;
  assign new_n9856 = ~new_n9853 & ~new_n9855 ;
  assign new_n9857 = new_n9783 & ~new_n9856 ;
  assign new_n9858 = new_n9783 & ~new_n9857 ;
  assign new_n9859 = new_n8572 & ~new_n9858 ;
  assign new_n9860 = ~new_n8572 & ~new_n9856 ;
  assign new_n9861 = ~new_n9783 & new_n9860 ;
  assign new_n9862 = ~new_n9859 & ~new_n9861 ;
  assign new_n9863 = new_n9776 & ~new_n9862 ;
  assign new_n9864 = new_n9776 & ~new_n9863 ;
  assign new_n9865 = new_n8446 & ~new_n9864 ;
  assign new_n9866 = ~new_n8446 & ~new_n9862 ;
  assign new_n9867 = ~new_n9776 & new_n9866 ;
  assign new_n9868 = ~new_n9865 & ~new_n9867 ;
  assign new_n9869 = new_n9769 & ~new_n9868 ;
  assign new_n9870 = new_n9769 & ~new_n9869 ;
  assign new_n9871 = new_n8324 & ~new_n9870 ;
  assign new_n9872 = ~new_n8324 & ~new_n9868 ;
  assign new_n9873 = ~new_n9769 & new_n9872 ;
  assign new_n9874 = ~new_n9871 & ~new_n9873 ;
  assign new_n9875 = new_n9762 & ~new_n9874 ;
  assign new_n9876 = new_n9762 & ~new_n9875 ;
  assign new_n9877 = new_n8192 & ~new_n9876 ;
  assign new_n9878 = ~new_n8192 & ~new_n9874 ;
  assign new_n9879 = ~new_n9762 & new_n9878 ;
  assign new_n9880 = ~new_n9877 & ~new_n9879 ;
  assign new_n9881 = new_n9755 & ~new_n9880 ;
  assign new_n9882 = new_n9755 & ~new_n9881 ;
  assign new_n9883 = new_n8064 & ~new_n9882 ;
  assign new_n9884 = ~new_n8064 & ~new_n9880 ;
  assign new_n9885 = ~new_n9755 & new_n9884 ;
  assign new_n9886 = ~new_n9883 & ~new_n9885 ;
  assign new_n9887 = new_n9748 & ~new_n9886 ;
  assign new_n9888 = new_n9748 & ~new_n9887 ;
  assign new_n9889 = new_n7923 & ~new_n9888 ;
  assign new_n9890 = ~new_n7923 & ~new_n9886 ;
  assign new_n9891 = ~new_n9748 & new_n9890 ;
  assign new_n9892 = ~new_n9889 & ~new_n9891 ;
  assign new_n9893 = new_n9741 & ~new_n9892 ;
  assign new_n9894 = new_n9741 & ~new_n9893 ;
  assign new_n9895 = new_n7799 & ~new_n9894 ;
  assign new_n9896 = ~new_n7799 & ~new_n9892 ;
  assign new_n9897 = ~new_n9741 & new_n9896 ;
  assign new_n9898 = ~new_n9895 & ~new_n9897 ;
  assign new_n9899 = new_n9734 & ~new_n9898 ;
  assign new_n9900 = new_n9734 & ~new_n9899 ;
  assign new_n9901 = new_n7675 & ~new_n9900 ;
  assign new_n9902 = ~new_n7675 & ~new_n9898 ;
  assign new_n9903 = ~new_n9734 & new_n9902 ;
  assign new_n9904 = ~new_n9901 & ~new_n9903 ;
  assign new_n9905 = new_n9727 & ~new_n9904 ;
  assign new_n9906 = new_n9727 & ~new_n9905 ;
  assign new_n9907 = new_n7551 & ~new_n9906 ;
  assign new_n9908 = ~new_n7551 & ~new_n9904 ;
  assign new_n9909 = ~new_n9727 & new_n9908 ;
  assign new_n9910 = ~new_n9907 & ~new_n9909 ;
  assign new_n9911 = new_n9720 & ~new_n9910 ;
  assign new_n9912 = new_n9720 & ~new_n9911 ;
  assign new_n9913 = new_n7420 & ~new_n9912 ;
  assign new_n9914 = ~new_n7420 & ~new_n9910 ;
  assign new_n9915 = ~new_n9720 & new_n9914 ;
  assign new_n9916 = ~new_n9913 & ~new_n9915 ;
  assign new_n9917 = new_n9713 & ~new_n9916 ;
  assign new_n9918 = new_n9713 & ~new_n9917 ;
  assign new_n9919 = new_n7290 & ~new_n9918 ;
  assign new_n9920 = ~new_n7290 & ~new_n9916 ;
  assign new_n9921 = ~new_n9713 & new_n9920 ;
  assign new_n9922 = ~new_n9919 & ~new_n9921 ;
  assign new_n9923 = new_n9706 & ~new_n9922 ;
  assign new_n9924 = new_n9706 & ~new_n9923 ;
  assign new_n9925 = new_n7165 & ~new_n9924 ;
  assign new_n9926 = ~new_n7165 & ~new_n9922 ;
  assign new_n9927 = ~new_n9706 & new_n9926 ;
  assign new_n9928 = ~new_n9925 & ~new_n9927 ;
  assign new_n9929 = new_n9699 & ~new_n9928 ;
  assign new_n9930 = new_n9699 & ~new_n9929 ;
  assign new_n9931 = new_n6942 & ~new_n9930 ;
  assign new_n9932 = ~new_n6942 & ~new_n9928 ;
  assign new_n9933 = ~new_n9699 & new_n9932 ;
  assign new_n9934 = ~new_n9931 & ~new_n9933 ;
  assign new_n9935 = new_n9692 & ~new_n9934 ;
  assign new_n9936 = new_n9692 & ~new_n9935 ;
  assign new_n9937 = new_n6717 & ~new_n9936 ;
  assign new_n9938 = ~new_n6717 & ~new_n9934 ;
  assign new_n9939 = ~new_n9692 & new_n9938 ;
  assign new_n9940 = ~new_n9937 & ~new_n9939 ;
  assign new_n9941 = new_n9685 & ~new_n9940 ;
  assign new_n9942 = new_n9685 & ~new_n9941 ;
  assign new_n9943 = new_n6487 & ~new_n9942 ;
  assign new_n9944 = ~new_n6487 & ~new_n9940 ;
  assign new_n9945 = ~new_n9685 & new_n9944 ;
  assign new_n9946 = ~new_n9943 & ~new_n9945 ;
  assign new_n9947 = new_n9678 & ~new_n9946 ;
  assign new_n9948 = new_n9678 & ~new_n9947 ;
  assign new_n9949 = new_n6252 & ~new_n9948 ;
  assign new_n9950 = ~new_n6252 & ~new_n9946 ;
  assign new_n9951 = ~new_n9678 & new_n9950 ;
  assign new_n9952 = ~new_n9949 & ~new_n9951 ;
  assign new_n9953 = new_n9671 & ~new_n9952 ;
  assign new_n9954 = new_n9671 & ~new_n9953 ;
  assign new_n9955 = new_n6022 & ~new_n9954 ;
  assign new_n9956 = ~new_n6022 & ~new_n9952 ;
  assign new_n9957 = ~new_n9671 & new_n9956 ;
  assign new_n9958 = ~new_n9955 & ~new_n9957 ;
  assign new_n9959 = new_n9664 & ~new_n9958 ;
  assign new_n9960 = new_n9664 & ~new_n9959 ;
  assign new_n9961 = new_n5796 & ~new_n9960 ;
  assign new_n9962 = ~new_n5796 & ~new_n9958 ;
  assign new_n9963 = ~new_n9664 & new_n9962 ;
  assign new_n9964 = ~new_n9961 & ~new_n9963 ;
  assign new_n9965 = new_n9657 & ~new_n9964 ;
  assign new_n9966 = new_n9657 & ~new_n9965 ;
  assign new_n9967 = new_n5570 & ~new_n9966 ;
  assign new_n9968 = ~new_n5570 & ~new_n9964 ;
  assign new_n9969 = ~new_n9657 & new_n9968 ;
  assign new_n9970 = ~new_n9967 & ~new_n9969 ;
  assign new_n9971 = new_n9650 & ~new_n9970 ;
  assign new_n9972 = new_n9650 & ~new_n9971 ;
  assign new_n9973 = new_n5286 & ~new_n9972 ;
  assign new_n9974 = ~new_n5286 & ~new_n9970 ;
  assign new_n9975 = ~new_n9650 & new_n9974 ;
  assign new_n9976 = ~new_n9973 & ~new_n9975 ;
  assign new_n9977 = new_n9643 & ~new_n9976 ;
  assign new_n9978 = new_n9643 & ~new_n9977 ;
  assign new_n9979 = new_n5002 & ~new_n9978 ;
  assign new_n9980 = ~new_n5002 & ~new_n9976 ;
  assign new_n9981 = ~new_n9643 & new_n9980 ;
  assign new_n9982 = ~new_n9979 & ~new_n9981 ;
  assign new_n9983 = new_n9636 & ~new_n9982 ;
  assign new_n9984 = new_n9636 & ~new_n9983 ;
  assign new_n9985 = new_n4640 & ~new_n9984 ;
  assign new_n9986 = ~new_n4640 & ~new_n9982 ;
  assign new_n9987 = ~new_n9636 & new_n9986 ;
  assign new_n9988 = ~new_n9985 & ~new_n9987 ;
  assign new_n9989 = new_n9629 & ~new_n9988 ;
  assign new_n9990 = new_n9629 & ~new_n9989 ;
  assign new_n9991 = new_n4278 & ~new_n9990 ;
  assign new_n9992 = ~new_n4278 & ~new_n9988 ;
  assign new_n9993 = ~new_n9629 & new_n9992 ;
  assign new_n9994 = ~new_n9991 & ~new_n9993 ;
  assign new_n9995 = new_n9622 & ~new_n9994 ;
  assign new_n9996 = new_n9622 & ~new_n9995 ;
  assign new_n9997 = new_n3919 & ~new_n9996 ;
  assign new_n9998 = ~new_n3919 & ~new_n9994 ;
  assign new_n9999 = ~new_n9622 & new_n9998 ;
  assign new_n10000 = ~new_n9997 & ~new_n9999 ;
  assign new_n10001 = new_n9615 & ~new_n10000 ;
  assign new_n10002 = new_n9615 & ~new_n10001 ;
  assign new_n10003 = new_n3554 & ~new_n10002 ;
  assign new_n10004 = ~new_n3554 & ~new_n10000 ;
  assign new_n10005 = ~new_n9615 & new_n10004 ;
  assign new_n10006 = ~new_n10003 & ~new_n10005 ;
  assign new_n10007 = new_n9608 & ~new_n10006 ;
  assign new_n10008 = new_n9608 & ~new_n10007 ;
  assign new_n10009 = new_n3098 & ~new_n10008 ;
  assign new_n10010 = ~new_n3098 & ~new_n10006 ;
  assign new_n10011 = ~new_n9608 & new_n10010 ;
  assign new_n10012 = ~new_n10009 & ~new_n10011 ;
  assign new_n10013 = ~lo0826 & ~new_n10012 ;
  assign new_n10014 = ~new_n9303 & new_n9825 ;
  assign new_n10015 = new_n9180 & new_n10014 ;
  assign new_n10016 = new_n9180 & ~new_n10015 ;
  assign new_n10017 = new_n9818 & ~new_n10016 ;
  assign new_n10018 = ~new_n9180 & new_n10014 ;
  assign new_n10019 = ~new_n9818 & new_n10018 ;
  assign new_n10020 = ~new_n10017 & ~new_n10019 ;
  assign new_n10021 = new_n9056 & ~new_n10020 ;
  assign new_n10022 = new_n9056 & ~new_n10021 ;
  assign new_n10023 = new_n9811 & ~new_n10022 ;
  assign new_n10024 = ~new_n9056 & ~new_n10020 ;
  assign new_n10025 = ~new_n9811 & new_n10024 ;
  assign new_n10026 = ~new_n10023 & ~new_n10025 ;
  assign new_n10027 = new_n8936 & ~new_n10026 ;
  assign new_n10028 = new_n8936 & ~new_n10027 ;
  assign new_n10029 = new_n9804 & ~new_n10028 ;
  assign new_n10030 = ~new_n8936 & ~new_n10026 ;
  assign new_n10031 = ~new_n9804 & new_n10030 ;
  assign new_n10032 = ~new_n10029 & ~new_n10031 ;
  assign new_n10033 = new_n8815 & ~new_n10032 ;
  assign new_n10034 = new_n8815 & ~new_n10033 ;
  assign new_n10035 = new_n9797 & ~new_n10034 ;
  assign new_n10036 = ~new_n8815 & ~new_n10032 ;
  assign new_n10037 = ~new_n9797 & new_n10036 ;
  assign new_n10038 = ~new_n10035 & ~new_n10037 ;
  assign new_n10039 = new_n8693 & ~new_n10038 ;
  assign new_n10040 = new_n8693 & ~new_n10039 ;
  assign new_n10041 = new_n9790 & ~new_n10040 ;
  assign new_n10042 = ~new_n8693 & ~new_n10038 ;
  assign new_n10043 = ~new_n9790 & new_n10042 ;
  assign new_n10044 = ~new_n10041 & ~new_n10043 ;
  assign new_n10045 = new_n8572 & ~new_n10044 ;
  assign new_n10046 = new_n8572 & ~new_n10045 ;
  assign new_n10047 = new_n9783 & ~new_n10046 ;
  assign new_n10048 = ~new_n8572 & ~new_n10044 ;
  assign new_n10049 = ~new_n9783 & new_n10048 ;
  assign new_n10050 = ~new_n10047 & ~new_n10049 ;
  assign new_n10051 = new_n8446 & ~new_n10050 ;
  assign new_n10052 = new_n8446 & ~new_n10051 ;
  assign new_n10053 = new_n9776 & ~new_n10052 ;
  assign new_n10054 = ~new_n8446 & ~new_n10050 ;
  assign new_n10055 = ~new_n9776 & new_n10054 ;
  assign new_n10056 = ~new_n10053 & ~new_n10055 ;
  assign new_n10057 = new_n8324 & ~new_n10056 ;
  assign new_n10058 = new_n8324 & ~new_n10057 ;
  assign new_n10059 = new_n9769 & ~new_n10058 ;
  assign new_n10060 = ~new_n8324 & ~new_n10056 ;
  assign new_n10061 = ~new_n9769 & new_n10060 ;
  assign new_n10062 = ~new_n10059 & ~new_n10061 ;
  assign new_n10063 = new_n8192 & ~new_n10062 ;
  assign new_n10064 = new_n8192 & ~new_n10063 ;
  assign new_n10065 = new_n9762 & ~new_n10064 ;
  assign new_n10066 = ~new_n8192 & ~new_n10062 ;
  assign new_n10067 = ~new_n9762 & new_n10066 ;
  assign new_n10068 = ~new_n10065 & ~new_n10067 ;
  assign new_n10069 = new_n8064 & ~new_n10068 ;
  assign new_n10070 = new_n8064 & ~new_n10069 ;
  assign new_n10071 = new_n9755 & ~new_n10070 ;
  assign new_n10072 = ~new_n8064 & ~new_n10068 ;
  assign new_n10073 = ~new_n9755 & new_n10072 ;
  assign new_n10074 = ~new_n10071 & ~new_n10073 ;
  assign new_n10075 = new_n7923 & ~new_n10074 ;
  assign new_n10076 = new_n7923 & ~new_n10075 ;
  assign new_n10077 = new_n9748 & ~new_n10076 ;
  assign new_n10078 = ~new_n7923 & ~new_n10074 ;
  assign new_n10079 = ~new_n9748 & new_n10078 ;
  assign new_n10080 = ~new_n10077 & ~new_n10079 ;
  assign new_n10081 = new_n7799 & ~new_n10080 ;
  assign new_n10082 = new_n7799 & ~new_n10081 ;
  assign new_n10083 = new_n9741 & ~new_n10082 ;
  assign new_n10084 = ~new_n7799 & ~new_n10080 ;
  assign new_n10085 = ~new_n9741 & new_n10084 ;
  assign new_n10086 = ~new_n10083 & ~new_n10085 ;
  assign new_n10087 = new_n7675 & ~new_n10086 ;
  assign new_n10088 = new_n7675 & ~new_n10087 ;
  assign new_n10089 = new_n9734 & ~new_n10088 ;
  assign new_n10090 = ~new_n7675 & ~new_n10086 ;
  assign new_n10091 = ~new_n9734 & new_n10090 ;
  assign new_n10092 = ~new_n10089 & ~new_n10091 ;
  assign new_n10093 = new_n7551 & ~new_n10092 ;
  assign new_n10094 = new_n7551 & ~new_n10093 ;
  assign new_n10095 = new_n9727 & ~new_n10094 ;
  assign new_n10096 = ~new_n7551 & ~new_n10092 ;
  assign new_n10097 = ~new_n9727 & new_n10096 ;
  assign new_n10098 = ~new_n10095 & ~new_n10097 ;
  assign new_n10099 = new_n7420 & ~new_n10098 ;
  assign new_n10100 = new_n7420 & ~new_n10099 ;
  assign new_n10101 = new_n9720 & ~new_n10100 ;
  assign new_n10102 = ~new_n7420 & ~new_n10098 ;
  assign new_n10103 = ~new_n9720 & new_n10102 ;
  assign new_n10104 = ~new_n10101 & ~new_n10103 ;
  assign new_n10105 = new_n7290 & ~new_n10104 ;
  assign new_n10106 = new_n7290 & ~new_n10105 ;
  assign new_n10107 = new_n9713 & ~new_n10106 ;
  assign new_n10108 = ~new_n7290 & ~new_n10104 ;
  assign new_n10109 = ~new_n9713 & new_n10108 ;
  assign new_n10110 = ~new_n10107 & ~new_n10109 ;
  assign new_n10111 = new_n7165 & ~new_n10110 ;
  assign new_n10112 = new_n7165 & ~new_n10111 ;
  assign new_n10113 = new_n9706 & ~new_n10112 ;
  assign new_n10114 = ~new_n7165 & ~new_n10110 ;
  assign new_n10115 = ~new_n9706 & new_n10114 ;
  assign new_n10116 = ~new_n10113 & ~new_n10115 ;
  assign new_n10117 = new_n6942 & ~new_n10116 ;
  assign new_n10118 = new_n6942 & ~new_n10117 ;
  assign new_n10119 = new_n9699 & ~new_n10118 ;
  assign new_n10120 = ~new_n6942 & ~new_n10116 ;
  assign new_n10121 = ~new_n9699 & new_n10120 ;
  assign new_n10122 = ~new_n10119 & ~new_n10121 ;
  assign new_n10123 = new_n6717 & ~new_n10122 ;
  assign new_n10124 = new_n6717 & ~new_n10123 ;
  assign new_n10125 = new_n9692 & ~new_n10124 ;
  assign new_n10126 = ~new_n6717 & ~new_n10122 ;
  assign new_n10127 = ~new_n9692 & new_n10126 ;
  assign new_n10128 = ~new_n10125 & ~new_n10127 ;
  assign new_n10129 = new_n6487 & ~new_n10128 ;
  assign new_n10130 = new_n6487 & ~new_n10129 ;
  assign new_n10131 = new_n9685 & ~new_n10130 ;
  assign new_n10132 = ~new_n6487 & ~new_n10128 ;
  assign new_n10133 = ~new_n9685 & new_n10132 ;
  assign new_n10134 = ~new_n10131 & ~new_n10133 ;
  assign new_n10135 = new_n6252 & ~new_n10134 ;
  assign new_n10136 = new_n6252 & ~new_n10135 ;
  assign new_n10137 = new_n9678 & ~new_n10136 ;
  assign new_n10138 = ~new_n6252 & ~new_n10134 ;
  assign new_n10139 = ~new_n9678 & new_n10138 ;
  assign new_n10140 = ~new_n10137 & ~new_n10139 ;
  assign new_n10141 = new_n6022 & ~new_n10140 ;
  assign new_n10142 = new_n6022 & ~new_n10141 ;
  assign new_n10143 = new_n9671 & ~new_n10142 ;
  assign new_n10144 = ~new_n6022 & ~new_n10140 ;
  assign new_n10145 = ~new_n9671 & new_n10144 ;
  assign new_n10146 = ~new_n10143 & ~new_n10145 ;
  assign new_n10147 = new_n5796 & ~new_n10146 ;
  assign new_n10148 = new_n5796 & ~new_n10147 ;
  assign new_n10149 = new_n9664 & ~new_n10148 ;
  assign new_n10150 = ~new_n5796 & ~new_n10146 ;
  assign new_n10151 = ~new_n9664 & new_n10150 ;
  assign new_n10152 = ~new_n10149 & ~new_n10151 ;
  assign new_n10153 = new_n5570 & ~new_n10152 ;
  assign new_n10154 = new_n5570 & ~new_n10153 ;
  assign new_n10155 = new_n9657 & ~new_n10154 ;
  assign new_n10156 = ~new_n5570 & ~new_n10152 ;
  assign new_n10157 = ~new_n9657 & new_n10156 ;
  assign new_n10158 = ~new_n10155 & ~new_n10157 ;
  assign new_n10159 = new_n5286 & ~new_n10158 ;
  assign new_n10160 = new_n5286 & ~new_n10159 ;
  assign new_n10161 = new_n9650 & ~new_n10160 ;
  assign new_n10162 = ~new_n5286 & ~new_n10158 ;
  assign new_n10163 = ~new_n9650 & new_n10162 ;
  assign new_n10164 = ~new_n10161 & ~new_n10163 ;
  assign new_n10165 = new_n5002 & ~new_n10164 ;
  assign new_n10166 = new_n5002 & ~new_n10165 ;
  assign new_n10167 = new_n9643 & ~new_n10166 ;
  assign new_n10168 = ~new_n5002 & ~new_n10164 ;
  assign new_n10169 = ~new_n9643 & new_n10168 ;
  assign new_n10170 = ~new_n10167 & ~new_n10169 ;
  assign new_n10171 = new_n4640 & ~new_n10170 ;
  assign new_n10172 = new_n4640 & ~new_n10171 ;
  assign new_n10173 = new_n9636 & ~new_n10172 ;
  assign new_n10174 = ~new_n4640 & ~new_n10170 ;
  assign new_n10175 = ~new_n9636 & new_n10174 ;
  assign new_n10176 = ~new_n10173 & ~new_n10175 ;
  assign new_n10177 = new_n4278 & ~new_n10176 ;
  assign new_n10178 = new_n4278 & ~new_n10177 ;
  assign new_n10179 = new_n9629 & ~new_n10178 ;
  assign new_n10180 = ~new_n4278 & ~new_n10176 ;
  assign new_n10181 = ~new_n9629 & new_n10180 ;
  assign new_n10182 = ~new_n10179 & ~new_n10181 ;
  assign new_n10183 = new_n3919 & ~new_n10182 ;
  assign new_n10184 = new_n3919 & ~new_n10183 ;
  assign new_n10185 = new_n9622 & ~new_n10184 ;
  assign new_n10186 = ~new_n3919 & ~new_n10182 ;
  assign new_n10187 = ~new_n9622 & new_n10186 ;
  assign new_n10188 = ~new_n10185 & ~new_n10187 ;
  assign new_n10189 = new_n3554 & ~new_n10188 ;
  assign new_n10190 = new_n3554 & ~new_n10189 ;
  assign new_n10191 = new_n9615 & ~new_n10190 ;
  assign new_n10192 = ~new_n3554 & ~new_n10188 ;
  assign new_n10193 = ~new_n9615 & new_n10192 ;
  assign new_n10194 = ~new_n10191 & ~new_n10193 ;
  assign new_n10195 = new_n3098 & ~new_n10194 ;
  assign new_n10196 = new_n3098 & ~new_n10195 ;
  assign new_n10197 = new_n9608 & ~new_n10196 ;
  assign new_n10198 = ~new_n3098 & ~new_n10194 ;
  assign new_n10199 = ~new_n9608 & new_n10198 ;
  assign new_n10200 = ~new_n10197 & ~new_n10199 ;
  assign new_n10201 = lo0826 & new_n10200 ;
  assign new_n10202 = ~new_n10013 & ~new_n10201 ;
  assign new_n10203 = ~lo0110 & ~new_n10202 ;
  assign new_n10204 = ~lo0826 & ~new_n10200 ;
  assign new_n10205 = lo0826 & new_n10012 ;
  assign new_n10206 = ~new_n10204 & ~new_n10205 ;
  assign new_n10207 = lo0110 & ~new_n10206 ;
  assign new_n10208 = ~new_n10203 & ~new_n10207 ;
  assign new_n10209 = new_n2739 & ~new_n10208 ;
  assign new_n10210 = ~lo0826 & new_n10012 ;
  assign new_n10211 = lo0826 & ~new_n10200 ;
  assign new_n10212 = ~new_n10210 & ~new_n10211 ;
  assign new_n10213 = ~lo0110 & ~new_n10212 ;
  assign new_n10214 = ~lo0826 & new_n10200 ;
  assign new_n10215 = lo0826 & ~new_n10012 ;
  assign new_n10216 = ~new_n10214 & ~new_n10215 ;
  assign new_n10217 = lo0110 & ~new_n10216 ;
  assign new_n10218 = ~new_n10213 & ~new_n10217 ;
  assign new_n10219 = ~new_n2739 & ~new_n10218 ;
  assign new_n10220 = ~new_n10209 & ~new_n10219 ;
  assign new_n10221 = lo0826 & new_n10220 ;
  assign new_n10222 = ~lo0826 & ~new_n10220 ;
  assign new_n10223 = lo0854 & ~new_n10222 ;
  assign new_n10224 = ~new_n10221 & new_n10223 ;
  assign new_n10225 = ~new_n2739 & new_n3281 ;
  assign new_n10226 = new_n2739 & ~new_n3281 ;
  assign new_n10227 = ~new_n10225 & ~new_n10226 ;
  assign new_n10228 = lo0855 & ~new_n10227 ;
  assign new_n10229 = lo0199 & lo0200 ;
  assign new_n10230 = new_n3113 & ~new_n10229 ;
  assign new_n10231 = ~new_n3116 & ~new_n10230 ;
  assign new_n10232 = ~new_n9165 & new_n10231 ;
  assign new_n10233 = ~new_n9825 & ~new_n10232 ;
  assign new_n10234 = ~lo0199 & lo0200 ;
  assign new_n10235 = lo0198 & new_n10234 ;
  assign new_n10236 = ~lo0199 & ~new_n10235 ;
  assign new_n10237 = new_n10234 & new_n10236 ;
  assign new_n10238 = ~new_n9405 & new_n10237 ;
  assign new_n10239 = ~new_n9305 & new_n10238 ;
  assign new_n10240 = new_n10234 & ~new_n10236 ;
  assign new_n10241 = ~new_n10234 & new_n10236 ;
  assign new_n10242 = ~new_n7385 & new_n10241 ;
  assign new_n10243 = ~new_n10240 & ~new_n10242 ;
  assign new_n10244 = ~new_n10239 & new_n10243 ;
  assign new_n10245 = new_n10236 & ~new_n10244 ;
  assign new_n10246 = ~new_n10236 & new_n10244 ;
  assign new_n10247 = ~new_n10245 & ~new_n10246 ;
  assign new_n10248 = ~new_n8425 & ~new_n10247 ;
  assign new_n10249 = new_n8425 & new_n10245 ;
  assign new_n10250 = ~new_n9305 & new_n9405 ;
  assign new_n10251 = new_n9305 & ~new_n9405 ;
  assign new_n10252 = ~new_n10250 & ~new_n10251 ;
  assign new_n10253 = ~new_n10236 & ~new_n10252 ;
  assign new_n10254 = ~new_n10244 & new_n10253 ;
  assign new_n10255 = ~new_n10249 & ~new_n10254 ;
  assign new_n10256 = ~new_n10248 & new_n10255 ;
  assign new_n10257 = ~lo0198 & new_n10229 ;
  assign new_n10258 = lo0197 & ~new_n10257 ;
  assign new_n10259 = lo0197 & new_n10229 ;
  assign new_n10260 = ~new_n3114 & ~new_n10259 ;
  assign new_n10261 = ~new_n10258 & new_n10260 ;
  assign new_n10262 = ~lo0196 & ~lo0200 ;
  assign new_n10263 = lo0198 & new_n10262 ;
  assign new_n10264 = ~new_n8013 & new_n10262 ;
  assign new_n10265 = lo0199 & new_n10264 ;
  assign new_n10266 = ~lo0196 & ~new_n10265 ;
  assign new_n10267 = ~new_n10264 & ~new_n10266 ;
  assign new_n10268 = ~new_n7293 & new_n10267 ;
  assign new_n10269 = new_n10264 & ~new_n10266 ;
  assign new_n10270 = ~new_n10264 & new_n10266 ;
  assign new_n10271 = ~new_n10269 & ~new_n10270 ;
  assign new_n10272 = ~new_n9405 & ~new_n10271 ;
  assign new_n10273 = new_n9405 & new_n10269 ;
  assign new_n10274 = ~new_n10272 & ~new_n10273 ;
  assign new_n10275 = ~new_n10268 & new_n10274 ;
  assign new_n10276 = ~new_n10263 & ~new_n10275 ;
  assign new_n10277 = new_n10263 & new_n10275 ;
  assign new_n10278 = ~new_n10276 & ~new_n10277 ;
  assign new_n10279 = ~new_n9305 & ~new_n10278 ;
  assign new_n10280 = new_n9305 & new_n10276 ;
  assign new_n10281 = new_n2586 & new_n10263 ;
  assign new_n10282 = ~new_n10275 & new_n10281 ;
  assign new_n10283 = ~new_n10280 & ~new_n10282 ;
  assign new_n10284 = ~new_n10279 & new_n10283 ;
  assign new_n10285 = new_n10261 & ~new_n10284 ;
  assign new_n10286 = new_n10258 & ~new_n10260 ;
  assign new_n10287 = ~new_n10258 & ~new_n10260 ;
  assign new_n10288 = new_n9305 & new_n9405 ;
  assign new_n10289 = new_n10287 & ~new_n10288 ;
  assign new_n10290 = ~new_n10286 & ~new_n10289 ;
  assign new_n10291 = ~new_n10285 & new_n10290 ;
  assign new_n10292 = ~new_n10258 & ~new_n10291 ;
  assign new_n10293 = new_n10258 & new_n10291 ;
  assign new_n10294 = ~new_n10292 & ~new_n10293 ;
  assign new_n10295 = ~new_n10256 & ~new_n10294 ;
  assign new_n10296 = new_n10256 & new_n10292 ;
  assign new_n10297 = new_n9405 & new_n10258 ;
  assign new_n10298 = ~new_n10291 & new_n10297 ;
  assign new_n10299 = ~new_n10296 & ~new_n10298 ;
  assign new_n10300 = ~new_n10295 & new_n10299 ;
  assign new_n10301 = new_n10232 & ~new_n10300 ;
  assign new_n10302 = ~new_n10233 & ~new_n10301 ;
  assign new_n10303 = lo0954 & new_n10302 ;
  assign new_n10304 = new_n10302 & ~new_n10303 ;
  assign new_n10305 = ~new_n9303 & ~new_n10304 ;
  assign new_n10306 = ~lo0954 & new_n9303 ;
  assign new_n10307 = ~new_n10302 & new_n10306 ;
  assign new_n10308 = ~new_n10305 & ~new_n10307 ;
  assign new_n10309 = lo0859 & ~new_n10308 ;
  assign new_n10310 = lo0760 & ~lo0859 ;
  assign new_n10311 = ~new_n10309 & ~new_n10310 ;
  assign new_n10312 = ~lo0858 & ~new_n10311 ;
  assign new_n10313 = lo0858 & new_n2586 ;
  assign new_n10314 = ~lo0857 & ~new_n10313 ;
  assign new_n10315 = ~new_n10312 & new_n10314 ;
  assign new_n10316 = ~lo0855 & ~lo0856 ;
  assign new_n10317 = ~new_n10315 & new_n10316 ;
  assign new_n10318 = ~new_n10228 & ~new_n10317 ;
  assign new_n10319 = ~lo0854 & ~new_n10318 ;
  assign new_n10320 = ~new_n10224 & ~new_n10319 ;
  assign new_n10321 = ~lo0853 & ~new_n10320 ;
  assign new_n10322 = ~new_n2742 & ~new_n10321 ;
  assign new_n10323 = ~lo0848 & ~lo0849 ;
  assign new_n10324 = ~lo0847 & new_n10323 ;
  assign new_n10325 = ~new_n10322 & new_n10324 ;
  assign new_n10326 = new_n3105 & ~new_n3292 ;
  assign new_n10327 = ~new_n9608 & new_n10326 ;
  assign new_n10328 = ~new_n3105 & new_n3292 ;
  assign new_n10329 = new_n9608 & new_n10328 ;
  assign new_n10330 = ~new_n10327 & ~new_n10329 ;
  assign new_n10331 = lo0200 & ~new_n10330 ;
  assign new_n10332 = new_n3105 & new_n3292 ;
  assign new_n10333 = ~new_n9608 & new_n10332 ;
  assign new_n10334 = ~new_n3105 & ~new_n3292 ;
  assign new_n10335 = new_n9608 & new_n10334 ;
  assign new_n10336 = ~new_n10333 & ~new_n10335 ;
  assign new_n10337 = ~lo0200 & ~new_n10336 ;
  assign new_n10338 = ~new_n10331 & ~new_n10337 ;
  assign new_n10339 = lo0199 & ~new_n10338 ;
  assign new_n10340 = new_n3295 & ~new_n9604 ;
  assign new_n10341 = ~new_n3105 & ~new_n10340 ;
  assign new_n10342 = new_n3105 & new_n9600 ;
  assign new_n10343 = ~new_n10341 & ~new_n10342 ;
  assign new_n10344 = ~lo0200 & new_n3111 ;
  assign new_n10345 = ~lo0200 & ~new_n10344 ;
  assign new_n10346 = new_n10343 & ~new_n10345 ;
  assign new_n10347 = new_n3112 & ~new_n10343 ;
  assign new_n10348 = ~new_n10346 & ~new_n10347 ;
  assign new_n10349 = ~lo0199 & ~new_n10348 ;
  assign new_n10350 = ~new_n10339 & ~new_n10349 ;
  assign new_n10351 = lo0848 & ~lo0849 ;
  assign new_n10352 = new_n3116 & new_n10351 ;
  assign new_n10353 = ~new_n9163 & new_n10352 ;
  assign new_n10354 = ~new_n10350 & new_n10353 ;
  assign new_n10355 = ~lo0198 & new_n3100 ;
  assign new_n10356 = new_n3117 & new_n10355 ;
  assign new_n10357 = ~lo0200 & ~new_n9143 ;
  assign new_n10358 = new_n3099 & ~new_n10357 ;
  assign new_n10359 = lo0196 & ~new_n10229 ;
  assign new_n10360 = ~lo0197 & ~new_n10359 ;
  assign new_n10361 = ~new_n10358 & ~new_n10360 ;
  assign new_n10362 = ~new_n10356 & ~new_n10361 ;
  assign new_n10363 = ~new_n10356 & ~new_n10362 ;
  assign new_n10364 = lo0197 & lo0200 ;
  assign new_n10365 = lo0196 & ~lo0198 ;
  assign new_n10366 = ~lo0197 & ~new_n10365 ;
  assign new_n10367 = ~new_n10364 & ~new_n10366 ;
  assign new_n10368 = new_n10362 & ~new_n10367 ;
  assign new_n10369 = ~new_n10363 & ~new_n10368 ;
  assign new_n10370 = ~new_n10362 & ~new_n10369 ;
  assign new_n10371 = ~new_n9608 & new_n10370 ;
  assign new_n10372 = new_n10362 & ~new_n10369 ;
  assign new_n10373 = ~new_n10362 & new_n10369 ;
  assign new_n10374 = ~new_n3292 & new_n10373 ;
  assign new_n10375 = ~new_n10372 & ~new_n10374 ;
  assign new_n10376 = ~new_n10371 & new_n10375 ;
  assign new_n10377 = ~new_n10362 & ~new_n10376 ;
  assign new_n10378 = new_n10362 & new_n10376 ;
  assign new_n10379 = ~new_n10377 & ~new_n10378 ;
  assign new_n10380 = ~new_n7523 & ~new_n10379 ;
  assign new_n10381 = new_n7523 & new_n10377 ;
  assign new_n10382 = ~lo0197 & new_n10262 ;
  assign new_n10383 = lo0197 & ~lo0198 ;
  assign new_n10384 = ~new_n10382 & ~new_n10383 ;
  assign new_n10385 = lo0199 & ~new_n10384 ;
  assign new_n10386 = ~new_n3113 & ~new_n10385 ;
  assign new_n10387 = ~lo0198 & new_n10386 ;
  assign new_n10388 = new_n10382 & ~new_n10387 ;
  assign new_n10389 = new_n10382 & ~new_n10386 ;
  assign new_n10390 = new_n3109 & ~new_n7523 ;
  assign new_n10391 = new_n8013 & ~new_n8551 ;
  assign new_n10392 = ~new_n10390 & ~new_n10391 ;
  assign new_n10393 = lo0197 & ~lo0199 ;
  assign new_n10394 = lo0197 & ~new_n9267 ;
  assign new_n10395 = ~new_n10332 & ~new_n10334 ;
  assign new_n10396 = ~new_n10393 & ~new_n10395 ;
  assign new_n10397 = ~new_n10326 & ~new_n10328 ;
  assign new_n10398 = ~new_n10396 & new_n10397 ;
  assign new_n10399 = new_n10394 & ~new_n10398 ;
  assign new_n10400 = new_n10393 & ~new_n10394 ;
  assign new_n10401 = new_n10334 & new_n10400 ;
  assign new_n10402 = ~new_n10399 & ~new_n10401 ;
  assign new_n10403 = new_n10393 & ~new_n10402 ;
  assign new_n10404 = ~new_n10393 & new_n10402 ;
  assign new_n10405 = ~new_n10403 & ~new_n10404 ;
  assign new_n10406 = ~new_n10392 & ~new_n10405 ;
  assign new_n10407 = new_n10392 & new_n10403 ;
  assign new_n10408 = new_n3292 & ~new_n10393 ;
  assign new_n10409 = ~new_n10402 & new_n10408 ;
  assign new_n10410 = ~new_n10407 & ~new_n10409 ;
  assign new_n10411 = ~new_n10406 & new_n10410 ;
  assign new_n10412 = new_n10389 & new_n10411 ;
  assign new_n10413 = ~new_n10382 & new_n10386 ;
  assign new_n10414 = ~new_n10389 & ~new_n10413 ;
  assign new_n10415 = ~new_n10411 & ~new_n10414 ;
  assign new_n10416 = ~new_n10382 & ~new_n10386 ;
  assign new_n10417 = ~new_n10332 & new_n10416 ;
  assign new_n10418 = ~new_n10415 & ~new_n10417 ;
  assign new_n10419 = ~new_n10412 & new_n10418 ;
  assign new_n10420 = ~new_n10388 & ~new_n10419 ;
  assign new_n10421 = new_n10388 & new_n10419 ;
  assign new_n10422 = ~new_n10420 & ~new_n10421 ;
  assign new_n10423 = ~new_n3105 & ~new_n10422 ;
  assign new_n10424 = new_n3105 & new_n10420 ;
  assign new_n10425 = new_n2718 & new_n10388 ;
  assign new_n10426 = ~new_n10419 & new_n10425 ;
  assign new_n10427 = ~new_n10424 & ~new_n10426 ;
  assign new_n10428 = ~new_n10423 & new_n10427 ;
  assign new_n10429 = new_n10362 & ~new_n10428 ;
  assign new_n10430 = ~new_n10376 & new_n10429 ;
  assign new_n10431 = ~new_n10381 & ~new_n10430 ;
  assign new_n10432 = ~new_n10380 & new_n10431 ;
  assign new_n10433 = ~new_n3650 & new_n10373 ;
  assign new_n10434 = new_n10362 & new_n10369 ;
  assign new_n10435 = ~new_n7648 & new_n10434 ;
  assign new_n10436 = ~new_n10372 & ~new_n10435 ;
  assign new_n10437 = ~new_n10433 & new_n10436 ;
  assign new_n10438 = new_n10369 & ~new_n10437 ;
  assign new_n10439 = new_n9615 & new_n10438 ;
  assign new_n10440 = ~new_n10369 & new_n10437 ;
  assign new_n10441 = ~new_n10438 & ~new_n10440 ;
  assign new_n10442 = ~new_n9615 & ~new_n10441 ;
  assign new_n10443 = new_n3557 & ~new_n3650 ;
  assign new_n10444 = ~new_n3557 & new_n3650 ;
  assign new_n10445 = ~new_n10443 & ~new_n10444 ;
  assign new_n10446 = ~new_n10393 & ~new_n10394 ;
  assign new_n10447 = ~new_n10392 & new_n10446 ;
  assign new_n10448 = ~new_n10393 & new_n10394 ;
  assign new_n10449 = ~new_n3557 & new_n10400 ;
  assign new_n10450 = ~new_n3650 & new_n10449 ;
  assign new_n10451 = ~new_n10448 & ~new_n10450 ;
  assign new_n10452 = ~new_n10447 & new_n10451 ;
  assign new_n10453 = new_n10394 & new_n10452 ;
  assign new_n10454 = ~new_n10394 & ~new_n10452 ;
  assign new_n10455 = ~new_n10453 & ~new_n10454 ;
  assign new_n10456 = ~new_n10445 & ~new_n10455 ;
  assign new_n10457 = new_n3650 & new_n10394 ;
  assign new_n10458 = ~new_n3650 & ~new_n10394 ;
  assign new_n10459 = ~new_n10457 & ~new_n10458 ;
  assign new_n10460 = ~new_n3557 & ~new_n10459 ;
  assign new_n10461 = new_n3557 & new_n3650 ;
  assign new_n10462 = ~new_n10460 & ~new_n10461 ;
  assign new_n10463 = ~new_n10452 & ~new_n10462 ;
  assign new_n10464 = ~new_n10456 & ~new_n10463 ;
  assign new_n10465 = new_n10389 & new_n10464 ;
  assign new_n10466 = ~new_n10414 & ~new_n10464 ;
  assign new_n10467 = new_n10416 & ~new_n10461 ;
  assign new_n10468 = ~new_n10466 & ~new_n10467 ;
  assign new_n10469 = ~new_n10465 & new_n10468 ;
  assign new_n10470 = ~new_n10388 & ~new_n10469 ;
  assign new_n10471 = new_n10388 & new_n10469 ;
  assign new_n10472 = ~new_n10470 & ~new_n10471 ;
  assign new_n10473 = ~new_n3557 & ~new_n10472 ;
  assign new_n10474 = new_n3557 & new_n10470 ;
  assign new_n10475 = new_n3081 & new_n10388 ;
  assign new_n10476 = ~new_n10469 & new_n10475 ;
  assign new_n10477 = ~new_n10474 & ~new_n10476 ;
  assign new_n10478 = ~new_n10473 & new_n10477 ;
  assign new_n10479 = ~new_n10369 & ~new_n10437 ;
  assign new_n10480 = ~new_n10478 & new_n10479 ;
  assign new_n10481 = ~new_n10442 & ~new_n10480 ;
  assign new_n10482 = ~new_n10439 & new_n10481 ;
  assign new_n10483 = ~new_n9622 & new_n10370 ;
  assign new_n10484 = ~new_n4014 & new_n10373 ;
  assign new_n10485 = ~new_n10372 & ~new_n10484 ;
  assign new_n10486 = ~new_n10483 & new_n10485 ;
  assign new_n10487 = ~new_n10362 & ~new_n10486 ;
  assign new_n10488 = new_n10362 & new_n10486 ;
  assign new_n10489 = ~new_n10487 & ~new_n10488 ;
  assign new_n10490 = ~new_n7772 & ~new_n10489 ;
  assign new_n10491 = new_n7772 & new_n10487 ;
  assign new_n10492 = ~new_n3922 & ~new_n4014 ;
  assign new_n10493 = new_n3922 & new_n4014 ;
  assign new_n10494 = ~new_n10492 & ~new_n10493 ;
  assign new_n10495 = ~new_n10393 & ~new_n10494 ;
  assign new_n10496 = ~new_n3922 & new_n4014 ;
  assign new_n10497 = new_n3922 & ~new_n4014 ;
  assign new_n10498 = ~new_n10496 & ~new_n10497 ;
  assign new_n10499 = ~new_n10495 & new_n10498 ;
  assign new_n10500 = new_n10394 & ~new_n10499 ;
  assign new_n10501 = new_n10400 & new_n10492 ;
  assign new_n10502 = ~new_n10500 & ~new_n10501 ;
  assign new_n10503 = new_n10393 & ~new_n10502 ;
  assign new_n10504 = ~new_n10393 & new_n10502 ;
  assign new_n10505 = ~new_n10503 & ~new_n10504 ;
  assign new_n10506 = ~new_n10392 & ~new_n10505 ;
  assign new_n10507 = new_n10392 & new_n10503 ;
  assign new_n10508 = new_n4014 & ~new_n10393 ;
  assign new_n10509 = ~new_n10502 & new_n10508 ;
  assign new_n10510 = ~new_n10507 & ~new_n10509 ;
  assign new_n10511 = ~new_n10506 & new_n10510 ;
  assign new_n10512 = new_n10389 & new_n10511 ;
  assign new_n10513 = ~new_n10414 & ~new_n10511 ;
  assign new_n10514 = new_n10416 & ~new_n10493 ;
  assign new_n10515 = ~new_n10513 & ~new_n10514 ;
  assign new_n10516 = ~new_n10512 & new_n10515 ;
  assign new_n10517 = ~new_n10388 & ~new_n10516 ;
  assign new_n10518 = new_n10388 & new_n10516 ;
  assign new_n10519 = ~new_n10517 & ~new_n10518 ;
  assign new_n10520 = ~new_n3922 & ~new_n10519 ;
  assign new_n10521 = new_n3922 & new_n10517 ;
  assign new_n10522 = new_n2990 & new_n10388 ;
  assign new_n10523 = ~new_n10516 & new_n10522 ;
  assign new_n10524 = ~new_n10521 & ~new_n10523 ;
  assign new_n10525 = ~new_n10520 & new_n10524 ;
  assign new_n10526 = new_n10362 & ~new_n10525 ;
  assign new_n10527 = ~new_n10486 & new_n10526 ;
  assign new_n10528 = ~new_n10491 & ~new_n10527 ;
  assign new_n10529 = ~new_n10490 & new_n10528 ;
  assign new_n10530 = ~new_n4373 & new_n10373 ;
  assign new_n10531 = ~new_n7894 & new_n10434 ;
  assign new_n10532 = ~new_n10372 & ~new_n10531 ;
  assign new_n10533 = ~new_n10530 & new_n10532 ;
  assign new_n10534 = new_n10369 & ~new_n10533 ;
  assign new_n10535 = new_n9629 & new_n10534 ;
  assign new_n10536 = ~new_n10369 & new_n10533 ;
  assign new_n10537 = ~new_n10534 & ~new_n10536 ;
  assign new_n10538 = ~new_n9629 & ~new_n10537 ;
  assign new_n10539 = new_n4281 & ~new_n4373 ;
  assign new_n10540 = ~new_n4281 & new_n4373 ;
  assign new_n10541 = ~new_n10539 & ~new_n10540 ;
  assign new_n10542 = ~new_n10447 & ~new_n10448 ;
  assign new_n10543 = ~new_n4373 & new_n10400 ;
  assign new_n10544 = ~new_n4281 & new_n10543 ;
  assign new_n10545 = new_n10542 & ~new_n10544 ;
  assign new_n10546 = new_n10394 & new_n10545 ;
  assign new_n10547 = ~new_n10394 & ~new_n10545 ;
  assign new_n10548 = ~new_n10546 & ~new_n10547 ;
  assign new_n10549 = ~new_n10541 & ~new_n10548 ;
  assign new_n10550 = new_n4373 & new_n10394 ;
  assign new_n10551 = ~new_n4373 & ~new_n10394 ;
  assign new_n10552 = ~new_n10550 & ~new_n10551 ;
  assign new_n10553 = ~new_n4281 & ~new_n10552 ;
  assign new_n10554 = new_n4281 & new_n4373 ;
  assign new_n10555 = ~new_n10553 & ~new_n10554 ;
  assign new_n10556 = ~new_n10545 & ~new_n10555 ;
  assign new_n10557 = ~new_n10549 & ~new_n10556 ;
  assign new_n10558 = new_n10389 & new_n10557 ;
  assign new_n10559 = ~new_n10414 & ~new_n10557 ;
  assign new_n10560 = new_n10416 & ~new_n10554 ;
  assign new_n10561 = ~new_n10559 & ~new_n10560 ;
  assign new_n10562 = ~new_n10558 & new_n10561 ;
  assign new_n10563 = ~new_n10388 & ~new_n10562 ;
  assign new_n10564 = new_n10388 & new_n10562 ;
  assign new_n10565 = ~new_n10563 & ~new_n10564 ;
  assign new_n10566 = ~new_n4281 & ~new_n10565 ;
  assign new_n10567 = new_n4281 & new_n10563 ;
  assign new_n10568 = new_n3453 & new_n10388 ;
  assign new_n10569 = ~new_n10562 & new_n10568 ;
  assign new_n10570 = ~new_n10567 & ~new_n10569 ;
  assign new_n10571 = ~new_n10566 & new_n10570 ;
  assign new_n10572 = ~new_n10369 & ~new_n10533 ;
  assign new_n10573 = ~new_n10571 & new_n10572 ;
  assign new_n10574 = ~new_n10538 & ~new_n10573 ;
  assign new_n10575 = ~new_n10535 & new_n10574 ;
  assign new_n10576 = ~new_n9636 & new_n10370 ;
  assign new_n10577 = ~new_n4735 & new_n10373 ;
  assign new_n10578 = ~new_n10372 & ~new_n10577 ;
  assign new_n10579 = ~new_n10576 & new_n10578 ;
  assign new_n10580 = ~new_n10362 & ~new_n10579 ;
  assign new_n10581 = new_n10362 & new_n10579 ;
  assign new_n10582 = ~new_n10580 & ~new_n10581 ;
  assign new_n10583 = ~new_n8035 & ~new_n10582 ;
  assign new_n10584 = new_n8035 & new_n10580 ;
  assign new_n10585 = ~new_n4643 & ~new_n4735 ;
  assign new_n10586 = new_n4643 & new_n4735 ;
  assign new_n10587 = ~new_n10585 & ~new_n10586 ;
  assign new_n10588 = ~new_n10393 & ~new_n10587 ;
  assign new_n10589 = ~new_n4643 & new_n4735 ;
  assign new_n10590 = new_n4643 & ~new_n4735 ;
  assign new_n10591 = ~new_n10589 & ~new_n10590 ;
  assign new_n10592 = ~new_n10588 & new_n10591 ;
  assign new_n10593 = new_n10394 & ~new_n10592 ;
  assign new_n10594 = new_n10400 & new_n10585 ;
  assign new_n10595 = ~new_n10593 & ~new_n10594 ;
  assign new_n10596 = new_n10393 & ~new_n10595 ;
  assign new_n10597 = ~new_n10393 & new_n10595 ;
  assign new_n10598 = ~new_n10596 & ~new_n10597 ;
  assign new_n10599 = ~new_n10392 & ~new_n10598 ;
  assign new_n10600 = new_n10392 & new_n10596 ;
  assign new_n10601 = new_n4735 & ~new_n10393 ;
  assign new_n10602 = ~new_n10595 & new_n10601 ;
  assign new_n10603 = ~new_n10600 & ~new_n10602 ;
  assign new_n10604 = ~new_n10599 & new_n10603 ;
  assign new_n10605 = new_n10389 & new_n10604 ;
  assign new_n10606 = ~new_n10414 & ~new_n10604 ;
  assign new_n10607 = new_n10416 & ~new_n10586 ;
  assign new_n10608 = ~new_n10606 & ~new_n10607 ;
  assign new_n10609 = ~new_n10605 & new_n10608 ;
  assign new_n10610 = ~new_n10388 & ~new_n10609 ;
  assign new_n10611 = new_n10388 & new_n10609 ;
  assign new_n10612 = ~new_n10610 & ~new_n10611 ;
  assign new_n10613 = ~new_n4643 & ~new_n10612 ;
  assign new_n10614 = new_n4643 & new_n10610 ;
  assign new_n10615 = new_n3806 & new_n10388 ;
  assign new_n10616 = ~new_n10609 & new_n10615 ;
  assign new_n10617 = ~new_n10614 & ~new_n10616 ;
  assign new_n10618 = ~new_n10613 & new_n10617 ;
  assign new_n10619 = new_n10362 & ~new_n10618 ;
  assign new_n10620 = ~new_n10579 & new_n10619 ;
  assign new_n10621 = ~new_n10584 & ~new_n10620 ;
  assign new_n10622 = ~new_n10583 & new_n10621 ;
  assign new_n10623 = ~new_n5097 & new_n10373 ;
  assign new_n10624 = ~new_n8163 & new_n10434 ;
  assign new_n10625 = ~new_n10372 & ~new_n10624 ;
  assign new_n10626 = ~new_n10623 & new_n10625 ;
  assign new_n10627 = new_n10369 & ~new_n10626 ;
  assign new_n10628 = new_n9643 & new_n10627 ;
  assign new_n10629 = ~new_n10369 & new_n10626 ;
  assign new_n10630 = ~new_n10627 & ~new_n10629 ;
  assign new_n10631 = ~new_n9643 & ~new_n10630 ;
  assign new_n10632 = new_n5005 & ~new_n5097 ;
  assign new_n10633 = ~new_n5005 & new_n5097 ;
  assign new_n10634 = ~new_n10632 & ~new_n10633 ;
  assign new_n10635 = ~new_n5097 & new_n10400 ;
  assign new_n10636 = ~new_n5005 & new_n10635 ;
  assign new_n10637 = new_n10542 & ~new_n10636 ;
  assign new_n10638 = new_n10394 & new_n10637 ;
  assign new_n10639 = ~new_n10394 & ~new_n10637 ;
  assign new_n10640 = ~new_n10638 & ~new_n10639 ;
  assign new_n10641 = ~new_n10634 & ~new_n10640 ;
  assign new_n10642 = new_n5097 & new_n10394 ;
  assign new_n10643 = ~new_n5097 & ~new_n10394 ;
  assign new_n10644 = ~new_n10642 & ~new_n10643 ;
  assign new_n10645 = ~new_n5005 & ~new_n10644 ;
  assign new_n10646 = new_n5005 & new_n5097 ;
  assign new_n10647 = ~new_n10645 & ~new_n10646 ;
  assign new_n10648 = ~new_n10637 & ~new_n10647 ;
  assign new_n10649 = ~new_n10641 & ~new_n10648 ;
  assign new_n10650 = new_n10389 & new_n10649 ;
  assign new_n10651 = ~new_n10414 & ~new_n10649 ;
  assign new_n10652 = new_n10416 & ~new_n10646 ;
  assign new_n10653 = ~new_n10651 & ~new_n10652 ;
  assign new_n10654 = ~new_n10650 & new_n10653 ;
  assign new_n10655 = ~new_n10388 & ~new_n10654 ;
  assign new_n10656 = new_n10388 & new_n10654 ;
  assign new_n10657 = ~new_n10655 & ~new_n10656 ;
  assign new_n10658 = ~new_n5005 & ~new_n10657 ;
  assign new_n10659 = new_n5005 & new_n10655 ;
  assign new_n10660 = new_n4086 & new_n10388 ;
  assign new_n10661 = ~new_n10654 & new_n10660 ;
  assign new_n10662 = ~new_n10659 & ~new_n10661 ;
  assign new_n10663 = ~new_n10658 & new_n10662 ;
  assign new_n10664 = ~new_n10369 & ~new_n10626 ;
  assign new_n10665 = ~new_n10663 & new_n10664 ;
  assign new_n10666 = ~new_n10631 & ~new_n10665 ;
  assign new_n10667 = ~new_n10628 & new_n10666 ;
  assign new_n10668 = ~new_n9650 & new_n10370 ;
  assign new_n10669 = ~new_n5381 & new_n10373 ;
  assign new_n10670 = ~new_n10372 & ~new_n10669 ;
  assign new_n10671 = ~new_n10668 & new_n10670 ;
  assign new_n10672 = ~new_n10362 & ~new_n10671 ;
  assign new_n10673 = new_n10362 & new_n10671 ;
  assign new_n10674 = ~new_n10672 & ~new_n10673 ;
  assign new_n10675 = ~new_n8295 & ~new_n10674 ;
  assign new_n10676 = new_n8295 & new_n10672 ;
  assign new_n10677 = ~new_n5289 & ~new_n5381 ;
  assign new_n10678 = new_n5289 & new_n5381 ;
  assign new_n10679 = ~new_n10677 & ~new_n10678 ;
  assign new_n10680 = ~new_n10393 & ~new_n10679 ;
  assign new_n10681 = ~new_n5289 & new_n5381 ;
  assign new_n10682 = new_n5289 & ~new_n5381 ;
  assign new_n10683 = ~new_n10681 & ~new_n10682 ;
  assign new_n10684 = ~new_n10680 & new_n10683 ;
  assign new_n10685 = new_n10394 & ~new_n10684 ;
  assign new_n10686 = new_n10400 & new_n10677 ;
  assign new_n10687 = ~new_n10685 & ~new_n10686 ;
  assign new_n10688 = new_n10393 & ~new_n10687 ;
  assign new_n10689 = ~new_n10393 & new_n10687 ;
  assign new_n10690 = ~new_n10688 & ~new_n10689 ;
  assign new_n10691 = ~new_n10392 & ~new_n10690 ;
  assign new_n10692 = new_n10392 & new_n10688 ;
  assign new_n10693 = new_n5381 & ~new_n10393 ;
  assign new_n10694 = ~new_n10687 & new_n10693 ;
  assign new_n10695 = ~new_n10692 & ~new_n10694 ;
  assign new_n10696 = ~new_n10691 & new_n10695 ;
  assign new_n10697 = new_n10389 & new_n10696 ;
  assign new_n10698 = ~new_n10414 & ~new_n10696 ;
  assign new_n10699 = new_n10416 & ~new_n10678 ;
  assign new_n10700 = ~new_n10698 & ~new_n10699 ;
  assign new_n10701 = ~new_n10697 & new_n10700 ;
  assign new_n10702 = ~new_n10388 & ~new_n10701 ;
  assign new_n10703 = new_n10388 & new_n10701 ;
  assign new_n10704 = ~new_n10702 & ~new_n10703 ;
  assign new_n10705 = ~new_n5289 & ~new_n10704 ;
  assign new_n10706 = new_n5289 & new_n10702 ;
  assign new_n10707 = new_n4530 & new_n10388 ;
  assign new_n10708 = ~new_n10701 & new_n10707 ;
  assign new_n10709 = ~new_n10706 & ~new_n10708 ;
  assign new_n10710 = ~new_n10705 & new_n10709 ;
  assign new_n10711 = new_n10362 & ~new_n10710 ;
  assign new_n10712 = ~new_n10671 & new_n10711 ;
  assign new_n10713 = ~new_n10676 & ~new_n10712 ;
  assign new_n10714 = ~new_n10675 & new_n10713 ;
  assign new_n10715 = ~new_n5665 & new_n10373 ;
  assign new_n10716 = ~new_n8425 & new_n10434 ;
  assign new_n10717 = ~new_n10372 & ~new_n10716 ;
  assign new_n10718 = ~new_n10715 & new_n10717 ;
  assign new_n10719 = new_n10369 & ~new_n10718 ;
  assign new_n10720 = new_n9657 & new_n10719 ;
  assign new_n10721 = ~new_n10369 & new_n10718 ;
  assign new_n10722 = ~new_n10719 & ~new_n10721 ;
  assign new_n10723 = ~new_n9657 & ~new_n10722 ;
  assign new_n10724 = new_n5573 & ~new_n5665 ;
  assign new_n10725 = ~new_n5573 & new_n5665 ;
  assign new_n10726 = ~new_n10724 & ~new_n10725 ;
  assign new_n10727 = ~new_n5665 & new_n10400 ;
  assign new_n10728 = ~new_n5573 & new_n10727 ;
  assign new_n10729 = new_n10542 & ~new_n10728 ;
  assign new_n10730 = new_n10394 & new_n10729 ;
  assign new_n10731 = ~new_n10394 & ~new_n10729 ;
  assign new_n10732 = ~new_n10730 & ~new_n10731 ;
  assign new_n10733 = ~new_n10726 & ~new_n10732 ;
  assign new_n10734 = new_n5665 & new_n10394 ;
  assign new_n10735 = ~new_n5665 & ~new_n10394 ;
  assign new_n10736 = ~new_n10734 & ~new_n10735 ;
  assign new_n10737 = ~new_n5573 & ~new_n10736 ;
  assign new_n10738 = new_n5573 & new_n5665 ;
  assign new_n10739 = ~new_n10737 & ~new_n10738 ;
  assign new_n10740 = ~new_n10729 & ~new_n10739 ;
  assign new_n10741 = ~new_n10733 & ~new_n10740 ;
  assign new_n10742 = new_n10389 & new_n10741 ;
  assign new_n10743 = ~new_n10414 & ~new_n10741 ;
  assign new_n10744 = new_n10416 & ~new_n10738 ;
  assign new_n10745 = ~new_n10743 & ~new_n10744 ;
  assign new_n10746 = ~new_n10742 & new_n10745 ;
  assign new_n10747 = ~new_n10388 & ~new_n10746 ;
  assign new_n10748 = new_n10388 & new_n10746 ;
  assign new_n10749 = ~new_n10747 & ~new_n10748 ;
  assign new_n10750 = ~new_n5573 & ~new_n10749 ;
  assign new_n10751 = new_n5573 & new_n10747 ;
  assign new_n10752 = new_n4807 & new_n10388 ;
  assign new_n10753 = ~new_n10746 & new_n10752 ;
  assign new_n10754 = ~new_n10751 & ~new_n10753 ;
  assign new_n10755 = ~new_n10750 & new_n10754 ;
  assign new_n10756 = ~new_n10369 & ~new_n10718 ;
  assign new_n10757 = ~new_n10755 & new_n10756 ;
  assign new_n10758 = ~new_n10723 & ~new_n10757 ;
  assign new_n10759 = ~new_n10720 & new_n10758 ;
  assign new_n10760 = ~new_n9664 & new_n10370 ;
  assign new_n10761 = ~new_n5891 & new_n10373 ;
  assign new_n10762 = ~new_n10372 & ~new_n10761 ;
  assign new_n10763 = ~new_n10760 & new_n10762 ;
  assign new_n10764 = ~new_n10362 & ~new_n10763 ;
  assign new_n10765 = new_n10362 & new_n10763 ;
  assign new_n10766 = ~new_n10764 & ~new_n10765 ;
  assign new_n10767 = ~new_n8551 & ~new_n10766 ;
  assign new_n10768 = new_n8551 & new_n10764 ;
  assign new_n10769 = ~new_n5799 & ~new_n5891 ;
  assign new_n10770 = new_n5799 & new_n5891 ;
  assign new_n10771 = ~new_n10769 & ~new_n10770 ;
  assign new_n10772 = ~new_n10393 & ~new_n10771 ;
  assign new_n10773 = new_n5799 & ~new_n5891 ;
  assign new_n10774 = ~new_n5799 & new_n5891 ;
  assign new_n10775 = ~new_n10773 & ~new_n10774 ;
  assign new_n10776 = ~new_n10772 & new_n10775 ;
  assign new_n10777 = new_n10394 & ~new_n10776 ;
  assign new_n10778 = new_n10400 & new_n10769 ;
  assign new_n10779 = ~new_n10777 & ~new_n10778 ;
  assign new_n10780 = new_n10393 & ~new_n10779 ;
  assign new_n10781 = ~new_n10393 & new_n10779 ;
  assign new_n10782 = ~new_n10780 & ~new_n10781 ;
  assign new_n10783 = ~new_n10392 & ~new_n10782 ;
  assign new_n10784 = new_n10392 & new_n10780 ;
  assign new_n10785 = new_n5891 & ~new_n10393 ;
  assign new_n10786 = ~new_n10779 & new_n10785 ;
  assign new_n10787 = ~new_n10784 & ~new_n10786 ;
  assign new_n10788 = ~new_n10783 & new_n10787 ;
  assign new_n10789 = new_n10389 & new_n10788 ;
  assign new_n10790 = ~new_n10414 & ~new_n10788 ;
  assign new_n10791 = new_n10416 & ~new_n10770 ;
  assign new_n10792 = ~new_n10790 & ~new_n10791 ;
  assign new_n10793 = ~new_n10789 & new_n10792 ;
  assign new_n10794 = ~new_n10388 & ~new_n10793 ;
  assign new_n10795 = new_n10388 & new_n10793 ;
  assign new_n10796 = ~new_n10794 & ~new_n10795 ;
  assign new_n10797 = ~new_n5799 & ~new_n10796 ;
  assign new_n10798 = new_n5799 & new_n10794 ;
  assign new_n10799 = new_n2813 & new_n10388 ;
  assign new_n10800 = ~new_n10793 & new_n10799 ;
  assign new_n10801 = ~new_n10798 & ~new_n10800 ;
  assign new_n10802 = ~new_n10797 & new_n10801 ;
  assign new_n10803 = new_n10362 & ~new_n10802 ;
  assign new_n10804 = ~new_n10763 & new_n10803 ;
  assign new_n10805 = ~new_n10768 & ~new_n10804 ;
  assign new_n10806 = ~new_n10767 & new_n10805 ;
  assign new_n10807 = ~new_n6117 & new_n10373 ;
  assign new_n10808 = ~new_n8672 & new_n10434 ;
  assign new_n10809 = ~new_n10372 & ~new_n10808 ;
  assign new_n10810 = ~new_n10807 & new_n10809 ;
  assign new_n10811 = new_n10369 & ~new_n10810 ;
  assign new_n10812 = new_n9671 & new_n10811 ;
  assign new_n10813 = ~new_n10369 & new_n10810 ;
  assign new_n10814 = ~new_n10811 & ~new_n10813 ;
  assign new_n10815 = ~new_n9671 & ~new_n10814 ;
  assign new_n10816 = new_n6025 & ~new_n6117 ;
  assign new_n10817 = ~new_n6025 & new_n6117 ;
  assign new_n10818 = ~new_n10816 & ~new_n10817 ;
  assign new_n10819 = ~new_n6117 & new_n10400 ;
  assign new_n10820 = ~new_n6025 & new_n10819 ;
  assign new_n10821 = new_n10542 & ~new_n10820 ;
  assign new_n10822 = new_n10394 & new_n10821 ;
  assign new_n10823 = ~new_n10394 & ~new_n10821 ;
  assign new_n10824 = ~new_n10822 & ~new_n10823 ;
  assign new_n10825 = ~new_n10818 & ~new_n10824 ;
  assign new_n10826 = new_n6117 & new_n10394 ;
  assign new_n10827 = ~new_n6117 & ~new_n10394 ;
  assign new_n10828 = ~new_n10826 & ~new_n10827 ;
  assign new_n10829 = ~new_n6025 & ~new_n10828 ;
  assign new_n10830 = new_n6025 & new_n6117 ;
  assign new_n10831 = ~new_n10829 & ~new_n10830 ;
  assign new_n10832 = ~new_n10821 & ~new_n10831 ;
  assign new_n10833 = ~new_n10825 & ~new_n10832 ;
  assign new_n10834 = new_n10389 & new_n10833 ;
  assign new_n10835 = ~new_n10414 & ~new_n10833 ;
  assign new_n10836 = new_n10416 & ~new_n10830 ;
  assign new_n10837 = ~new_n10835 & ~new_n10836 ;
  assign new_n10838 = ~new_n10834 & new_n10837 ;
  assign new_n10839 = ~new_n10388 & ~new_n10838 ;
  assign new_n10840 = new_n10388 & new_n10838 ;
  assign new_n10841 = ~new_n10839 & ~new_n10840 ;
  assign new_n10842 = ~new_n6025 & ~new_n10841 ;
  assign new_n10843 = new_n6025 & new_n10839 ;
  assign new_n10844 = new_n3538 & new_n10388 ;
  assign new_n10845 = ~new_n10838 & new_n10844 ;
  assign new_n10846 = ~new_n10843 & ~new_n10845 ;
  assign new_n10847 = ~new_n10842 & new_n10846 ;
  assign new_n10848 = ~new_n10369 & ~new_n10810 ;
  assign new_n10849 = ~new_n10847 & new_n10848 ;
  assign new_n10850 = ~new_n10815 & ~new_n10849 ;
  assign new_n10851 = ~new_n10812 & new_n10850 ;
  assign new_n10852 = ~new_n9678 & new_n10370 ;
  assign new_n10853 = ~new_n6347 & new_n10373 ;
  assign new_n10854 = ~new_n10372 & ~new_n10853 ;
  assign new_n10855 = ~new_n10852 & new_n10854 ;
  assign new_n10856 = ~new_n10362 & ~new_n10855 ;
  assign new_n10857 = new_n10362 & new_n10855 ;
  assign new_n10858 = ~new_n10856 & ~new_n10857 ;
  assign new_n10859 = ~new_n8794 & ~new_n10858 ;
  assign new_n10860 = new_n8794 & new_n10856 ;
  assign new_n10861 = ~new_n6255 & ~new_n6347 ;
  assign new_n10862 = new_n6255 & new_n6347 ;
  assign new_n10863 = ~new_n10861 & ~new_n10862 ;
  assign new_n10864 = ~new_n10393 & ~new_n10863 ;
  assign new_n10865 = new_n6255 & ~new_n6347 ;
  assign new_n10866 = ~new_n6255 & new_n6347 ;
  assign new_n10867 = ~new_n10865 & ~new_n10866 ;
  assign new_n10868 = ~new_n10864 & new_n10867 ;
  assign new_n10869 = new_n10394 & ~new_n10868 ;
  assign new_n10870 = new_n10400 & new_n10861 ;
  assign new_n10871 = ~new_n10869 & ~new_n10870 ;
  assign new_n10872 = new_n10393 & ~new_n10871 ;
  assign new_n10873 = ~new_n10393 & new_n10871 ;
  assign new_n10874 = ~new_n10872 & ~new_n10873 ;
  assign new_n10875 = ~new_n10392 & ~new_n10874 ;
  assign new_n10876 = new_n10392 & new_n10872 ;
  assign new_n10877 = new_n6347 & ~new_n10393 ;
  assign new_n10878 = ~new_n10871 & new_n10877 ;
  assign new_n10879 = ~new_n10876 & ~new_n10878 ;
  assign new_n10880 = ~new_n10875 & new_n10879 ;
  assign new_n10881 = new_n10389 & new_n10880 ;
  assign new_n10882 = ~new_n10414 & ~new_n10880 ;
  assign new_n10883 = new_n10416 & ~new_n10862 ;
  assign new_n10884 = ~new_n10882 & ~new_n10883 ;
  assign new_n10885 = ~new_n10881 & new_n10884 ;
  assign new_n10886 = ~new_n10388 & ~new_n10885 ;
  assign new_n10887 = new_n10388 & new_n10885 ;
  assign new_n10888 = ~new_n10886 & ~new_n10887 ;
  assign new_n10889 = ~new_n6255 & ~new_n10888 ;
  assign new_n10890 = new_n6255 & new_n10886 ;
  assign new_n10891 = new_n3897 & new_n10388 ;
  assign new_n10892 = ~new_n10885 & new_n10891 ;
  assign new_n10893 = ~new_n10890 & ~new_n10892 ;
  assign new_n10894 = ~new_n10889 & new_n10893 ;
  assign new_n10895 = new_n10362 & ~new_n10894 ;
  assign new_n10896 = ~new_n10855 & new_n10895 ;
  assign new_n10897 = ~new_n10860 & ~new_n10896 ;
  assign new_n10898 = ~new_n10859 & new_n10897 ;
  assign new_n10899 = ~new_n6582 & new_n10373 ;
  assign new_n10900 = ~new_n8915 & new_n10434 ;
  assign new_n10901 = ~new_n10372 & ~new_n10900 ;
  assign new_n10902 = ~new_n10899 & new_n10901 ;
  assign new_n10903 = new_n10369 & ~new_n10902 ;
  assign new_n10904 = new_n9685 & new_n10903 ;
  assign new_n10905 = ~new_n10369 & new_n10902 ;
  assign new_n10906 = ~new_n10903 & ~new_n10905 ;
  assign new_n10907 = ~new_n9685 & ~new_n10906 ;
  assign new_n10908 = new_n6490 & ~new_n6582 ;
  assign new_n10909 = ~new_n6490 & new_n6582 ;
  assign new_n10910 = ~new_n10908 & ~new_n10909 ;
  assign new_n10911 = ~new_n6582 & new_n10400 ;
  assign new_n10912 = ~new_n6490 & new_n10911 ;
  assign new_n10913 = new_n10542 & ~new_n10912 ;
  assign new_n10914 = new_n10394 & new_n10913 ;
  assign new_n10915 = ~new_n10394 & ~new_n10913 ;
  assign new_n10916 = ~new_n10914 & ~new_n10915 ;
  assign new_n10917 = ~new_n10910 & ~new_n10916 ;
  assign new_n10918 = new_n6582 & new_n10394 ;
  assign new_n10919 = ~new_n6582 & ~new_n10394 ;
  assign new_n10920 = ~new_n10918 & ~new_n10919 ;
  assign new_n10921 = ~new_n6490 & ~new_n10920 ;
  assign new_n10922 = new_n6490 & new_n6582 ;
  assign new_n10923 = ~new_n10921 & ~new_n10922 ;
  assign new_n10924 = ~new_n10913 & ~new_n10923 ;
  assign new_n10925 = ~new_n10917 & ~new_n10924 ;
  assign new_n10926 = new_n10389 & new_n10925 ;
  assign new_n10927 = ~new_n10414 & ~new_n10925 ;
  assign new_n10928 = new_n10416 & ~new_n10922 ;
  assign new_n10929 = ~new_n10927 & ~new_n10928 ;
  assign new_n10930 = ~new_n10926 & new_n10929 ;
  assign new_n10931 = ~new_n10388 & ~new_n10930 ;
  assign new_n10932 = new_n10388 & new_n10930 ;
  assign new_n10933 = ~new_n10931 & ~new_n10932 ;
  assign new_n10934 = ~new_n6490 & ~new_n10933 ;
  assign new_n10935 = new_n6490 & new_n10931 ;
  assign new_n10936 = new_n4257 & new_n10388 ;
  assign new_n10937 = ~new_n10930 & new_n10936 ;
  assign new_n10938 = ~new_n10935 & ~new_n10937 ;
  assign new_n10939 = ~new_n10934 & new_n10938 ;
  assign new_n10940 = ~new_n10369 & ~new_n10902 ;
  assign new_n10941 = ~new_n10939 & new_n10940 ;
  assign new_n10942 = ~new_n10907 & ~new_n10941 ;
  assign new_n10943 = ~new_n10904 & new_n10942 ;
  assign new_n10944 = ~new_n9692 & new_n10370 ;
  assign new_n10945 = ~new_n6812 & new_n10373 ;
  assign new_n10946 = ~new_n10372 & ~new_n10945 ;
  assign new_n10947 = ~new_n10944 & new_n10946 ;
  assign new_n10948 = ~new_n10362 & ~new_n10947 ;
  assign new_n10949 = new_n10362 & new_n10947 ;
  assign new_n10950 = ~new_n10948 & ~new_n10949 ;
  assign new_n10951 = ~new_n9035 & ~new_n10950 ;
  assign new_n10952 = new_n9035 & new_n10948 ;
  assign new_n10953 = ~new_n6720 & ~new_n6812 ;
  assign new_n10954 = new_n6720 & new_n6812 ;
  assign new_n10955 = ~new_n10953 & ~new_n10954 ;
  assign new_n10956 = ~new_n10393 & ~new_n10955 ;
  assign new_n10957 = new_n6720 & ~new_n6812 ;
  assign new_n10958 = ~new_n6720 & new_n6812 ;
  assign new_n10959 = ~new_n10957 & ~new_n10958 ;
  assign new_n10960 = ~new_n10956 & new_n10959 ;
  assign new_n10961 = new_n10394 & ~new_n10960 ;
  assign new_n10962 = new_n10400 & new_n10953 ;
  assign new_n10963 = ~new_n10961 & ~new_n10962 ;
  assign new_n10964 = new_n10393 & ~new_n10963 ;
  assign new_n10965 = ~new_n10393 & new_n10963 ;
  assign new_n10966 = ~new_n10964 & ~new_n10965 ;
  assign new_n10967 = ~new_n10392 & ~new_n10966 ;
  assign new_n10968 = new_n10392 & new_n10964 ;
  assign new_n10969 = new_n6812 & ~new_n10393 ;
  assign new_n10970 = ~new_n10963 & new_n10969 ;
  assign new_n10971 = ~new_n10968 & ~new_n10970 ;
  assign new_n10972 = ~new_n10967 & new_n10971 ;
  assign new_n10973 = new_n10389 & new_n10972 ;
  assign new_n10974 = ~new_n10414 & ~new_n10972 ;
  assign new_n10975 = new_n10416 & ~new_n10954 ;
  assign new_n10976 = ~new_n10974 & ~new_n10975 ;
  assign new_n10977 = ~new_n10973 & new_n10976 ;
  assign new_n10978 = ~new_n10388 & ~new_n10977 ;
  assign new_n10979 = new_n10388 & new_n10977 ;
  assign new_n10980 = ~new_n10978 & ~new_n10979 ;
  assign new_n10981 = ~new_n6720 & ~new_n10980 ;
  assign new_n10982 = new_n6720 & new_n10978 ;
  assign new_n10983 = new_n4619 & new_n10388 ;
  assign new_n10984 = ~new_n10977 & new_n10983 ;
  assign new_n10985 = ~new_n10982 & ~new_n10984 ;
  assign new_n10986 = ~new_n10981 & new_n10985 ;
  assign new_n10987 = new_n10362 & ~new_n10986 ;
  assign new_n10988 = ~new_n10947 & new_n10987 ;
  assign new_n10989 = ~new_n10952 & ~new_n10988 ;
  assign new_n10990 = ~new_n10951 & new_n10989 ;
  assign new_n10991 = ~new_n7037 & new_n10373 ;
  assign new_n10992 = ~new_n9159 & new_n10434 ;
  assign new_n10993 = ~new_n10372 & ~new_n10992 ;
  assign new_n10994 = ~new_n10991 & new_n10993 ;
  assign new_n10995 = new_n10369 & ~new_n10994 ;
  assign new_n10996 = new_n9699 & new_n10995 ;
  assign new_n10997 = ~new_n10369 & new_n10994 ;
  assign new_n10998 = ~new_n10995 & ~new_n10997 ;
  assign new_n10999 = ~new_n9699 & ~new_n10998 ;
  assign new_n11000 = new_n6945 & ~new_n7037 ;
  assign new_n11001 = ~new_n6945 & new_n7037 ;
  assign new_n11002 = ~new_n11000 & ~new_n11001 ;
  assign new_n11003 = ~new_n7037 & new_n10400 ;
  assign new_n11004 = ~new_n6945 & new_n11003 ;
  assign new_n11005 = new_n10542 & ~new_n11004 ;
  assign new_n11006 = new_n10394 & new_n11005 ;
  assign new_n11007 = ~new_n10394 & ~new_n11005 ;
  assign new_n11008 = ~new_n11006 & ~new_n11007 ;
  assign new_n11009 = ~new_n11002 & ~new_n11008 ;
  assign new_n11010 = new_n7037 & new_n10394 ;
  assign new_n11011 = ~new_n7037 & ~new_n10394 ;
  assign new_n11012 = ~new_n11010 & ~new_n11011 ;
  assign new_n11013 = ~new_n6945 & ~new_n11012 ;
  assign new_n11014 = new_n6945 & new_n7037 ;
  assign new_n11015 = ~new_n11013 & ~new_n11014 ;
  assign new_n11016 = ~new_n11005 & ~new_n11015 ;
  assign new_n11017 = ~new_n11009 & ~new_n11016 ;
  assign new_n11018 = new_n10389 & new_n11017 ;
  assign new_n11019 = ~new_n10414 & ~new_n11017 ;
  assign new_n11020 = new_n10416 & ~new_n11014 ;
  assign new_n11021 = ~new_n11019 & ~new_n11020 ;
  assign new_n11022 = ~new_n11018 & new_n11021 ;
  assign new_n11023 = ~new_n10388 & ~new_n11022 ;
  assign new_n11024 = new_n10388 & new_n11022 ;
  assign new_n11025 = ~new_n11023 & ~new_n11024 ;
  assign new_n11026 = ~new_n6945 & ~new_n11025 ;
  assign new_n11027 = new_n6945 & new_n11023 ;
  assign new_n11028 = new_n4981 & new_n10388 ;
  assign new_n11029 = ~new_n11022 & new_n11028 ;
  assign new_n11030 = ~new_n11027 & ~new_n11029 ;
  assign new_n11031 = ~new_n11026 & new_n11030 ;
  assign new_n11032 = ~new_n10369 & ~new_n10994 ;
  assign new_n11033 = ~new_n11031 & new_n11032 ;
  assign new_n11034 = ~new_n10999 & ~new_n11033 ;
  assign new_n11035 = ~new_n10996 & new_n11034 ;
  assign new_n11036 = ~new_n9706 & new_n10370 ;
  assign new_n11037 = ~new_n7260 & new_n10373 ;
  assign new_n11038 = ~new_n10372 & ~new_n11037 ;
  assign new_n11039 = ~new_n11036 & new_n11038 ;
  assign new_n11040 = ~new_n10362 & ~new_n11039 ;
  assign new_n11041 = new_n10362 & new_n11039 ;
  assign new_n11042 = ~new_n11040 & ~new_n11041 ;
  assign new_n11043 = ~new_n9283 & ~new_n11042 ;
  assign new_n11044 = new_n9283 & new_n11040 ;
  assign new_n11045 = ~new_n7168 & ~new_n7260 ;
  assign new_n11046 = new_n7168 & new_n7260 ;
  assign new_n11047 = ~new_n11045 & ~new_n11046 ;
  assign new_n11048 = ~new_n10393 & ~new_n11047 ;
  assign new_n11049 = new_n7168 & ~new_n7260 ;
  assign new_n11050 = ~new_n7168 & new_n7260 ;
  assign new_n11051 = ~new_n11049 & ~new_n11050 ;
  assign new_n11052 = ~new_n11048 & new_n11051 ;
  assign new_n11053 = new_n10394 & ~new_n11052 ;
  assign new_n11054 = new_n10400 & new_n11045 ;
  assign new_n11055 = ~new_n11053 & ~new_n11054 ;
  assign new_n11056 = new_n10393 & ~new_n11055 ;
  assign new_n11057 = ~new_n10393 & new_n11055 ;
  assign new_n11058 = ~new_n11056 & ~new_n11057 ;
  assign new_n11059 = ~new_n10392 & ~new_n11058 ;
  assign new_n11060 = new_n10392 & new_n11056 ;
  assign new_n11061 = new_n7260 & ~new_n10393 ;
  assign new_n11062 = ~new_n11055 & new_n11061 ;
  assign new_n11063 = ~new_n11060 & ~new_n11062 ;
  assign new_n11064 = ~new_n11059 & new_n11063 ;
  assign new_n11065 = new_n10389 & new_n11064 ;
  assign new_n11066 = ~new_n10414 & ~new_n11064 ;
  assign new_n11067 = new_n10416 & ~new_n11046 ;
  assign new_n11068 = ~new_n11066 & ~new_n11067 ;
  assign new_n11069 = ~new_n11065 & new_n11068 ;
  assign new_n11070 = ~new_n10388 & ~new_n11069 ;
  assign new_n11071 = new_n10388 & new_n11069 ;
  assign new_n11072 = ~new_n11070 & ~new_n11071 ;
  assign new_n11073 = ~new_n7168 & ~new_n11072 ;
  assign new_n11074 = new_n7168 & new_n11070 ;
  assign new_n11075 = new_n5265 & new_n10388 ;
  assign new_n11076 = ~new_n11069 & new_n11075 ;
  assign new_n11077 = ~new_n11074 & ~new_n11076 ;
  assign new_n11078 = ~new_n11073 & new_n11077 ;
  assign new_n11079 = new_n10362 & ~new_n11078 ;
  assign new_n11080 = ~new_n11039 & new_n11079 ;
  assign new_n11081 = ~new_n11044 & ~new_n11080 ;
  assign new_n11082 = ~new_n11043 & new_n11081 ;
  assign new_n11083 = ~lo0199 & ~new_n9720 ;
  assign new_n11084 = new_n3109 & ~new_n7423 ;
  assign new_n11085 = ~new_n3105 & new_n8013 ;
  assign new_n11086 = ~new_n10390 & ~new_n11085 ;
  assign new_n11087 = ~new_n11084 & new_n11086 ;
  assign new_n11088 = ~new_n11083 & new_n11087 ;
  assign new_n11089 = new_n3116 & ~new_n9720 ;
  assign new_n11090 = lo0198 & ~new_n7523 ;
  assign new_n11091 = ~new_n10391 & ~new_n11090 ;
  assign new_n11092 = ~lo0196 & ~lo0197 ;
  assign new_n11093 = ~new_n11091 & new_n11092 ;
  assign new_n11094 = ~new_n3099 & ~new_n11093 ;
  assign new_n11095 = ~new_n11089 & new_n11094 ;
  assign new_n11096 = ~lo0196 & ~new_n11095 ;
  assign new_n11097 = lo0196 & new_n11095 ;
  assign new_n11098 = ~new_n11096 & ~new_n11097 ;
  assign new_n11099 = ~new_n11088 & ~new_n11098 ;
  assign new_n11100 = new_n11088 & new_n11096 ;
  assign new_n11101 = lo0198 & new_n7523 ;
  assign new_n11102 = ~lo0198 & ~new_n7523 ;
  assign new_n11103 = ~new_n11101 & ~new_n11102 ;
  assign new_n11104 = ~lo0199 & ~new_n7423 ;
  assign new_n11105 = ~lo0199 & ~new_n11104 ;
  assign new_n11106 = ~new_n11103 & ~new_n11105 ;
  assign new_n11107 = ~lo0199 & new_n11090 ;
  assign new_n11108 = new_n7423 & new_n11107 ;
  assign new_n11109 = new_n7523 & new_n8013 ;
  assign new_n11110 = ~new_n7423 & new_n11109 ;
  assign new_n11111 = ~new_n11108 & ~new_n11110 ;
  assign new_n11112 = ~new_n11106 & new_n11111 ;
  assign new_n11113 = lo0196 & ~new_n11112 ;
  assign new_n11114 = ~new_n11095 & new_n11113 ;
  assign new_n11115 = ~new_n11100 & ~new_n11114 ;
  assign new_n11116 = ~new_n11099 & new_n11115 ;
  assign new_n11117 = lo0200 & ~new_n11116 ;
  assign new_n11118 = ~lo0199 & ~new_n3292 ;
  assign new_n11119 = lo0199 & ~new_n8551 ;
  assign new_n11120 = ~new_n11118 & ~new_n11119 ;
  assign new_n11121 = lo0196 & ~new_n9163 ;
  assign new_n11122 = ~new_n11120 & new_n11121 ;
  assign new_n11123 = ~new_n7423 & new_n9143 ;
  assign new_n11124 = lo0198 & new_n2899 ;
  assign new_n11125 = ~new_n11102 & ~new_n11124 ;
  assign new_n11126 = lo0199 & ~new_n11125 ;
  assign new_n11127 = ~new_n11123 & ~new_n11126 ;
  assign new_n11128 = ~lo0196 & ~new_n11127 ;
  assign new_n11129 = ~new_n11122 & ~new_n11128 ;
  assign new_n11130 = new_n3117 & ~new_n11129 ;
  assign new_n11131 = lo0196 & new_n9163 ;
  assign new_n11132 = new_n3117 & ~new_n11131 ;
  assign new_n11133 = ~new_n9720 & ~new_n11132 ;
  assign new_n11134 = ~new_n11130 & ~new_n11133 ;
  assign new_n11135 = ~lo0200 & ~new_n11134 ;
  assign new_n11136 = ~new_n11117 & ~new_n11135 ;
  assign new_n11137 = ~new_n7385 & new_n10373 ;
  assign new_n11138 = ~new_n9405 & new_n10434 ;
  assign new_n11139 = ~new_n10372 & ~new_n11138 ;
  assign new_n11140 = ~new_n11137 & new_n11139 ;
  assign new_n11141 = new_n10369 & ~new_n11140 ;
  assign new_n11142 = new_n9713 & new_n11141 ;
  assign new_n11143 = ~new_n10369 & new_n11140 ;
  assign new_n11144 = ~new_n11141 & ~new_n11143 ;
  assign new_n11145 = ~new_n9713 & ~new_n11144 ;
  assign new_n11146 = new_n7293 & ~new_n7385 ;
  assign new_n11147 = ~new_n7293 & new_n7385 ;
  assign new_n11148 = ~new_n11146 & ~new_n11147 ;
  assign new_n11149 = ~new_n7385 & new_n10400 ;
  assign new_n11150 = ~new_n7293 & new_n11149 ;
  assign new_n11151 = new_n10542 & ~new_n11150 ;
  assign new_n11152 = new_n10394 & new_n11151 ;
  assign new_n11153 = ~new_n10394 & ~new_n11151 ;
  assign new_n11154 = ~new_n11152 & ~new_n11153 ;
  assign new_n11155 = ~new_n11148 & ~new_n11154 ;
  assign new_n11156 = new_n7385 & new_n10394 ;
  assign new_n11157 = ~new_n7385 & ~new_n10394 ;
  assign new_n11158 = ~new_n11156 & ~new_n11157 ;
  assign new_n11159 = ~new_n7293 & ~new_n11158 ;
  assign new_n11160 = new_n7293 & new_n7385 ;
  assign new_n11161 = ~new_n11159 & ~new_n11160 ;
  assign new_n11162 = ~new_n11151 & ~new_n11161 ;
  assign new_n11163 = ~new_n11155 & ~new_n11162 ;
  assign new_n11164 = new_n10389 & new_n11163 ;
  assign new_n11165 = ~new_n10414 & ~new_n11163 ;
  assign new_n11166 = new_n10416 & ~new_n11160 ;
  assign new_n11167 = ~new_n11165 & ~new_n11166 ;
  assign new_n11168 = ~new_n11164 & new_n11167 ;
  assign new_n11169 = ~new_n10388 & ~new_n11168 ;
  assign new_n11170 = new_n10388 & new_n11168 ;
  assign new_n11171 = ~new_n11169 & ~new_n11170 ;
  assign new_n11172 = ~new_n7293 & ~new_n11171 ;
  assign new_n11173 = new_n7293 & new_n11169 ;
  assign new_n11174 = new_n5549 & new_n10388 ;
  assign new_n11175 = ~new_n11168 & new_n11174 ;
  assign new_n11176 = ~new_n11173 & ~new_n11175 ;
  assign new_n11177 = ~new_n11172 & new_n11176 ;
  assign new_n11178 = ~new_n10369 & ~new_n11140 ;
  assign new_n11179 = ~new_n11177 & new_n11178 ;
  assign new_n11180 = ~new_n11145 & ~new_n11179 ;
  assign new_n11181 = ~new_n11142 & new_n11180 ;
  assign new_n11182 = ~new_n9727 & ~new_n10232 ;
  assign new_n11183 = ~new_n3113 & ~new_n10259 ;
  assign new_n11184 = ~lo0197 & lo0198 ;
  assign new_n11185 = ~new_n10383 & ~new_n11184 ;
  assign new_n11186 = ~new_n11183 & ~new_n11185 ;
  assign new_n11187 = new_n10232 & new_n11186 ;
  assign new_n11188 = new_n7554 & new_n7648 ;
  assign new_n11189 = new_n11187 & ~new_n11188 ;
  assign new_n11190 = new_n10232 & ~new_n11186 ;
  assign new_n11191 = lo0198 & lo0200 ;
  assign new_n11192 = ~new_n10355 & ~new_n11191 ;
  assign new_n11193 = lo0199 & new_n11192 ;
  assign new_n11194 = ~new_n9267 & ~new_n11193 ;
  assign new_n11195 = lo0200 & new_n11193 ;
  assign new_n11196 = new_n11192 & ~new_n11195 ;
  assign new_n11197 = ~new_n11194 & ~new_n11196 ;
  assign new_n11198 = new_n7554 & new_n11197 ;
  assign new_n11199 = new_n11194 & new_n11196 ;
  assign new_n11200 = ~new_n11197 & ~new_n11199 ;
  assign new_n11201 = ~new_n7554 & ~new_n11200 ;
  assign new_n11202 = new_n11194 & ~new_n11196 ;
  assign new_n11203 = ~new_n7648 & new_n11202 ;
  assign new_n11204 = ~new_n11201 & ~new_n11203 ;
  assign new_n11205 = ~new_n11198 & new_n11204 ;
  assign new_n11206 = ~new_n11193 & ~new_n11205 ;
  assign new_n11207 = new_n11193 & new_n11205 ;
  assign new_n11208 = ~new_n11206 & ~new_n11207 ;
  assign new_n11209 = ~new_n3372 & ~new_n11208 ;
  assign new_n11210 = new_n3372 & new_n11206 ;
  assign new_n11211 = ~new_n8551 & new_n11193 ;
  assign new_n11212 = ~new_n11205 & new_n11211 ;
  assign new_n11213 = ~new_n11210 & ~new_n11212 ;
  assign new_n11214 = ~new_n11209 & new_n11213 ;
  assign new_n11215 = ~lo0197 & new_n11183 ;
  assign new_n11216 = ~new_n11214 & new_n11215 ;
  assign new_n11217 = lo0197 & ~new_n11183 ;
  assign new_n11218 = ~new_n7648 & new_n10237 ;
  assign new_n11219 = ~new_n7554 & new_n11218 ;
  assign new_n11220 = ~new_n3650 & new_n10241 ;
  assign new_n11221 = ~new_n10240 & ~new_n11220 ;
  assign new_n11222 = ~new_n11219 & new_n11221 ;
  assign new_n11223 = new_n10236 & ~new_n11222 ;
  assign new_n11224 = ~new_n10236 & new_n11222 ;
  assign new_n11225 = ~new_n11223 & ~new_n11224 ;
  assign new_n11226 = ~new_n8672 & ~new_n11225 ;
  assign new_n11227 = new_n8672 & new_n11223 ;
  assign new_n11228 = ~new_n7554 & new_n7648 ;
  assign new_n11229 = new_n7554 & ~new_n7648 ;
  assign new_n11230 = ~new_n11228 & ~new_n11229 ;
  assign new_n11231 = ~new_n10236 & ~new_n11230 ;
  assign new_n11232 = ~new_n11222 & new_n11231 ;
  assign new_n11233 = ~new_n11227 & ~new_n11232 ;
  assign new_n11234 = ~new_n11226 & new_n11233 ;
  assign new_n11235 = lo0197 & new_n11183 ;
  assign new_n11236 = ~new_n11234 & new_n11235 ;
  assign new_n11237 = ~new_n11217 & ~new_n11236 ;
  assign new_n11238 = ~new_n11216 & new_n11237 ;
  assign new_n11239 = new_n11183 & ~new_n11238 ;
  assign new_n11240 = ~new_n11183 & new_n11238 ;
  assign new_n11241 = ~new_n11239 & ~new_n11240 ;
  assign new_n11242 = ~new_n3557 & ~new_n11241 ;
  assign new_n11243 = new_n3557 & new_n11239 ;
  assign new_n11244 = new_n7648 & ~new_n11183 ;
  assign new_n11245 = ~new_n11238 & new_n11244 ;
  assign new_n11246 = ~new_n11243 & ~new_n11245 ;
  assign new_n11247 = ~new_n11242 & new_n11246 ;
  assign new_n11248 = new_n11190 & ~new_n11247 ;
  assign new_n11249 = ~new_n11189 & ~new_n11248 ;
  assign new_n11250 = ~new_n11182 & new_n11249 ;
  assign new_n11251 = ~new_n9734 & ~new_n10232 ;
  assign new_n11252 = new_n7678 & new_n7772 ;
  assign new_n11253 = new_n11187 & ~new_n11252 ;
  assign new_n11254 = new_n7678 & new_n11197 ;
  assign new_n11255 = ~new_n7678 & ~new_n11200 ;
  assign new_n11256 = ~new_n7772 & new_n11202 ;
  assign new_n11257 = ~new_n11255 & ~new_n11256 ;
  assign new_n11258 = ~new_n11254 & new_n11257 ;
  assign new_n11259 = ~new_n11193 & ~new_n11258 ;
  assign new_n11260 = new_n11193 & new_n11258 ;
  assign new_n11261 = ~new_n11259 & ~new_n11260 ;
  assign new_n11262 = ~new_n3723 & ~new_n11261 ;
  assign new_n11263 = new_n3723 & new_n11259 ;
  assign new_n11264 = new_n11211 & ~new_n11258 ;
  assign new_n11265 = ~new_n11263 & ~new_n11264 ;
  assign new_n11266 = ~new_n11262 & new_n11265 ;
  assign new_n11267 = new_n11215 & ~new_n11266 ;
  assign new_n11268 = ~new_n4014 & new_n10241 ;
  assign new_n11269 = ~new_n10234 & ~new_n10236 ;
  assign new_n11270 = ~new_n8794 & new_n11269 ;
  assign new_n11271 = ~new_n10240 & ~new_n11270 ;
  assign new_n11272 = ~new_n11268 & new_n11271 ;
  assign new_n11273 = ~new_n7678 & ~new_n7772 ;
  assign new_n11274 = ~new_n11252 & ~new_n11273 ;
  assign new_n11275 = ~new_n10234 & ~new_n11274 ;
  assign new_n11276 = new_n7678 & ~new_n7772 ;
  assign new_n11277 = ~new_n7678 & new_n7772 ;
  assign new_n11278 = ~new_n11276 & ~new_n11277 ;
  assign new_n11279 = ~new_n11275 & new_n11278 ;
  assign new_n11280 = ~new_n11272 & ~new_n11279 ;
  assign new_n11281 = new_n10234 & new_n11272 ;
  assign new_n11282 = new_n11273 & new_n11281 ;
  assign new_n11283 = ~new_n11280 & ~new_n11282 ;
  assign new_n11284 = new_n11235 & ~new_n11283 ;
  assign new_n11285 = ~new_n11217 & ~new_n11284 ;
  assign new_n11286 = ~new_n11267 & new_n11285 ;
  assign new_n11287 = new_n11183 & ~new_n11286 ;
  assign new_n11288 = ~new_n11183 & new_n11286 ;
  assign new_n11289 = ~new_n11287 & ~new_n11288 ;
  assign new_n11290 = ~new_n3922 & ~new_n11289 ;
  assign new_n11291 = new_n3922 & new_n11287 ;
  assign new_n11292 = new_n7772 & ~new_n11183 ;
  assign new_n11293 = ~new_n11286 & new_n11292 ;
  assign new_n11294 = ~new_n11291 & ~new_n11293 ;
  assign new_n11295 = ~new_n11290 & new_n11294 ;
  assign new_n11296 = new_n11190 & ~new_n11295 ;
  assign new_n11297 = ~new_n11253 & ~new_n11296 ;
  assign new_n11298 = ~new_n11251 & new_n11297 ;
  assign new_n11299 = ~new_n9741 & ~new_n10232 ;
  assign new_n11300 = new_n7802 & new_n7894 ;
  assign new_n11301 = new_n11187 & ~new_n11300 ;
  assign new_n11302 = new_n7802 & new_n11197 ;
  assign new_n11303 = ~new_n7802 & ~new_n11200 ;
  assign new_n11304 = ~new_n7894 & new_n11202 ;
  assign new_n11305 = ~new_n11303 & ~new_n11304 ;
  assign new_n11306 = ~new_n11302 & new_n11305 ;
  assign new_n11307 = ~new_n11193 & ~new_n11306 ;
  assign new_n11308 = new_n11193 & new_n11306 ;
  assign new_n11309 = ~new_n11307 & ~new_n11308 ;
  assign new_n11310 = ~new_n4168 & ~new_n11309 ;
  assign new_n11311 = new_n4168 & new_n11307 ;
  assign new_n11312 = new_n11211 & ~new_n11306 ;
  assign new_n11313 = ~new_n11311 & ~new_n11312 ;
  assign new_n11314 = ~new_n11310 & new_n11313 ;
  assign new_n11315 = new_n11215 & ~new_n11314 ;
  assign new_n11316 = ~new_n7894 & new_n10237 ;
  assign new_n11317 = ~new_n7802 & new_n11316 ;
  assign new_n11318 = ~new_n4373 & new_n10241 ;
  assign new_n11319 = ~new_n10240 & ~new_n11318 ;
  assign new_n11320 = ~new_n11317 & new_n11319 ;
  assign new_n11321 = new_n10236 & ~new_n11320 ;
  assign new_n11322 = ~new_n10236 & new_n11320 ;
  assign new_n11323 = ~new_n11321 & ~new_n11322 ;
  assign new_n11324 = ~new_n8915 & ~new_n11323 ;
  assign new_n11325 = new_n8915 & new_n11321 ;
  assign new_n11326 = ~new_n7802 & new_n7894 ;
  assign new_n11327 = new_n7802 & ~new_n7894 ;
  assign new_n11328 = ~new_n11326 & ~new_n11327 ;
  assign new_n11329 = ~new_n10236 & ~new_n11328 ;
  assign new_n11330 = ~new_n11320 & new_n11329 ;
  assign new_n11331 = ~new_n11325 & ~new_n11330 ;
  assign new_n11332 = ~new_n11324 & new_n11331 ;
  assign new_n11333 = new_n11235 & ~new_n11332 ;
  assign new_n11334 = ~new_n11217 & ~new_n11333 ;
  assign new_n11335 = ~new_n11315 & new_n11334 ;
  assign new_n11336 = new_n11183 & ~new_n11335 ;
  assign new_n11337 = ~new_n11183 & new_n11335 ;
  assign new_n11338 = ~new_n11336 & ~new_n11337 ;
  assign new_n11339 = ~new_n4281 & ~new_n11338 ;
  assign new_n11340 = new_n4281 & new_n11336 ;
  assign new_n11341 = new_n7894 & ~new_n11183 ;
  assign new_n11342 = ~new_n11335 & new_n11341 ;
  assign new_n11343 = ~new_n11340 & ~new_n11342 ;
  assign new_n11344 = ~new_n11339 & new_n11343 ;
  assign new_n11345 = new_n11190 & ~new_n11344 ;
  assign new_n11346 = ~new_n11301 & ~new_n11345 ;
  assign new_n11347 = ~new_n11299 & new_n11346 ;
  assign new_n11348 = ~new_n9748 & ~new_n10232 ;
  assign new_n11349 = new_n7926 & new_n8035 ;
  assign new_n11350 = new_n11187 & ~new_n11349 ;
  assign new_n11351 = new_n7926 & new_n11197 ;
  assign new_n11352 = ~new_n7926 & ~new_n11200 ;
  assign new_n11353 = ~new_n8035 & new_n11202 ;
  assign new_n11354 = ~new_n11352 & ~new_n11353 ;
  assign new_n11355 = ~new_n11351 & new_n11354 ;
  assign new_n11356 = ~new_n11193 & ~new_n11355 ;
  assign new_n11357 = new_n11193 & new_n11355 ;
  assign new_n11358 = ~new_n11356 & ~new_n11357 ;
  assign new_n11359 = ~new_n4446 & ~new_n11358 ;
  assign new_n11360 = new_n4446 & new_n11356 ;
  assign new_n11361 = new_n11211 & ~new_n11355 ;
  assign new_n11362 = ~new_n11360 & ~new_n11361 ;
  assign new_n11363 = ~new_n11359 & new_n11362 ;
  assign new_n11364 = new_n11215 & ~new_n11363 ;
  assign new_n11365 = ~new_n4735 & new_n10241 ;
  assign new_n11366 = ~new_n9035 & new_n11269 ;
  assign new_n11367 = ~new_n10240 & ~new_n11366 ;
  assign new_n11368 = ~new_n11365 & new_n11367 ;
  assign new_n11369 = ~new_n7926 & ~new_n8035 ;
  assign new_n11370 = ~new_n11349 & ~new_n11369 ;
  assign new_n11371 = ~new_n10234 & ~new_n11370 ;
  assign new_n11372 = new_n7926 & ~new_n8035 ;
  assign new_n11373 = ~new_n7926 & new_n8035 ;
  assign new_n11374 = ~new_n11372 & ~new_n11373 ;
  assign new_n11375 = ~new_n11371 & new_n11374 ;
  assign new_n11376 = ~new_n11368 & ~new_n11375 ;
  assign new_n11377 = new_n10234 & new_n11368 ;
  assign new_n11378 = new_n11369 & new_n11377 ;
  assign new_n11379 = ~new_n11376 & ~new_n11378 ;
  assign new_n11380 = new_n11235 & ~new_n11379 ;
  assign new_n11381 = ~new_n11217 & ~new_n11380 ;
  assign new_n11382 = ~new_n11364 & new_n11381 ;
  assign new_n11383 = new_n11183 & ~new_n11382 ;
  assign new_n11384 = ~new_n11183 & new_n11382 ;
  assign new_n11385 = ~new_n11383 & ~new_n11384 ;
  assign new_n11386 = ~new_n4643 & ~new_n11385 ;
  assign new_n11387 = new_n4643 & new_n11383 ;
  assign new_n11388 = new_n8035 & ~new_n11183 ;
  assign new_n11389 = ~new_n11382 & new_n11388 ;
  assign new_n11390 = ~new_n11387 & ~new_n11389 ;
  assign new_n11391 = ~new_n11386 & new_n11390 ;
  assign new_n11392 = new_n11190 & ~new_n11391 ;
  assign new_n11393 = ~new_n11350 & ~new_n11392 ;
  assign new_n11394 = ~new_n11348 & new_n11393 ;
  assign new_n11395 = ~new_n9755 & ~new_n10232 ;
  assign new_n11396 = new_n8067 & new_n8163 ;
  assign new_n11397 = new_n11187 & ~new_n11396 ;
  assign new_n11398 = new_n8067 & new_n11197 ;
  assign new_n11399 = ~new_n8067 & ~new_n11200 ;
  assign new_n11400 = ~new_n8163 & new_n11202 ;
  assign new_n11401 = ~new_n11399 & ~new_n11400 ;
  assign new_n11402 = ~new_n11398 & new_n11401 ;
  assign new_n11403 = ~new_n11193 & ~new_n11402 ;
  assign new_n11404 = new_n11193 & new_n11402 ;
  assign new_n11405 = ~new_n11403 & ~new_n11404 ;
  assign new_n11406 = ~new_n4889 & ~new_n11405 ;
  assign new_n11407 = new_n4889 & new_n11403 ;
  assign new_n11408 = new_n11211 & ~new_n11402 ;
  assign new_n11409 = ~new_n11407 & ~new_n11408 ;
  assign new_n11410 = ~new_n11406 & new_n11409 ;
  assign new_n11411 = new_n11215 & ~new_n11410 ;
  assign new_n11412 = ~new_n8163 & new_n10237 ;
  assign new_n11413 = ~new_n8067 & new_n11412 ;
  assign new_n11414 = ~new_n5097 & new_n10241 ;
  assign new_n11415 = ~new_n10240 & ~new_n11414 ;
  assign new_n11416 = ~new_n11413 & new_n11415 ;
  assign new_n11417 = new_n10236 & ~new_n11416 ;
  assign new_n11418 = ~new_n10236 & new_n11416 ;
  assign new_n11419 = ~new_n11417 & ~new_n11418 ;
  assign new_n11420 = ~new_n9159 & ~new_n11419 ;
  assign new_n11421 = new_n9159 & new_n11417 ;
  assign new_n11422 = ~new_n8067 & new_n8163 ;
  assign new_n11423 = new_n8067 & ~new_n8163 ;
  assign new_n11424 = ~new_n11422 & ~new_n11423 ;
  assign new_n11425 = ~new_n10236 & ~new_n11424 ;
  assign new_n11426 = ~new_n11416 & new_n11425 ;
  assign new_n11427 = ~new_n11421 & ~new_n11426 ;
  assign new_n11428 = ~new_n11420 & new_n11427 ;
  assign new_n11429 = new_n11235 & ~new_n11428 ;
  assign new_n11430 = ~new_n11217 & ~new_n11429 ;
  assign new_n11431 = ~new_n11411 & new_n11430 ;
  assign new_n11432 = new_n11183 & ~new_n11431 ;
  assign new_n11433 = ~new_n11183 & new_n11431 ;
  assign new_n11434 = ~new_n11432 & ~new_n11433 ;
  assign new_n11435 = ~new_n5005 & ~new_n11434 ;
  assign new_n11436 = new_n5005 & new_n11432 ;
  assign new_n11437 = new_n8163 & ~new_n11183 ;
  assign new_n11438 = ~new_n11431 & new_n11437 ;
  assign new_n11439 = ~new_n11436 & ~new_n11438 ;
  assign new_n11440 = ~new_n11435 & new_n11439 ;
  assign new_n11441 = new_n11190 & ~new_n11440 ;
  assign new_n11442 = ~new_n11397 & ~new_n11441 ;
  assign new_n11443 = ~new_n11395 & new_n11442 ;
  assign new_n11444 = ~new_n9762 & ~new_n10232 ;
  assign new_n11445 = new_n8195 & new_n8295 ;
  assign new_n11446 = new_n11187 & ~new_n11445 ;
  assign new_n11447 = new_n8195 & new_n11197 ;
  assign new_n11448 = ~new_n8195 & ~new_n11200 ;
  assign new_n11449 = ~new_n8295 & new_n11202 ;
  assign new_n11450 = ~new_n11448 & ~new_n11449 ;
  assign new_n11451 = ~new_n11447 & new_n11450 ;
  assign new_n11452 = ~new_n11193 & ~new_n11451 ;
  assign new_n11453 = new_n11193 & new_n11451 ;
  assign new_n11454 = ~new_n11452 & ~new_n11453 ;
  assign new_n11455 = ~new_n5170 & ~new_n11454 ;
  assign new_n11456 = new_n5170 & new_n11452 ;
  assign new_n11457 = new_n11211 & ~new_n11451 ;
  assign new_n11458 = ~new_n11456 & ~new_n11457 ;
  assign new_n11459 = ~new_n11455 & new_n11458 ;
  assign new_n11460 = new_n11215 & ~new_n11459 ;
  assign new_n11461 = ~new_n5381 & new_n10241 ;
  assign new_n11462 = ~new_n9283 & new_n11269 ;
  assign new_n11463 = ~new_n10240 & ~new_n11462 ;
  assign new_n11464 = ~new_n11461 & new_n11463 ;
  assign new_n11465 = ~new_n8195 & ~new_n8295 ;
  assign new_n11466 = ~new_n11445 & ~new_n11465 ;
  assign new_n11467 = ~new_n10234 & ~new_n11466 ;
  assign new_n11468 = new_n8195 & ~new_n8295 ;
  assign new_n11469 = ~new_n8195 & new_n8295 ;
  assign new_n11470 = ~new_n11468 & ~new_n11469 ;
  assign new_n11471 = ~new_n11467 & new_n11470 ;
  assign new_n11472 = ~new_n11464 & ~new_n11471 ;
  assign new_n11473 = new_n10234 & new_n11464 ;
  assign new_n11474 = new_n11465 & new_n11473 ;
  assign new_n11475 = ~new_n11472 & ~new_n11474 ;
  assign new_n11476 = new_n11235 & ~new_n11475 ;
  assign new_n11477 = ~new_n11217 & ~new_n11476 ;
  assign new_n11478 = ~new_n11460 & new_n11477 ;
  assign new_n11479 = new_n11183 & ~new_n11478 ;
  assign new_n11480 = ~new_n11183 & new_n11478 ;
  assign new_n11481 = ~new_n11479 & ~new_n11480 ;
  assign new_n11482 = ~new_n5289 & ~new_n11481 ;
  assign new_n11483 = new_n5289 & new_n11479 ;
  assign new_n11484 = new_n8295 & ~new_n11183 ;
  assign new_n11485 = ~new_n11478 & new_n11484 ;
  assign new_n11486 = ~new_n11483 & ~new_n11485 ;
  assign new_n11487 = ~new_n11482 & new_n11486 ;
  assign new_n11488 = new_n11190 & ~new_n11487 ;
  assign new_n11489 = ~new_n11446 & ~new_n11488 ;
  assign new_n11490 = ~new_n11444 & new_n11489 ;
  assign new_n11491 = ~new_n9769 & ~new_n10232 ;
  assign new_n11492 = new_n8327 & new_n8425 ;
  assign new_n11493 = new_n11187 & ~new_n11492 ;
  assign new_n11494 = new_n8327 & new_n11197 ;
  assign new_n11495 = ~new_n8327 & ~new_n11200 ;
  assign new_n11496 = ~new_n8425 & new_n11202 ;
  assign new_n11497 = ~new_n11495 & ~new_n11496 ;
  assign new_n11498 = ~new_n11494 & new_n11497 ;
  assign new_n11499 = ~new_n11193 & ~new_n11498 ;
  assign new_n11500 = new_n11193 & new_n11498 ;
  assign new_n11501 = ~new_n11499 & ~new_n11500 ;
  assign new_n11502 = ~new_n5455 & ~new_n11501 ;
  assign new_n11503 = new_n5455 & new_n11499 ;
  assign new_n11504 = new_n11211 & ~new_n11498 ;
  assign new_n11505 = ~new_n11503 & ~new_n11504 ;
  assign new_n11506 = ~new_n11502 & new_n11505 ;
  assign new_n11507 = new_n11215 & ~new_n11506 ;
  assign new_n11508 = ~new_n8425 & new_n10237 ;
  assign new_n11509 = ~new_n8327 & new_n11508 ;
  assign new_n11510 = ~new_n5665 & new_n10241 ;
  assign new_n11511 = ~new_n10240 & ~new_n11510 ;
  assign new_n11512 = ~new_n11509 & new_n11511 ;
  assign new_n11513 = new_n10236 & ~new_n11512 ;
  assign new_n11514 = ~new_n10236 & new_n11512 ;
  assign new_n11515 = ~new_n11513 & ~new_n11514 ;
  assign new_n11516 = ~new_n9405 & ~new_n11515 ;
  assign new_n11517 = new_n9405 & new_n11513 ;
  assign new_n11518 = new_n8327 & ~new_n8425 ;
  assign new_n11519 = ~new_n8327 & new_n8425 ;
  assign new_n11520 = ~new_n11518 & ~new_n11519 ;
  assign new_n11521 = ~new_n10236 & ~new_n11520 ;
  assign new_n11522 = ~new_n11512 & new_n11521 ;
  assign new_n11523 = ~new_n11517 & ~new_n11522 ;
  assign new_n11524 = ~new_n11516 & new_n11523 ;
  assign new_n11525 = new_n11235 & ~new_n11524 ;
  assign new_n11526 = ~new_n11217 & ~new_n11525 ;
  assign new_n11527 = ~new_n11507 & new_n11526 ;
  assign new_n11528 = new_n11183 & ~new_n11527 ;
  assign new_n11529 = ~new_n11183 & new_n11527 ;
  assign new_n11530 = ~new_n11528 & ~new_n11529 ;
  assign new_n11531 = ~new_n5573 & ~new_n11530 ;
  assign new_n11532 = new_n5573 & new_n11528 ;
  assign new_n11533 = new_n8425 & ~new_n11183 ;
  assign new_n11534 = ~new_n11527 & new_n11533 ;
  assign new_n11535 = ~new_n11532 & ~new_n11534 ;
  assign new_n11536 = ~new_n11531 & new_n11535 ;
  assign new_n11537 = new_n11190 & ~new_n11536 ;
  assign new_n11538 = ~new_n11493 & ~new_n11537 ;
  assign new_n11539 = ~new_n11491 & new_n11538 ;
  assign new_n11540 = ~new_n9776 & ~new_n10232 ;
  assign new_n11541 = ~new_n5799 & new_n10267 ;
  assign new_n11542 = ~new_n8551 & ~new_n10271 ;
  assign new_n11543 = new_n8551 & new_n10269 ;
  assign new_n11544 = ~new_n11542 & ~new_n11543 ;
  assign new_n11545 = ~new_n11541 & new_n11544 ;
  assign new_n11546 = ~new_n10263 & ~new_n11545 ;
  assign new_n11547 = new_n10263 & new_n11545 ;
  assign new_n11548 = ~new_n11546 & ~new_n11547 ;
  assign new_n11549 = ~new_n8449 & ~new_n11548 ;
  assign new_n11550 = new_n8449 & new_n11546 ;
  assign new_n11551 = ~new_n5743 & new_n10263 ;
  assign new_n11552 = ~new_n11545 & new_n11551 ;
  assign new_n11553 = ~new_n11550 & ~new_n11552 ;
  assign new_n11554 = ~new_n11549 & new_n11553 ;
  assign new_n11555 = new_n10261 & ~new_n11554 ;
  assign new_n11556 = new_n10258 & new_n10260 ;
  assign new_n11557 = ~new_n5891 & new_n10241 ;
  assign new_n11558 = ~new_n7523 & new_n11269 ;
  assign new_n11559 = ~new_n10240 & ~new_n11558 ;
  assign new_n11560 = ~new_n11557 & new_n11559 ;
  assign new_n11561 = ~new_n8449 & ~new_n8551 ;
  assign new_n11562 = new_n8449 & new_n8551 ;
  assign new_n11563 = ~new_n11561 & ~new_n11562 ;
  assign new_n11564 = ~new_n10234 & ~new_n11563 ;
  assign new_n11565 = new_n8449 & ~new_n8551 ;
  assign new_n11566 = ~new_n8449 & new_n8551 ;
  assign new_n11567 = ~new_n11565 & ~new_n11566 ;
  assign new_n11568 = ~new_n11564 & new_n11567 ;
  assign new_n11569 = ~new_n11560 & ~new_n11568 ;
  assign new_n11570 = new_n10234 & new_n11560 ;
  assign new_n11571 = new_n11561 & new_n11570 ;
  assign new_n11572 = ~new_n11569 & ~new_n11571 ;
  assign new_n11573 = new_n11556 & ~new_n11572 ;
  assign new_n11574 = ~new_n10286 & ~new_n11573 ;
  assign new_n11575 = ~new_n11555 & new_n11574 ;
  assign new_n11576 = new_n8551 & ~new_n11575 ;
  assign new_n11577 = ~new_n8551 & new_n11575 ;
  assign new_n11578 = ~new_n11576 & ~new_n11577 ;
  assign new_n11579 = new_n8449 & ~new_n11578 ;
  assign new_n11580 = ~new_n8449 & new_n11576 ;
  assign new_n11581 = ~new_n11579 & ~new_n11580 ;
  assign new_n11582 = ~new_n10260 & ~new_n11581 ;
  assign new_n11583 = ~new_n10260 & new_n11575 ;
  assign new_n11584 = new_n10260 & ~new_n11575 ;
  assign new_n11585 = ~new_n11583 & ~new_n11584 ;
  assign new_n11586 = ~new_n8449 & ~new_n11585 ;
  assign new_n11587 = new_n8449 & new_n11584 ;
  assign new_n11588 = ~new_n11586 & ~new_n11587 ;
  assign new_n11589 = ~new_n11582 & new_n11588 ;
  assign new_n11590 = new_n10232 & ~new_n11589 ;
  assign new_n11591 = ~new_n11540 & ~new_n11590 ;
  assign new_n11592 = ~new_n9783 & ~new_n10232 ;
  assign new_n11593 = ~new_n8672 & new_n10237 ;
  assign new_n11594 = ~new_n8575 & new_n11593 ;
  assign new_n11595 = ~new_n6117 & new_n10241 ;
  assign new_n11596 = ~new_n10240 & ~new_n11595 ;
  assign new_n11597 = ~new_n11594 & new_n11596 ;
  assign new_n11598 = new_n10236 & ~new_n11597 ;
  assign new_n11599 = ~new_n10236 & new_n11597 ;
  assign new_n11600 = ~new_n11598 & ~new_n11599 ;
  assign new_n11601 = ~new_n7648 & ~new_n11600 ;
  assign new_n11602 = new_n7648 & new_n11598 ;
  assign new_n11603 = ~new_n8575 & new_n8672 ;
  assign new_n11604 = new_n8575 & ~new_n8672 ;
  assign new_n11605 = ~new_n11603 & ~new_n11604 ;
  assign new_n11606 = ~new_n10236 & ~new_n11605 ;
  assign new_n11607 = ~new_n11597 & new_n11606 ;
  assign new_n11608 = ~new_n11602 & ~new_n11607 ;
  assign new_n11609 = ~new_n11601 & new_n11608 ;
  assign new_n11610 = ~new_n6025 & new_n10267 ;
  assign new_n11611 = ~new_n8672 & ~new_n10271 ;
  assign new_n11612 = new_n8672 & new_n10269 ;
  assign new_n11613 = ~new_n11611 & ~new_n11612 ;
  assign new_n11614 = ~new_n11610 & new_n11613 ;
  assign new_n11615 = ~new_n10263 & ~new_n11614 ;
  assign new_n11616 = new_n10263 & new_n11614 ;
  assign new_n11617 = ~new_n11615 & ~new_n11616 ;
  assign new_n11618 = ~new_n8575 & ~new_n11617 ;
  assign new_n11619 = new_n8575 & new_n11615 ;
  assign new_n11620 = new_n5977 & new_n10263 ;
  assign new_n11621 = ~new_n11614 & new_n11620 ;
  assign new_n11622 = ~new_n11619 & ~new_n11621 ;
  assign new_n11623 = ~new_n11618 & new_n11622 ;
  assign new_n11624 = new_n10261 & ~new_n11623 ;
  assign new_n11625 = new_n8575 & new_n8672 ;
  assign new_n11626 = new_n10287 & ~new_n11625 ;
  assign new_n11627 = ~new_n10286 & ~new_n11626 ;
  assign new_n11628 = ~new_n11624 & new_n11627 ;
  assign new_n11629 = ~new_n10258 & ~new_n11628 ;
  assign new_n11630 = new_n10258 & new_n11628 ;
  assign new_n11631 = ~new_n11629 & ~new_n11630 ;
  assign new_n11632 = ~new_n11609 & ~new_n11631 ;
  assign new_n11633 = new_n11609 & new_n11629 ;
  assign new_n11634 = new_n8672 & new_n10258 ;
  assign new_n11635 = ~new_n11628 & new_n11634 ;
  assign new_n11636 = ~new_n11633 & ~new_n11635 ;
  assign new_n11637 = ~new_n11632 & new_n11636 ;
  assign new_n11638 = new_n10232 & ~new_n11637 ;
  assign new_n11639 = ~new_n11592 & ~new_n11638 ;
  assign new_n11640 = ~new_n9790 & ~new_n10232 ;
  assign new_n11641 = ~new_n6255 & new_n10267 ;
  assign new_n11642 = ~new_n8794 & ~new_n10271 ;
  assign new_n11643 = new_n8794 & new_n10269 ;
  assign new_n11644 = ~new_n11642 & ~new_n11643 ;
  assign new_n11645 = ~new_n11641 & new_n11644 ;
  assign new_n11646 = ~new_n10263 & ~new_n11645 ;
  assign new_n11647 = new_n10263 & new_n11645 ;
  assign new_n11648 = ~new_n11646 & ~new_n11647 ;
  assign new_n11649 = ~new_n8696 & ~new_n11648 ;
  assign new_n11650 = new_n8696 & new_n11646 ;
  assign new_n11651 = new_n6202 & new_n10263 ;
  assign new_n11652 = ~new_n11645 & new_n11651 ;
  assign new_n11653 = ~new_n11650 & ~new_n11652 ;
  assign new_n11654 = ~new_n11649 & new_n11653 ;
  assign new_n11655 = new_n10261 & ~new_n11654 ;
  assign new_n11656 = ~new_n6347 & new_n10241 ;
  assign new_n11657 = ~new_n7772 & new_n11269 ;
  assign new_n11658 = ~new_n10240 & ~new_n11657 ;
  assign new_n11659 = ~new_n11656 & new_n11658 ;
  assign new_n11660 = ~new_n8696 & ~new_n8794 ;
  assign new_n11661 = new_n8696 & new_n8794 ;
  assign new_n11662 = ~new_n11660 & ~new_n11661 ;
  assign new_n11663 = ~new_n10234 & ~new_n11662 ;
  assign new_n11664 = ~new_n8696 & new_n8794 ;
  assign new_n11665 = new_n8696 & ~new_n8794 ;
  assign new_n11666 = ~new_n11664 & ~new_n11665 ;
  assign new_n11667 = ~new_n11663 & new_n11666 ;
  assign new_n11668 = ~new_n11659 & ~new_n11667 ;
  assign new_n11669 = new_n10234 & new_n11659 ;
  assign new_n11670 = new_n11660 & new_n11669 ;
  assign new_n11671 = ~new_n11668 & ~new_n11670 ;
  assign new_n11672 = new_n11556 & ~new_n11671 ;
  assign new_n11673 = ~new_n10286 & ~new_n11672 ;
  assign new_n11674 = ~new_n11655 & new_n11673 ;
  assign new_n11675 = new_n8794 & ~new_n11674 ;
  assign new_n11676 = ~new_n8794 & new_n11674 ;
  assign new_n11677 = ~new_n11675 & ~new_n11676 ;
  assign new_n11678 = new_n8696 & ~new_n11677 ;
  assign new_n11679 = ~new_n8696 & new_n11675 ;
  assign new_n11680 = ~new_n11678 & ~new_n11679 ;
  assign new_n11681 = ~new_n10260 & ~new_n11680 ;
  assign new_n11682 = ~new_n10260 & new_n11674 ;
  assign new_n11683 = new_n10260 & ~new_n11674 ;
  assign new_n11684 = ~new_n11682 & ~new_n11683 ;
  assign new_n11685 = ~new_n8696 & ~new_n11684 ;
  assign new_n11686 = new_n8696 & new_n11683 ;
  assign new_n11687 = ~new_n11685 & ~new_n11686 ;
  assign new_n11688 = ~new_n11681 & new_n11687 ;
  assign new_n11689 = new_n10232 & ~new_n11688 ;
  assign new_n11690 = ~new_n11640 & ~new_n11689 ;
  assign new_n11691 = ~new_n9818 & ~new_n10232 ;
  assign new_n11692 = ~new_n7168 & new_n10267 ;
  assign new_n11693 = ~new_n9283 & ~new_n10271 ;
  assign new_n11694 = new_n9283 & new_n10269 ;
  assign new_n11695 = ~new_n11693 & ~new_n11694 ;
  assign new_n11696 = ~new_n11692 & new_n11695 ;
  assign new_n11697 = ~new_n10263 & ~new_n11696 ;
  assign new_n11698 = new_n10263 & new_n11696 ;
  assign new_n11699 = ~new_n11697 & ~new_n11698 ;
  assign new_n11700 = ~new_n9182 & ~new_n11699 ;
  assign new_n11701 = new_n9182 & new_n11697 ;
  assign new_n11702 = new_n7122 & new_n10263 ;
  assign new_n11703 = ~new_n11696 & new_n11702 ;
  assign new_n11704 = ~new_n11701 & ~new_n11703 ;
  assign new_n11705 = ~new_n11700 & new_n11704 ;
  assign new_n11706 = new_n10261 & ~new_n11705 ;
  assign new_n11707 = ~new_n7260 & new_n10241 ;
  assign new_n11708 = ~new_n8295 & new_n11269 ;
  assign new_n11709 = ~new_n10240 & ~new_n11708 ;
  assign new_n11710 = ~new_n11707 & new_n11709 ;
  assign new_n11711 = ~new_n9182 & ~new_n9283 ;
  assign new_n11712 = new_n9182 & new_n9283 ;
  assign new_n11713 = ~new_n11711 & ~new_n11712 ;
  assign new_n11714 = ~new_n10234 & ~new_n11713 ;
  assign new_n11715 = ~new_n9182 & new_n9283 ;
  assign new_n11716 = new_n9182 & ~new_n9283 ;
  assign new_n11717 = ~new_n11715 & ~new_n11716 ;
  assign new_n11718 = ~new_n11714 & new_n11717 ;
  assign new_n11719 = ~new_n11710 & ~new_n11718 ;
  assign new_n11720 = new_n10234 & new_n11710 ;
  assign new_n11721 = new_n11711 & new_n11720 ;
  assign new_n11722 = ~new_n11719 & ~new_n11721 ;
  assign new_n11723 = new_n11556 & ~new_n11722 ;
  assign new_n11724 = ~new_n10286 & ~new_n11723 ;
  assign new_n11725 = ~new_n11706 & new_n11724 ;
  assign new_n11726 = new_n9283 & ~new_n11725 ;
  assign new_n11727 = ~new_n9283 & new_n11725 ;
  assign new_n11728 = ~new_n11726 & ~new_n11727 ;
  assign new_n11729 = new_n9182 & ~new_n11728 ;
  assign new_n11730 = ~new_n9182 & new_n11726 ;
  assign new_n11731 = ~new_n11729 & ~new_n11730 ;
  assign new_n11732 = ~new_n10260 & ~new_n11731 ;
  assign new_n11733 = ~new_n10260 & new_n11725 ;
  assign new_n11734 = new_n10260 & ~new_n11725 ;
  assign new_n11735 = ~new_n11733 & ~new_n11734 ;
  assign new_n11736 = ~new_n9182 & ~new_n11735 ;
  assign new_n11737 = new_n9182 & new_n11734 ;
  assign new_n11738 = ~new_n11736 & ~new_n11737 ;
  assign new_n11739 = ~new_n11732 & new_n11738 ;
  assign new_n11740 = new_n10232 & ~new_n11739 ;
  assign new_n11741 = ~new_n11691 & ~new_n11740 ;
  assign new_n11742 = ~new_n9804 & ~new_n10232 ;
  assign new_n11743 = ~new_n6720 & new_n10267 ;
  assign new_n11744 = ~new_n9035 & ~new_n10271 ;
  assign new_n11745 = new_n9035 & new_n10269 ;
  assign new_n11746 = ~new_n11744 & ~new_n11745 ;
  assign new_n11747 = ~new_n11743 & new_n11746 ;
  assign new_n11748 = ~new_n10263 & ~new_n11747 ;
  assign new_n11749 = new_n10263 & new_n11747 ;
  assign new_n11750 = ~new_n11748 & ~new_n11749 ;
  assign new_n11751 = ~new_n8939 & ~new_n11750 ;
  assign new_n11752 = new_n8939 & new_n11748 ;
  assign new_n11753 = new_n6667 & new_n10263 ;
  assign new_n11754 = ~new_n11747 & new_n11753 ;
  assign new_n11755 = ~new_n11752 & ~new_n11754 ;
  assign new_n11756 = ~new_n11751 & new_n11755 ;
  assign new_n11757 = new_n10261 & ~new_n11756 ;
  assign new_n11758 = ~new_n6812 & new_n10241 ;
  assign new_n11759 = ~new_n8035 & new_n11269 ;
  assign new_n11760 = ~new_n10240 & ~new_n11759 ;
  assign new_n11761 = ~new_n11758 & new_n11760 ;
  assign new_n11762 = ~new_n8939 & ~new_n9035 ;
  assign new_n11763 = new_n8939 & new_n9035 ;
  assign new_n11764 = ~new_n11762 & ~new_n11763 ;
  assign new_n11765 = ~new_n10234 & ~new_n11764 ;
  assign new_n11766 = ~new_n8939 & new_n9035 ;
  assign new_n11767 = new_n8939 & ~new_n9035 ;
  assign new_n11768 = ~new_n11766 & ~new_n11767 ;
  assign new_n11769 = ~new_n11765 & new_n11768 ;
  assign new_n11770 = ~new_n11761 & ~new_n11769 ;
  assign new_n11771 = new_n10234 & new_n11761 ;
  assign new_n11772 = new_n11762 & new_n11771 ;
  assign new_n11773 = ~new_n11770 & ~new_n11772 ;
  assign new_n11774 = new_n11556 & ~new_n11773 ;
  assign new_n11775 = ~new_n10286 & ~new_n11774 ;
  assign new_n11776 = ~new_n11757 & new_n11775 ;
  assign new_n11777 = new_n9035 & ~new_n11776 ;
  assign new_n11778 = ~new_n9035 & new_n11776 ;
  assign new_n11779 = ~new_n11777 & ~new_n11778 ;
  assign new_n11780 = new_n8939 & ~new_n11779 ;
  assign new_n11781 = ~new_n8939 & new_n11777 ;
  assign new_n11782 = ~new_n11780 & ~new_n11781 ;
  assign new_n11783 = ~new_n10260 & ~new_n11782 ;
  assign new_n11784 = ~new_n10260 & new_n11776 ;
  assign new_n11785 = new_n10260 & ~new_n11776 ;
  assign new_n11786 = ~new_n11784 & ~new_n11785 ;
  assign new_n11787 = ~new_n8939 & ~new_n11786 ;
  assign new_n11788 = new_n8939 & new_n11785 ;
  assign new_n11789 = ~new_n11787 & ~new_n11788 ;
  assign new_n11790 = ~new_n11783 & new_n11789 ;
  assign new_n11791 = new_n10232 & ~new_n11790 ;
  assign new_n11792 = ~new_n11742 & ~new_n11791 ;
  assign new_n11793 = ~new_n9797 & ~new_n10232 ;
  assign new_n11794 = ~new_n8915 & new_n10237 ;
  assign new_n11795 = ~new_n8818 & new_n11794 ;
  assign new_n11796 = ~new_n6582 & new_n10241 ;
  assign new_n11797 = ~new_n10240 & ~new_n11796 ;
  assign new_n11798 = ~new_n11795 & new_n11797 ;
  assign new_n11799 = new_n10236 & ~new_n11798 ;
  assign new_n11800 = ~new_n10236 & new_n11798 ;
  assign new_n11801 = ~new_n11799 & ~new_n11800 ;
  assign new_n11802 = ~new_n7894 & ~new_n11801 ;
  assign new_n11803 = new_n7894 & new_n11799 ;
  assign new_n11804 = ~new_n8818 & new_n8915 ;
  assign new_n11805 = new_n8818 & ~new_n8915 ;
  assign new_n11806 = ~new_n11804 & ~new_n11805 ;
  assign new_n11807 = ~new_n10236 & ~new_n11806 ;
  assign new_n11808 = ~new_n11798 & new_n11807 ;
  assign new_n11809 = ~new_n11803 & ~new_n11808 ;
  assign new_n11810 = ~new_n11802 & new_n11809 ;
  assign new_n11811 = ~new_n6490 & new_n10267 ;
  assign new_n11812 = ~new_n8915 & ~new_n10271 ;
  assign new_n11813 = new_n8915 & new_n10269 ;
  assign new_n11814 = ~new_n11812 & ~new_n11813 ;
  assign new_n11815 = ~new_n11811 & new_n11814 ;
  assign new_n11816 = ~new_n10263 & ~new_n11815 ;
  assign new_n11817 = new_n10263 & new_n11815 ;
  assign new_n11818 = ~new_n11816 & ~new_n11817 ;
  assign new_n11819 = ~new_n8818 & ~new_n11818 ;
  assign new_n11820 = new_n8818 & new_n11816 ;
  assign new_n11821 = new_n6433 & new_n10263 ;
  assign new_n11822 = ~new_n11815 & new_n11821 ;
  assign new_n11823 = ~new_n11820 & ~new_n11822 ;
  assign new_n11824 = ~new_n11819 & new_n11823 ;
  assign new_n11825 = new_n10261 & ~new_n11824 ;
  assign new_n11826 = new_n8818 & new_n8915 ;
  assign new_n11827 = new_n10287 & ~new_n11826 ;
  assign new_n11828 = ~new_n10286 & ~new_n11827 ;
  assign new_n11829 = ~new_n11825 & new_n11828 ;
  assign new_n11830 = ~new_n10258 & ~new_n11829 ;
  assign new_n11831 = new_n10258 & new_n11829 ;
  assign new_n11832 = ~new_n11830 & ~new_n11831 ;
  assign new_n11833 = ~new_n11810 & ~new_n11832 ;
  assign new_n11834 = new_n11810 & new_n11830 ;
  assign new_n11835 = new_n8915 & new_n10258 ;
  assign new_n11836 = ~new_n11829 & new_n11835 ;
  assign new_n11837 = ~new_n11834 & ~new_n11836 ;
  assign new_n11838 = ~new_n11833 & new_n11837 ;
  assign new_n11839 = new_n10232 & ~new_n11838 ;
  assign new_n11840 = ~new_n11793 & ~new_n11839 ;
  assign new_n11841 = lo0200 & new_n3115 ;
  assign new_n11842 = lo0847 & new_n10323 ;
  assign new_n11843 = ~new_n11841 & new_n11842 ;
  assign new_n11844 = new_n11840 & new_n11843 ;
  assign new_n11845 = ~new_n9811 & ~new_n10232 ;
  assign new_n11846 = ~new_n9159 & new_n10237 ;
  assign new_n11847 = ~new_n9059 & new_n11846 ;
  assign new_n11848 = ~new_n7037 & new_n10241 ;
  assign new_n11849 = ~new_n10240 & ~new_n11848 ;
  assign new_n11850 = ~new_n11847 & new_n11849 ;
  assign new_n11851 = new_n10236 & ~new_n11850 ;
  assign new_n11852 = ~new_n10236 & new_n11850 ;
  assign new_n11853 = ~new_n11851 & ~new_n11852 ;
  assign new_n11854 = ~new_n8163 & ~new_n11853 ;
  assign new_n11855 = new_n8163 & new_n11851 ;
  assign new_n11856 = ~new_n9059 & new_n9159 ;
  assign new_n11857 = new_n9059 & ~new_n9159 ;
  assign new_n11858 = ~new_n11856 & ~new_n11857 ;
  assign new_n11859 = ~new_n10236 & ~new_n11858 ;
  assign new_n11860 = ~new_n11850 & new_n11859 ;
  assign new_n11861 = ~new_n11855 & ~new_n11860 ;
  assign new_n11862 = ~new_n11854 & new_n11861 ;
  assign new_n11863 = ~new_n6945 & new_n10267 ;
  assign new_n11864 = ~new_n9159 & ~new_n10271 ;
  assign new_n11865 = new_n9159 & new_n10269 ;
  assign new_n11866 = ~new_n11864 & ~new_n11865 ;
  assign new_n11867 = ~new_n11863 & new_n11866 ;
  assign new_n11868 = ~new_n10263 & ~new_n11867 ;
  assign new_n11869 = new_n10263 & new_n11867 ;
  assign new_n11870 = ~new_n11868 & ~new_n11869 ;
  assign new_n11871 = ~new_n9059 & ~new_n11870 ;
  assign new_n11872 = new_n9059 & new_n11868 ;
  assign new_n11873 = new_n6899 & new_n10263 ;
  assign new_n11874 = ~new_n11867 & new_n11873 ;
  assign new_n11875 = ~new_n11872 & ~new_n11874 ;
  assign new_n11876 = ~new_n11871 & new_n11875 ;
  assign new_n11877 = new_n10261 & ~new_n11876 ;
  assign new_n11878 = new_n9059 & new_n9159 ;
  assign new_n11879 = new_n10287 & ~new_n11878 ;
  assign new_n11880 = ~new_n10286 & ~new_n11879 ;
  assign new_n11881 = ~new_n11877 & new_n11880 ;
  assign new_n11882 = ~new_n10258 & ~new_n11881 ;
  assign new_n11883 = new_n10258 & new_n11881 ;
  assign new_n11884 = ~new_n11882 & ~new_n11883 ;
  assign new_n11885 = ~new_n11862 & ~new_n11884 ;
  assign new_n11886 = new_n11862 & new_n11882 ;
  assign new_n11887 = new_n9159 & new_n10258 ;
  assign new_n11888 = ~new_n11881 & new_n11887 ;
  assign new_n11889 = ~new_n11886 & ~new_n11888 ;
  assign new_n11890 = ~new_n11885 & new_n11889 ;
  assign new_n11891 = new_n10232 & ~new_n11890 ;
  assign new_n11892 = ~new_n11845 & ~new_n11891 ;
  assign new_n11893 = new_n10302 & new_n11892 ;
  assign new_n11894 = new_n11844 & new_n11893 ;
  assign new_n11895 = new_n11792 & new_n11894 ;
  assign new_n11896 = new_n11741 & new_n11895 ;
  assign new_n11897 = new_n11690 & new_n11896 ;
  assign new_n11898 = new_n11639 & new_n11897 ;
  assign new_n11899 = new_n11591 & new_n11898 ;
  assign new_n11900 = new_n11539 & new_n11899 ;
  assign new_n11901 = new_n11490 & new_n11900 ;
  assign new_n11902 = new_n11443 & new_n11901 ;
  assign new_n11903 = new_n11394 & new_n11902 ;
  assign new_n11904 = new_n11347 & new_n11903 ;
  assign new_n11905 = new_n11298 & new_n11904 ;
  assign new_n11906 = new_n11250 & new_n11905 ;
  assign new_n11907 = new_n11181 & new_n11906 ;
  assign new_n11908 = new_n11136 & new_n11907 ;
  assign new_n11909 = new_n11082 & new_n11908 ;
  assign new_n11910 = new_n11035 & new_n11909 ;
  assign new_n11911 = new_n10990 & new_n11910 ;
  assign new_n11912 = new_n10943 & new_n11911 ;
  assign new_n11913 = new_n10898 & new_n11912 ;
  assign new_n11914 = new_n10851 & new_n11913 ;
  assign new_n11915 = new_n10806 & new_n11914 ;
  assign new_n11916 = new_n10759 & new_n11915 ;
  assign new_n11917 = new_n10714 & new_n11916 ;
  assign new_n11918 = new_n10667 & new_n11917 ;
  assign new_n11919 = new_n10622 & new_n11918 ;
  assign new_n11920 = new_n10575 & new_n11919 ;
  assign new_n11921 = new_n10529 & new_n11920 ;
  assign new_n11922 = new_n10482 & new_n11921 ;
  assign new_n11923 = new_n10432 & new_n11922 ;
  assign new_n11924 = new_n5766 & new_n6690 ;
  assign new_n11925 = new_n4541 & new_n11924 ;
  assign new_n11926 = new_n2910 & new_n5996 ;
  assign new_n11927 = new_n3549 & new_n6917 ;
  assign new_n11928 = new_n11926 & new_n11927 ;
  assign new_n11929 = new_n4992 & new_n6461 ;
  assign new_n11930 = new_n3464 & new_n4630 ;
  assign new_n11931 = new_n11929 & new_n11930 ;
  assign new_n11932 = new_n11928 & new_n11931 ;
  assign new_n11933 = new_n11925 & new_n11932 ;
  assign new_n11934 = new_n11841 & new_n11842 ;
  assign new_n11935 = new_n5187 & new_n11934 ;
  assign new_n11936 = new_n5276 & new_n5472 ;
  assign new_n11937 = new_n2619 & new_n4818 ;
  assign new_n11938 = new_n11936 & new_n11937 ;
  assign new_n11939 = new_n11935 & new_n11938 ;
  assign new_n11940 = new_n2824 & new_n3734 ;
  assign new_n11941 = new_n4461 & new_n4904 ;
  assign new_n11942 = new_n11940 & new_n11941 ;
  assign new_n11943 = new_n4097 & new_n7138 ;
  assign new_n11944 = new_n3817 & new_n5560 ;
  assign new_n11945 = new_n11943 & new_n11944 ;
  assign new_n11946 = new_n11942 & new_n11945 ;
  assign new_n11947 = new_n3383 & new_n4268 ;
  assign new_n11948 = new_n3908 & new_n4179 ;
  assign new_n11949 = new_n11947 & new_n11948 ;
  assign new_n11950 = new_n3092 & new_n6225 ;
  assign new_n11951 = new_n2739 & new_n3001 ;
  assign new_n11952 = new_n11950 & new_n11951 ;
  assign new_n11953 = new_n11949 & new_n11952 ;
  assign new_n11954 = new_n11946 & new_n11953 ;
  assign new_n11955 = new_n11939 & new_n11954 ;
  assign new_n11956 = new_n11933 & new_n11955 ;
  assign new_n11957 = ~new_n4097 & new_n5086 ;
  assign new_n11958 = new_n4097 & ~new_n5086 ;
  assign new_n11959 = ~new_n11957 & ~new_n11958 ;
  assign new_n11960 = ~new_n3092 & new_n3639 ;
  assign new_n11961 = new_n3092 & ~new_n3639 ;
  assign new_n11962 = ~new_n11960 & ~new_n11961 ;
  assign new_n11963 = ~new_n4541 & new_n5370 ;
  assign new_n11964 = new_n4541 & ~new_n5370 ;
  assign new_n11965 = ~new_n11963 & ~new_n11964 ;
  assign new_n11966 = new_n11962 & new_n11965 ;
  assign new_n11967 = new_n11959 & new_n11966 ;
  assign new_n11968 = ~new_n3817 & new_n4724 ;
  assign new_n11969 = new_n3817 & ~new_n4724 ;
  assign new_n11970 = ~new_n11968 & ~new_n11969 ;
  assign new_n11971 = new_n3464 & ~new_n4362 ;
  assign new_n11972 = new_n4818 & ~new_n5654 ;
  assign new_n11973 = ~new_n11971 & ~new_n11972 ;
  assign new_n11974 = new_n11970 & new_n11973 ;
  assign new_n11975 = ~new_n3464 & new_n4362 ;
  assign new_n11976 = ~new_n4818 & new_n5654 ;
  assign new_n11977 = ~new_n11975 & ~new_n11976 ;
  assign new_n11978 = ~new_n3001 & new_n4003 ;
  assign new_n11979 = new_n3001 & ~new_n4003 ;
  assign new_n11980 = ~new_n11978 & ~new_n11979 ;
  assign new_n11981 = new_n11977 & new_n11980 ;
  assign new_n11982 = new_n11974 & new_n11981 ;
  assign new_n11983 = new_n11967 & new_n11982 ;
  assign new_n11984 = ~new_n6461 & new_n8902 ;
  assign new_n11985 = new_n6461 & ~new_n8902 ;
  assign new_n11986 = ~new_n11984 & ~new_n11985 ;
  assign new_n11987 = ~new_n6225 & new_n8780 ;
  assign new_n11988 = new_n6690 & ~new_n9021 ;
  assign new_n11989 = ~new_n11987 & ~new_n11988 ;
  assign new_n11990 = new_n11986 & new_n11989 ;
  assign new_n11991 = ~new_n6917 & new_n9141 ;
  assign new_n11992 = new_n6917 & ~new_n9141 ;
  assign new_n11993 = ~new_n11991 & ~new_n11992 ;
  assign new_n11994 = ~new_n5996 & new_n8659 ;
  assign new_n11995 = new_n5996 & ~new_n8659 ;
  assign new_n11996 = ~new_n11994 & ~new_n11995 ;
  assign new_n11997 = new_n11993 & new_n11996 ;
  assign new_n11998 = new_n11990 & new_n11997 ;
  assign new_n11999 = ~new_n7138 & new_n9266 ;
  assign new_n12000 = new_n7138 & ~new_n9266 ;
  assign new_n12001 = ~new_n11999 & ~new_n12000 ;
  assign new_n12002 = new_n6225 & ~new_n8780 ;
  assign new_n12003 = ~new_n6690 & new_n9021 ;
  assign new_n12004 = ~new_n12002 & ~new_n12003 ;
  assign new_n12005 = new_n12001 & new_n12004 ;
  assign new_n12006 = new_n2619 & ~new_n9389 ;
  assign new_n12007 = ~new_n2619 & new_n9389 ;
  assign new_n12008 = ~new_n12006 & ~new_n12007 ;
  assign new_n12009 = ~new_n5766 & new_n8533 ;
  assign new_n12010 = new_n5766 & ~new_n8533 ;
  assign new_n12011 = ~new_n12009 & ~new_n12010 ;
  assign new_n12012 = new_n12008 & new_n12011 ;
  assign new_n12013 = new_n12005 & new_n12012 ;
  assign new_n12014 = new_n11998 & new_n12013 ;
  assign new_n12015 = new_n11983 & new_n12014 ;
  assign new_n12016 = ~new_n4179 & new_n7883 ;
  assign new_n12017 = new_n4179 & ~new_n7883 ;
  assign new_n12018 = ~new_n12016 & ~new_n12017 ;
  assign new_n12019 = ~new_n5187 & new_n8281 ;
  assign new_n12020 = new_n4461 & ~new_n8008 ;
  assign new_n12021 = ~new_n12019 & ~new_n12020 ;
  assign new_n12022 = new_n12018 & new_n12021 ;
  assign new_n12023 = ~new_n4904 & new_n8149 ;
  assign new_n12024 = new_n4904 & ~new_n8149 ;
  assign new_n12025 = ~new_n12023 & ~new_n12024 ;
  assign new_n12026 = ~new_n3383 & new_n7637 ;
  assign new_n12027 = new_n3383 & ~new_n7637 ;
  assign new_n12028 = ~new_n12026 & ~new_n12027 ;
  assign new_n12029 = new_n12025 & new_n12028 ;
  assign new_n12030 = new_n12022 & new_n12029 ;
  assign new_n12031 = ~new_n2910 & new_n7512 ;
  assign new_n12032 = new_n2910 & ~new_n7512 ;
  assign new_n12033 = ~new_n12031 & ~new_n12032 ;
  assign new_n12034 = new_n5187 & ~new_n8281 ;
  assign new_n12035 = ~new_n4461 & new_n8008 ;
  assign new_n12036 = ~new_n12034 & ~new_n12035 ;
  assign new_n12037 = new_n12033 & new_n12036 ;
  assign new_n12038 = ~new_n3734 & new_n7761 ;
  assign new_n12039 = new_n3734 & ~new_n7761 ;
  assign new_n12040 = ~new_n12038 & ~new_n12039 ;
  assign new_n12041 = ~new_n5472 & new_n8411 ;
  assign new_n12042 = new_n5472 & ~new_n8411 ;
  assign new_n12043 = ~new_n12041 & ~new_n12042 ;
  assign new_n12044 = new_n12040 & new_n12043 ;
  assign new_n12045 = new_n12037 & new_n12044 ;
  assign new_n12046 = new_n12030 & new_n12045 ;
  assign new_n12047 = ~new_n4268 & new_n6571 ;
  assign new_n12048 = new_n4268 & ~new_n6571 ;
  assign new_n12049 = ~new_n12047 & ~new_n12048 ;
  assign new_n12050 = ~new_n5276 & new_n7249 ;
  assign new_n12051 = new_n4630 & ~new_n6801 ;
  assign new_n12052 = ~new_n12050 & ~new_n12051 ;
  assign new_n12053 = new_n12049 & new_n12052 ;
  assign new_n12054 = ~new_n4992 & new_n7026 ;
  assign new_n12055 = new_n4992 & ~new_n7026 ;
  assign new_n12056 = ~new_n12054 & ~new_n12055 ;
  assign new_n12057 = ~new_n3549 & new_n6106 ;
  assign new_n12058 = new_n3549 & ~new_n6106 ;
  assign new_n12059 = ~new_n12057 & ~new_n12058 ;
  assign new_n12060 = new_n12056 & new_n12059 ;
  assign new_n12061 = new_n12053 & new_n12060 ;
  assign new_n12062 = ~new_n2824 & new_n5880 ;
  assign new_n12063 = new_n2824 & ~new_n5880 ;
  assign new_n12064 = ~new_n12062 & ~new_n12063 ;
  assign new_n12065 = new_n5276 & ~new_n7249 ;
  assign new_n12066 = ~new_n4630 & new_n6801 ;
  assign new_n12067 = ~new_n12065 & ~new_n12066 ;
  assign new_n12068 = new_n12064 & new_n12067 ;
  assign new_n12069 = ~new_n3908 & new_n6336 ;
  assign new_n12070 = new_n3908 & ~new_n6336 ;
  assign new_n12071 = ~new_n12069 & ~new_n12070 ;
  assign new_n12072 = ~new_n5560 & new_n7374 ;
  assign new_n12073 = new_n5560 & ~new_n7374 ;
  assign new_n12074 = ~new_n12072 & ~new_n12073 ;
  assign new_n12075 = new_n12071 & new_n12074 ;
  assign new_n12076 = new_n12068 & new_n12075 ;
  assign new_n12077 = new_n12061 & new_n12076 ;
  assign new_n12078 = new_n12046 & new_n12077 ;
  assign new_n12079 = new_n12015 & new_n12078 ;
  assign new_n12080 = new_n10227 & new_n12079 ;
  assign new_n12081 = new_n2739 & ~new_n12080 ;
  assign new_n12082 = new_n7138 & new_n12007 ;
  assign new_n12083 = new_n7138 & ~new_n12082 ;
  assign new_n12084 = new_n9266 & ~new_n12083 ;
  assign new_n12085 = ~new_n7138 & ~new_n9266 ;
  assign new_n12086 = new_n12007 & new_n12085 ;
  assign new_n12087 = ~new_n12084 & ~new_n12086 ;
  assign new_n12088 = new_n6917 & ~new_n12087 ;
  assign new_n12089 = new_n6917 & ~new_n12088 ;
  assign new_n12090 = new_n9141 & ~new_n12089 ;
  assign new_n12091 = ~new_n6917 & ~new_n9141 ;
  assign new_n12092 = ~new_n12087 & new_n12091 ;
  assign new_n12093 = ~new_n12090 & ~new_n12092 ;
  assign new_n12094 = new_n6690 & ~new_n12093 ;
  assign new_n12095 = new_n6690 & ~new_n12094 ;
  assign new_n12096 = new_n9021 & ~new_n12095 ;
  assign new_n12097 = ~new_n6690 & ~new_n9021 ;
  assign new_n12098 = ~new_n12093 & new_n12097 ;
  assign new_n12099 = ~new_n12096 & ~new_n12098 ;
  assign new_n12100 = new_n6461 & ~new_n12099 ;
  assign new_n12101 = new_n6461 & ~new_n12100 ;
  assign new_n12102 = new_n8902 & ~new_n12101 ;
  assign new_n12103 = ~new_n6461 & ~new_n8902 ;
  assign new_n12104 = ~new_n12099 & new_n12103 ;
  assign new_n12105 = ~new_n12102 & ~new_n12104 ;
  assign new_n12106 = new_n6225 & ~new_n12105 ;
  assign new_n12107 = new_n6225 & ~new_n12106 ;
  assign new_n12108 = new_n8780 & ~new_n12107 ;
  assign new_n12109 = ~new_n6225 & ~new_n8780 ;
  assign new_n12110 = ~new_n12105 & new_n12109 ;
  assign new_n12111 = ~new_n12108 & ~new_n12110 ;
  assign new_n12112 = new_n5996 & ~new_n12111 ;
  assign new_n12113 = new_n5996 & ~new_n12112 ;
  assign new_n12114 = new_n8659 & ~new_n12113 ;
  assign new_n12115 = ~new_n5996 & ~new_n8659 ;
  assign new_n12116 = ~new_n12111 & new_n12115 ;
  assign new_n12117 = ~new_n12114 & ~new_n12116 ;
  assign new_n12118 = new_n5766 & ~new_n12117 ;
  assign new_n12119 = new_n5766 & ~new_n12118 ;
  assign new_n12120 = new_n8533 & ~new_n12119 ;
  assign new_n12121 = ~new_n5766 & ~new_n8533 ;
  assign new_n12122 = ~new_n12117 & new_n12121 ;
  assign new_n12123 = ~new_n12120 & ~new_n12122 ;
  assign new_n12124 = new_n5472 & ~new_n12123 ;
  assign new_n12125 = new_n5472 & ~new_n12124 ;
  assign new_n12126 = new_n8411 & ~new_n12125 ;
  assign new_n12127 = ~new_n5472 & ~new_n8411 ;
  assign new_n12128 = ~new_n12123 & new_n12127 ;
  assign new_n12129 = ~new_n12126 & ~new_n12128 ;
  assign new_n12130 = new_n5187 & ~new_n12129 ;
  assign new_n12131 = new_n5187 & ~new_n12130 ;
  assign new_n12132 = new_n8281 & ~new_n12131 ;
  assign new_n12133 = ~new_n5187 & ~new_n8281 ;
  assign new_n12134 = ~new_n12129 & new_n12133 ;
  assign new_n12135 = ~new_n12132 & ~new_n12134 ;
  assign new_n12136 = new_n4904 & ~new_n12135 ;
  assign new_n12137 = new_n4904 & ~new_n12136 ;
  assign new_n12138 = new_n8149 & ~new_n12137 ;
  assign new_n12139 = ~new_n4904 & ~new_n8149 ;
  assign new_n12140 = ~new_n12135 & new_n12139 ;
  assign new_n12141 = ~new_n12138 & ~new_n12140 ;
  assign new_n12142 = new_n4461 & ~new_n12141 ;
  assign new_n12143 = new_n4461 & ~new_n12142 ;
  assign new_n12144 = new_n8008 & ~new_n12143 ;
  assign new_n12145 = ~new_n4461 & ~new_n8008 ;
  assign new_n12146 = ~new_n12141 & new_n12145 ;
  assign new_n12147 = ~new_n12144 & ~new_n12146 ;
  assign new_n12148 = new_n4179 & ~new_n12147 ;
  assign new_n12149 = new_n4179 & ~new_n12148 ;
  assign new_n12150 = new_n7883 & ~new_n12149 ;
  assign new_n12151 = ~new_n4179 & ~new_n7883 ;
  assign new_n12152 = ~new_n12147 & new_n12151 ;
  assign new_n12153 = ~new_n12150 & ~new_n12152 ;
  assign new_n12154 = new_n3734 & ~new_n12153 ;
  assign new_n12155 = new_n3734 & ~new_n12154 ;
  assign new_n12156 = new_n7761 & ~new_n12155 ;
  assign new_n12157 = ~new_n3734 & ~new_n7761 ;
  assign new_n12158 = ~new_n12153 & new_n12157 ;
  assign new_n12159 = ~new_n12156 & ~new_n12158 ;
  assign new_n12160 = new_n3383 & ~new_n12159 ;
  assign new_n12161 = new_n3383 & ~new_n12160 ;
  assign new_n12162 = new_n7637 & ~new_n12161 ;
  assign new_n12163 = ~new_n3383 & ~new_n7637 ;
  assign new_n12164 = ~new_n12159 & new_n12163 ;
  assign new_n12165 = ~new_n12162 & ~new_n12164 ;
  assign new_n12166 = new_n2910 & ~new_n12165 ;
  assign new_n12167 = new_n2910 & ~new_n12166 ;
  assign new_n12168 = new_n7512 & ~new_n12167 ;
  assign new_n12169 = ~new_n2910 & ~new_n7512 ;
  assign new_n12170 = ~new_n12165 & new_n12169 ;
  assign new_n12171 = ~new_n12168 & ~new_n12170 ;
  assign new_n12172 = new_n5560 & ~new_n12171 ;
  assign new_n12173 = new_n5560 & ~new_n12172 ;
  assign new_n12174 = new_n7374 & ~new_n12173 ;
  assign new_n12175 = ~new_n5560 & ~new_n7374 ;
  assign new_n12176 = ~new_n12171 & new_n12175 ;
  assign new_n12177 = ~new_n12174 & ~new_n12176 ;
  assign new_n12178 = new_n5276 & ~new_n12177 ;
  assign new_n12179 = new_n5276 & ~new_n12178 ;
  assign new_n12180 = new_n7249 & ~new_n12179 ;
  assign new_n12181 = ~new_n5276 & ~new_n7249 ;
  assign new_n12182 = ~new_n12177 & new_n12181 ;
  assign new_n12183 = ~new_n12180 & ~new_n12182 ;
  assign new_n12184 = new_n4992 & ~new_n12183 ;
  assign new_n12185 = new_n4992 & ~new_n12184 ;
  assign new_n12186 = new_n7026 & ~new_n12185 ;
  assign new_n12187 = ~new_n4992 & ~new_n7026 ;
  assign new_n12188 = ~new_n12183 & new_n12187 ;
  assign new_n12189 = ~new_n12186 & ~new_n12188 ;
  assign new_n12190 = new_n4630 & ~new_n12189 ;
  assign new_n12191 = new_n4630 & ~new_n12190 ;
  assign new_n12192 = new_n6801 & ~new_n12191 ;
  assign new_n12193 = ~new_n4630 & ~new_n6801 ;
  assign new_n12194 = ~new_n12189 & new_n12193 ;
  assign new_n12195 = ~new_n12192 & ~new_n12194 ;
  assign new_n12196 = new_n4268 & ~new_n12195 ;
  assign new_n12197 = new_n4268 & ~new_n12196 ;
  assign new_n12198 = new_n6571 & ~new_n12197 ;
  assign new_n12199 = ~new_n4268 & ~new_n6571 ;
  assign new_n12200 = ~new_n12195 & new_n12199 ;
  assign new_n12201 = ~new_n12198 & ~new_n12200 ;
  assign new_n12202 = new_n3908 & ~new_n12201 ;
  assign new_n12203 = new_n3908 & ~new_n12202 ;
  assign new_n12204 = new_n6336 & ~new_n12203 ;
  assign new_n12205 = ~new_n3908 & ~new_n6336 ;
  assign new_n12206 = ~new_n12201 & new_n12205 ;
  assign new_n12207 = ~new_n12204 & ~new_n12206 ;
  assign new_n12208 = new_n3549 & ~new_n12207 ;
  assign new_n12209 = new_n3549 & ~new_n12208 ;
  assign new_n12210 = new_n6106 & ~new_n12209 ;
  assign new_n12211 = ~new_n3549 & ~new_n6106 ;
  assign new_n12212 = ~new_n12207 & new_n12211 ;
  assign new_n12213 = ~new_n12210 & ~new_n12212 ;
  assign new_n12214 = new_n2824 & ~new_n12213 ;
  assign new_n12215 = new_n2824 & ~new_n12214 ;
  assign new_n12216 = new_n5880 & ~new_n12215 ;
  assign new_n12217 = ~new_n2824 & ~new_n5880 ;
  assign new_n12218 = ~new_n12213 & new_n12217 ;
  assign new_n12219 = ~new_n12216 & ~new_n12218 ;
  assign new_n12220 = new_n4818 & ~new_n12219 ;
  assign new_n12221 = new_n4818 & ~new_n12220 ;
  assign new_n12222 = new_n5654 & ~new_n12221 ;
  assign new_n12223 = ~new_n4818 & ~new_n5654 ;
  assign new_n12224 = ~new_n12219 & new_n12223 ;
  assign new_n12225 = ~new_n12222 & ~new_n12224 ;
  assign new_n12226 = new_n4541 & ~new_n12225 ;
  assign new_n12227 = new_n4541 & ~new_n12226 ;
  assign new_n12228 = new_n5370 & ~new_n12227 ;
  assign new_n12229 = ~new_n4541 & ~new_n5370 ;
  assign new_n12230 = ~new_n12225 & new_n12229 ;
  assign new_n12231 = ~new_n12228 & ~new_n12230 ;
  assign new_n12232 = new_n4097 & ~new_n12231 ;
  assign new_n12233 = new_n4097 & ~new_n12232 ;
  assign new_n12234 = new_n5086 & ~new_n12233 ;
  assign new_n12235 = ~new_n4097 & ~new_n5086 ;
  assign new_n12236 = ~new_n12231 & new_n12235 ;
  assign new_n12237 = ~new_n12234 & ~new_n12236 ;
  assign new_n12238 = new_n3817 & ~new_n12237 ;
  assign new_n12239 = new_n3817 & ~new_n12238 ;
  assign new_n12240 = new_n4724 & ~new_n12239 ;
  assign new_n12241 = ~new_n3817 & ~new_n4724 ;
  assign new_n12242 = ~new_n12237 & new_n12241 ;
  assign new_n12243 = ~new_n12240 & ~new_n12242 ;
  assign new_n12244 = new_n3464 & ~new_n12243 ;
  assign new_n12245 = new_n3464 & ~new_n12244 ;
  assign new_n12246 = new_n4362 & ~new_n12245 ;
  assign new_n12247 = ~new_n3464 & ~new_n4362 ;
  assign new_n12248 = ~new_n12243 & new_n12247 ;
  assign new_n12249 = ~new_n12246 & ~new_n12248 ;
  assign new_n12250 = new_n3001 & ~new_n12249 ;
  assign new_n12251 = new_n3001 & ~new_n12250 ;
  assign new_n12252 = new_n4003 & ~new_n12251 ;
  assign new_n12253 = ~new_n3001 & ~new_n4003 ;
  assign new_n12254 = ~new_n12249 & new_n12253 ;
  assign new_n12255 = ~new_n12252 & ~new_n12254 ;
  assign new_n12256 = new_n3092 & ~new_n12255 ;
  assign new_n12257 = new_n3092 & ~new_n12256 ;
  assign new_n12258 = new_n3639 & ~new_n12257 ;
  assign new_n12259 = ~new_n3092 & ~new_n3639 ;
  assign new_n12260 = ~new_n12255 & new_n12259 ;
  assign new_n12261 = ~new_n12258 & ~new_n12260 ;
  assign new_n12262 = new_n10227 & ~new_n12261 ;
  assign new_n12263 = ~new_n10225 & ~new_n12262 ;
  assign new_n12264 = ~lo0851 & lo0852 ;
  assign new_n12265 = ~new_n12263 & new_n12264 ;
  assign new_n12266 = lo0851 & lo0852 ;
  assign new_n12267 = new_n10227 & new_n11983 ;
  assign new_n12268 = ~new_n12046 & ~new_n12077 ;
  assign new_n12269 = ~new_n12014 & new_n12268 ;
  assign new_n12270 = ~new_n12267 & new_n12269 ;
  assign new_n12271 = ~lo0851 & ~lo0852 ;
  assign new_n12272 = ~new_n12270 & new_n12271 ;
  assign new_n12273 = ~new_n12266 & ~new_n12272 ;
  assign new_n12274 = ~new_n12265 & new_n12273 ;
  assign new_n12275 = ~lo0851 & ~new_n12274 ;
  assign new_n12276 = lo0851 & new_n12274 ;
  assign new_n12277 = ~new_n12275 & ~new_n12276 ;
  assign new_n12278 = new_n12081 & ~new_n12277 ;
  assign new_n12279 = ~new_n12081 & new_n12275 ;
  assign new_n12280 = ~new_n10226 & ~new_n12262 ;
  assign new_n12281 = lo0851 & ~new_n12280 ;
  assign new_n12282 = ~new_n12274 & new_n12281 ;
  assign new_n12283 = ~new_n12279 & ~new_n12282 ;
  assign new_n12284 = ~new_n12278 & new_n12283 ;
  assign new_n12285 = lo0850 & ~new_n12284 ;
  assign new_n12286 = ~new_n12079 & new_n12261 ;
  assign new_n12287 = new_n10227 & ~new_n12286 ;
  assign new_n12288 = ~new_n10225 & ~new_n12287 ;
  assign new_n12289 = lo0852 & ~new_n12080 ;
  assign new_n12290 = ~new_n12080 & ~new_n12289 ;
  assign new_n12291 = lo0851 & ~new_n12290 ;
  assign new_n12292 = new_n12080 & new_n12271 ;
  assign new_n12293 = lo0851 & ~lo0852 ;
  assign new_n12294 = new_n12081 & new_n12293 ;
  assign new_n12295 = ~new_n12292 & ~new_n12294 ;
  assign new_n12296 = ~new_n12291 & new_n12295 ;
  assign new_n12297 = ~lo0852 & ~new_n12296 ;
  assign new_n12298 = new_n12288 & new_n12297 ;
  assign new_n12299 = lo0852 & new_n12296 ;
  assign new_n12300 = ~new_n12297 & ~new_n12299 ;
  assign new_n12301 = ~new_n12288 & ~new_n12300 ;
  assign new_n12302 = ~new_n10226 & ~new_n12287 ;
  assign new_n12303 = lo0852 & ~new_n12296 ;
  assign new_n12304 = ~new_n12302 & new_n12303 ;
  assign new_n12305 = ~new_n12301 & ~new_n12304 ;
  assign new_n12306 = ~new_n12298 & new_n12305 ;
  assign new_n12307 = ~lo0850 & ~new_n12306 ;
  assign new_n12308 = ~new_n12285 & ~new_n12307 ;
  assign new_n12309 = lo0849 & ~new_n12308 ;
  assign new_n12310 = ~new_n11956 & ~new_n12309 ;
  assign new_n12311 = ~new_n11923 & new_n12310 ;
  assign new_n12312 = ~new_n10354 & new_n12311 ;
  assign new_n12313 = ~new_n10325 & new_n12312 ;
  assign new_n12314 = ~new_n2465 & new_n12313 ;
  assign new_n12315 = new_n2465 & ~new_n12313 ;
  assign new_n12316 = ~new_n12314 & ~new_n12315 ;
  assign new_n12317 = ~lo1292 & ~new_n12316 ;
  assign new_n12318 = new_n2456 & ~new_n12317 ;
  assign new_n12319 = ~new_n2412 & new_n2442 ;
  assign new_n12320 = new_n2298 & ~new_n2402 ;
  assign new_n12321 = ~new_n2442 & ~new_n12320 ;
  assign new_n12322 = ~new_n12319 & ~new_n12321 ;
  assign new_n12323 = new_n2265 & ~new_n12322 ;
  assign new_n12324 = lo0193 & ~new_n2265 ;
  assign new_n12325 = ~new_n12323 & ~new_n12324 ;
  assign new_n12326 = lo0191 & ~new_n2265 ;
  assign new_n12327 = new_n2285 & new_n2443 ;
  assign new_n12328 = new_n2265 & ~new_n12327 ;
  assign new_n12329 = ~new_n12326 & ~new_n12328 ;
  assign new_n12330 = lo1291 & lo1292 ;
  assign new_n12331 = new_n2262 & new_n12330 ;
  assign new_n12332 = ~lo1293 & lo1294 ;
  assign new_n12333 = ~lo1293 & ~new_n12332 ;
  assign new_n12334 = ~new_n12331 & new_n12333 ;
  assign new_n12335 = new_n12325 & new_n12334 ;
  assign new_n12336 = new_n12329 & new_n12335 ;
  assign new_n12337 = ~new_n12325 & ~new_n12329 ;
  assign new_n12338 = lo1291 & ~lo1292 ;
  assign new_n12339 = ~lo1291 & lo1292 ;
  assign new_n12340 = ~new_n12338 & ~new_n12339 ;
  assign new_n12341 = ~lo1294 & ~new_n12340 ;
  assign new_n12342 = lo1293 & new_n12341 ;
  assign new_n12343 = new_n12325 & new_n12342 ;
  assign new_n12344 = ~new_n12329 & new_n12343 ;
  assign new_n12345 = ~new_n12337 & ~new_n12344 ;
  assign new_n12346 = ~new_n12336 & new_n12345 ;
  assign new_n12347 = new_n12325 & ~new_n12346 ;
  assign new_n12348 = ~new_n12325 & new_n12346 ;
  assign new_n12349 = ~new_n12347 & ~new_n12348 ;
  assign new_n12350 = new_n12318 & ~new_n12349 ;
  assign new_n12351 = ~new_n12318 & new_n12347 ;
  assign new_n12352 = lo0192 & ~new_n2265 ;
  assign new_n12353 = lo0129 & ~new_n2395 ;
  assign new_n12354 = new_n2292 & ~new_n12353 ;
  assign new_n12355 = ~new_n2442 & ~new_n12354 ;
  assign new_n12356 = new_n2265 & new_n12355 ;
  assign new_n12357 = ~new_n12352 & ~new_n12356 ;
  assign new_n12358 = new_n12325 & new_n12357 ;
  assign new_n12359 = new_n2408 & new_n2442 ;
  assign new_n12360 = ~new_n2317 & ~new_n2402 ;
  assign new_n12361 = ~lo0129 & new_n2402 ;
  assign new_n12362 = ~new_n12360 & ~new_n12361 ;
  assign new_n12363 = ~new_n2442 & ~new_n12362 ;
  assign new_n12364 = ~new_n12359 & ~new_n12363 ;
  assign new_n12365 = new_n2265 & ~new_n12364 ;
  assign new_n12366 = lo0195 & ~new_n2265 ;
  assign new_n12367 = ~new_n12365 & ~new_n12366 ;
  assign new_n12368 = ~new_n2465 & ~new_n12367 ;
  assign new_n12369 = new_n12358 & new_n12368 ;
  assign new_n12370 = ~new_n12325 & ~new_n12357 ;
  assign new_n12371 = ~new_n12369 & ~new_n12370 ;
  assign new_n12372 = ~new_n12329 & ~new_n12371 ;
  assign new_n12373 = ~new_n12357 & ~new_n12367 ;
  assign new_n12374 = new_n12329 & new_n12373 ;
  assign new_n12375 = ~new_n12372 & ~new_n12374 ;
  assign new_n12376 = lo1291 & new_n2263 ;
  assign new_n12377 = ~new_n12325 & new_n12376 ;
  assign new_n12378 = ~new_n12346 & new_n12377 ;
  assign new_n12379 = ~new_n12375 & ~new_n12378 ;
  assign new_n12380 = ~new_n12351 & new_n12379 ;
  assign new_n12381 = ~new_n12350 & new_n12380 ;
  assign new_n12382 = new_n2455 & ~new_n12381 ;
  assign new_n12383 = lo1292 & new_n2456 ;
  assign new_n12384 = new_n12329 & new_n12383 ;
  assign new_n12385 = new_n2465 & ~new_n12325 ;
  assign new_n12386 = new_n12357 & ~new_n12385 ;
  assign new_n12387 = lo1293 & ~lo1294 ;
  assign new_n12388 = lo1291 & new_n12387 ;
  assign new_n12389 = ~new_n12386 & new_n12388 ;
  assign new_n12390 = new_n12330 & new_n12387 ;
  assign new_n12391 = ~lo1291 & ~lo1292 ;
  assign new_n12392 = new_n12332 & new_n12391 ;
  assign new_n12393 = ~new_n12390 & ~new_n12392 ;
  assign new_n12394 = new_n12325 & ~new_n12393 ;
  assign new_n12395 = ~new_n2465 & ~new_n12325 ;
  assign new_n12396 = new_n12342 & new_n12395 ;
  assign new_n12397 = ~new_n12394 & ~new_n12396 ;
  assign new_n12398 = new_n12357 & ~new_n12397 ;
  assign new_n12399 = ~new_n12389 & ~new_n12398 ;
  assign new_n12400 = ~new_n12329 & ~new_n12399 ;
  assign new_n12401 = ~new_n12384 & ~new_n12400 ;
  assign new_n12402 = ~new_n2450 & ~new_n2454 ;
  assign new_n12403 = ~new_n12401 & new_n12402 ;
  assign new_n12404 = new_n2450 & ~new_n2454 ;
  assign new_n12405 = ~new_n2450 & new_n2454 ;
  assign new_n12406 = new_n12329 & ~new_n12383 ;
  assign new_n12407 = new_n12405 & ~new_n12406 ;
  assign new_n12408 = ~new_n12404 & ~new_n12407 ;
  assign new_n12409 = ~new_n12403 & new_n12408 ;
  assign new_n12410 = ~new_n12382 & new_n12409 ;
  assign new_n12411 = ~new_n2446 & ~new_n12410 ;
  assign new_n12412 = ~new_n2279 & new_n2443 ;
  assign new_n12413 = ~lo0176 & ~new_n2414 ;
  assign new_n12414 = lo0860 & new_n2414 ;
  assign new_n12415 = ~new_n12413 & ~new_n12414 ;
  assign new_n12416 = new_n2442 & ~new_n12415 ;
  assign new_n12417 = ~new_n12412 & ~new_n12416 ;
  assign new_n12418 = new_n2265 & ~new_n12417 ;
  assign new_n12419 = lo0861 & ~new_n2265 ;
  assign new_n12420 = ~new_n12418 & ~new_n12419 ;
  assign new_n12421 = ~new_n2362 & new_n2443 ;
  assign new_n12422 = ~lo0175 & ~lo0862 ;
  assign new_n12423 = ~lo0180 & new_n12422 ;
  assign new_n12424 = new_n2403 & ~new_n12423 ;
  assign new_n12425 = new_n2442 & new_n12424 ;
  assign new_n12426 = ~new_n12421 & ~new_n12425 ;
  assign new_n12427 = new_n2265 & ~new_n12426 ;
  assign new_n12428 = lo0863 & ~new_n2265 ;
  assign new_n12429 = ~new_n12427 & ~new_n12428 ;
  assign new_n12430 = ~lo0180 & ~lo0864 ;
  assign new_n12431 = ~lo0175 & ~new_n12430 ;
  assign new_n12432 = new_n2403 & ~new_n12431 ;
  assign new_n12433 = new_n2442 & ~new_n12432 ;
  assign new_n12434 = ~new_n2375 & ~new_n2402 ;
  assign new_n12435 = lo0129 & new_n2402 ;
  assign new_n12436 = ~new_n12434 & ~new_n12435 ;
  assign new_n12437 = ~new_n2442 & ~new_n12436 ;
  assign new_n12438 = ~new_n12433 & ~new_n12437 ;
  assign new_n12439 = new_n2265 & ~new_n12438 ;
  assign new_n12440 = lo0865 & ~new_n2265 ;
  assign new_n12441 = ~new_n12439 & ~new_n12440 ;
  assign new_n12442 = ~new_n12429 & ~new_n12441 ;
  assign new_n12443 = ~new_n12420 & new_n12442 ;
  assign new_n12444 = ~new_n12383 & new_n12443 ;
  assign new_n12445 = new_n2414 & new_n2442 ;
  assign new_n12446 = lo0866 & new_n12445 ;
  assign new_n12447 = new_n2329 & ~new_n2402 ;
  assign new_n12448 = ~new_n2442 & ~new_n12447 ;
  assign new_n12449 = ~new_n12446 & ~new_n12448 ;
  assign new_n12450 = new_n2265 & ~new_n12449 ;
  assign new_n12451 = lo0867 & ~new_n2265 ;
  assign new_n12452 = ~new_n12450 & ~new_n12451 ;
  assign new_n12453 = lo0868 & ~new_n2265 ;
  assign new_n12454 = ~new_n2443 & ~new_n12445 ;
  assign new_n12455 = ~new_n2356 & ~new_n2442 ;
  assign new_n12456 = lo0869 & new_n2442 ;
  assign new_n12457 = ~new_n12455 & ~new_n12456 ;
  assign new_n12458 = ~new_n12454 & ~new_n12457 ;
  assign new_n12459 = new_n2265 & new_n12458 ;
  assign new_n12460 = ~new_n12453 & ~new_n12459 ;
  assign new_n12461 = lo0870 & ~new_n2265 ;
  assign new_n12462 = ~lo0871 & new_n2442 ;
  assign new_n12463 = new_n2305 & ~new_n2442 ;
  assign new_n12464 = ~new_n12462 & ~new_n12463 ;
  assign new_n12465 = ~new_n12454 & new_n12464 ;
  assign new_n12466 = new_n2265 & new_n12465 ;
  assign new_n12467 = ~new_n12461 & ~new_n12466 ;
  assign new_n12468 = new_n12460 & new_n12467 ;
  assign new_n12469 = ~new_n12420 & ~new_n12468 ;
  assign new_n12470 = new_n12383 & ~new_n12469 ;
  assign new_n12471 = lo1291 & new_n2262 ;
  assign new_n12472 = lo1292 & new_n12471 ;
  assign new_n12473 = ~new_n12420 & new_n12472 ;
  assign new_n12474 = ~new_n12468 & new_n12473 ;
  assign new_n12475 = new_n12442 & ~new_n12474 ;
  assign new_n12476 = ~new_n12470 & new_n12475 ;
  assign new_n12477 = new_n12329 & new_n12452 ;
  assign new_n12478 = ~new_n12476 & new_n12477 ;
  assign new_n12479 = ~new_n12329 & ~new_n12452 ;
  assign new_n12480 = ~new_n12420 & ~new_n12460 ;
  assign new_n12481 = new_n12383 & ~new_n12480 ;
  assign new_n12482 = new_n12467 & ~new_n12472 ;
  assign new_n12483 = new_n12480 & ~new_n12482 ;
  assign new_n12484 = new_n12442 & ~new_n12483 ;
  assign new_n12485 = ~new_n12481 & new_n12484 ;
  assign new_n12486 = ~new_n12329 & new_n12452 ;
  assign new_n12487 = ~new_n12485 & new_n12486 ;
  assign new_n12488 = ~new_n12479 & ~new_n12487 ;
  assign new_n12489 = ~new_n12478 & new_n12488 ;
  assign new_n12490 = new_n12452 & ~new_n12489 ;
  assign new_n12491 = ~new_n12452 & new_n12489 ;
  assign new_n12492 = ~new_n12490 & ~new_n12491 ;
  assign new_n12493 = ~new_n12444 & ~new_n12492 ;
  assign new_n12494 = new_n12444 & new_n12490 ;
  assign new_n12495 = new_n12376 & new_n12420 ;
  assign new_n12496 = new_n12383 & ~new_n12420 ;
  assign new_n12497 = new_n12442 & ~new_n12496 ;
  assign new_n12498 = ~new_n12495 & new_n12497 ;
  assign new_n12499 = ~new_n12452 & ~new_n12498 ;
  assign new_n12500 = ~new_n12489 & new_n12499 ;
  assign new_n12501 = new_n2455 & ~new_n12500 ;
  assign new_n12502 = ~new_n12494 & new_n12501 ;
  assign new_n12503 = ~new_n12493 & new_n12502 ;
  assign new_n12504 = new_n2446 & ~new_n12503 ;
  assign new_n12505 = ~new_n12411 & ~new_n12504 ;
  assign new_n12506 = new_n2264 & ~new_n12367 ;
  assign new_n12507 = ~new_n12357 & new_n12506 ;
  assign new_n12508 = new_n2446 & new_n12329 ;
  assign new_n12509 = ~new_n12420 & new_n12452 ;
  assign new_n12510 = ~new_n12467 & new_n12509 ;
  assign new_n12511 = ~new_n12313 & new_n12510 ;
  assign new_n12512 = ~new_n12420 & new_n12441 ;
  assign new_n12513 = new_n12420 & ~new_n12441 ;
  assign new_n12514 = ~new_n12512 & ~new_n12513 ;
  assign new_n12515 = ~new_n12429 & ~new_n12514 ;
  assign new_n12516 = new_n12511 & new_n12515 ;
  assign new_n12517 = new_n12420 & new_n12452 ;
  assign new_n12518 = new_n2264 & new_n12517 ;
  assign new_n12519 = new_n12515 & new_n12518 ;
  assign new_n12520 = ~new_n12516 & ~new_n12519 ;
  assign new_n12521 = new_n12508 & ~new_n12520 ;
  assign new_n12522 = ~new_n2446 & ~new_n12329 ;
  assign new_n12523 = ~new_n12460 & new_n12467 ;
  assign new_n12524 = new_n12429 & new_n12441 ;
  assign new_n12525 = new_n12523 & new_n12524 ;
  assign new_n12526 = new_n2446 & ~new_n12329 ;
  assign new_n12527 = new_n12517 & new_n12526 ;
  assign new_n12528 = new_n12525 & new_n12527 ;
  assign new_n12529 = ~new_n12522 & ~new_n12528 ;
  assign new_n12530 = ~new_n12521 & new_n12529 ;
  assign new_n12531 = new_n2446 & ~new_n12530 ;
  assign new_n12532 = ~new_n2446 & new_n12530 ;
  assign new_n12533 = ~new_n12531 & ~new_n12532 ;
  assign new_n12534 = new_n12507 & ~new_n12533 ;
  assign new_n12535 = ~new_n12507 & new_n12531 ;
  assign new_n12536 = new_n12357 & new_n12368 ;
  assign new_n12537 = new_n12325 & ~new_n12376 ;
  assign new_n12538 = new_n12536 & ~new_n12537 ;
  assign new_n12539 = ~new_n2263 & ~new_n12325 ;
  assign new_n12540 = ~new_n12357 & ~new_n12539 ;
  assign new_n12541 = ~new_n12538 & ~new_n12540 ;
  assign new_n12542 = ~new_n2446 & ~new_n12541 ;
  assign new_n12543 = ~new_n12530 & new_n12542 ;
  assign new_n12544 = ~new_n12535 & ~new_n12543 ;
  assign new_n12545 = ~new_n12534 & new_n12544 ;
  assign new_n12546 = new_n2455 & ~new_n12545 ;
  assign new_n12547 = new_n2264 & new_n12329 ;
  assign new_n12548 = ~new_n2446 & new_n12547 ;
  assign new_n12549 = ~new_n12429 & new_n12441 ;
  assign new_n12550 = new_n12429 & ~new_n12441 ;
  assign new_n12551 = ~new_n12549 & ~new_n12550 ;
  assign new_n12552 = ~new_n12329 & ~new_n12551 ;
  assign new_n12553 = new_n12420 & ~new_n12452 ;
  assign new_n12554 = new_n12329 & ~new_n12524 ;
  assign new_n12555 = new_n12553 & ~new_n12554 ;
  assign new_n12556 = ~new_n12552 & new_n12555 ;
  assign new_n12557 = ~new_n12509 & ~new_n12556 ;
  assign new_n12558 = new_n2446 & ~new_n12557 ;
  assign new_n12559 = ~new_n12548 & ~new_n12558 ;
  assign new_n12560 = new_n12405 & ~new_n12559 ;
  assign new_n12561 = ~new_n12402 & ~new_n12560 ;
  assign new_n12562 = ~new_n12546 & new_n12561 ;
  assign new_n12563 = new_n2454 & ~new_n12562 ;
  assign new_n12564 = ~new_n2454 & new_n12562 ;
  assign new_n12565 = ~new_n12563 & ~new_n12564 ;
  assign new_n12566 = ~new_n2446 & ~new_n12565 ;
  assign new_n12567 = new_n2446 & new_n12563 ;
  assign new_n12568 = ~new_n12420 & ~new_n12549 ;
  assign new_n12569 = new_n12524 & new_n12553 ;
  assign new_n12570 = new_n12329 & ~new_n12569 ;
  assign new_n12571 = ~new_n12568 & new_n12570 ;
  assign new_n12572 = new_n2446 & ~new_n12571 ;
  assign new_n12573 = new_n12325 & new_n12386 ;
  assign new_n12574 = ~lo1292 & lo1293 ;
  assign new_n12575 = lo1292 & ~lo1293 ;
  assign new_n12576 = ~new_n12574 & ~new_n12575 ;
  assign new_n12577 = ~lo1291 & ~lo1294 ;
  assign new_n12578 = ~new_n12576 & new_n12577 ;
  assign new_n12579 = new_n12573 & new_n12578 ;
  assign new_n12580 = ~new_n12386 & new_n12472 ;
  assign new_n12581 = ~new_n12579 & ~new_n12580 ;
  assign new_n12582 = ~new_n12329 & ~new_n12581 ;
  assign new_n12583 = ~new_n12547 & ~new_n12582 ;
  assign new_n12584 = ~new_n2446 & ~new_n12583 ;
  assign new_n12585 = ~new_n12572 & ~new_n12584 ;
  assign new_n12586 = ~new_n2454 & ~new_n12585 ;
  assign new_n12587 = ~new_n12562 & new_n12586 ;
  assign new_n12588 = ~new_n12567 & ~new_n12587 ;
  assign new_n12589 = ~new_n12566 & new_n12588 ;
  assign new_n12590 = ~new_n2446 & new_n12329 ;
  assign new_n12591 = new_n2465 & new_n12357 ;
  assign new_n12592 = new_n12460 & ~new_n12467 ;
  assign new_n12593 = new_n2456 & new_n12443 ;
  assign new_n12594 = new_n12592 & new_n12593 ;
  assign new_n12595 = new_n12452 & new_n12594 ;
  assign new_n12596 = new_n2456 & ~new_n12420 ;
  assign new_n12597 = new_n12442 & ~new_n12596 ;
  assign new_n12598 = ~new_n12452 & ~new_n12597 ;
  assign new_n12599 = ~new_n12595 & ~new_n12598 ;
  assign new_n12600 = new_n12508 & ~new_n12599 ;
  assign new_n12601 = ~new_n12522 & ~new_n12600 ;
  assign new_n12602 = new_n2264 & ~new_n12441 ;
  assign new_n12603 = ~new_n12429 & new_n12602 ;
  assign new_n12604 = ~new_n12550 & ~new_n12603 ;
  assign new_n12605 = new_n12420 & ~new_n12604 ;
  assign new_n12606 = new_n12452 & new_n12523 ;
  assign new_n12607 = new_n12376 & new_n12606 ;
  assign new_n12608 = new_n2456 & ~new_n12452 ;
  assign new_n12609 = ~new_n12607 & ~new_n12608 ;
  assign new_n12610 = new_n12443 & ~new_n12609 ;
  assign new_n12611 = ~new_n12605 & ~new_n12610 ;
  assign new_n12612 = new_n12526 & ~new_n12611 ;
  assign new_n12613 = new_n12601 & ~new_n12612 ;
  assign new_n12614 = new_n2446 & ~new_n12613 ;
  assign new_n12615 = ~new_n2446 & new_n12613 ;
  assign new_n12616 = ~new_n12614 & ~new_n12615 ;
  assign new_n12617 = new_n12591 & ~new_n12616 ;
  assign new_n12618 = ~new_n12591 & new_n12614 ;
  assign new_n12619 = new_n2456 & new_n12325 ;
  assign new_n12620 = ~new_n12371 & ~new_n12377 ;
  assign new_n12621 = ~new_n12619 & new_n12620 ;
  assign new_n12622 = ~new_n2446 & ~new_n12621 ;
  assign new_n12623 = ~new_n12613 & new_n12622 ;
  assign new_n12624 = ~new_n12618 & ~new_n12623 ;
  assign new_n12625 = ~new_n12617 & new_n12624 ;
  assign new_n12626 = new_n2455 & ~new_n12625 ;
  assign new_n12627 = ~new_n12420 & new_n12549 ;
  assign new_n12628 = new_n12420 & ~new_n12551 ;
  assign new_n12629 = ~new_n12627 & ~new_n12628 ;
  assign new_n12630 = ~new_n12477 & ~new_n12479 ;
  assign new_n12631 = ~new_n12420 & ~new_n12630 ;
  assign new_n12632 = new_n12420 & new_n12479 ;
  assign new_n12633 = new_n12486 & new_n12512 ;
  assign new_n12634 = ~new_n12632 & ~new_n12633 ;
  assign new_n12635 = ~new_n12631 & new_n12634 ;
  assign new_n12636 = new_n12452 & ~new_n12635 ;
  assign new_n12637 = ~new_n12452 & new_n12635 ;
  assign new_n12638 = ~new_n12636 & ~new_n12637 ;
  assign new_n12639 = ~new_n12629 & ~new_n12638 ;
  assign new_n12640 = new_n12629 & new_n12636 ;
  assign new_n12641 = ~new_n12442 & new_n12551 ;
  assign new_n12642 = new_n12553 & ~new_n12641 ;
  assign new_n12643 = ~new_n12635 & new_n12642 ;
  assign new_n12644 = ~new_n12640 & ~new_n12643 ;
  assign new_n12645 = ~new_n12639 & new_n12644 ;
  assign new_n12646 = new_n2446 & new_n12405 ;
  assign new_n12647 = ~new_n12645 & new_n12646 ;
  assign new_n12648 = ~new_n12402 & ~new_n12647 ;
  assign new_n12649 = ~new_n12626 & new_n12648 ;
  assign new_n12650 = new_n2454 & ~new_n12649 ;
  assign new_n12651 = ~new_n2454 & new_n12649 ;
  assign new_n12652 = ~new_n12650 & ~new_n12651 ;
  assign new_n12653 = ~new_n12590 & ~new_n12652 ;
  assign new_n12654 = new_n12590 & new_n12650 ;
  assign new_n12655 = ~new_n12526 & ~new_n12590 ;
  assign new_n12656 = ~new_n2454 & new_n12655 ;
  assign new_n12657 = new_n2446 & new_n12569 ;
  assign new_n12658 = ~new_n2465 & new_n12357 ;
  assign new_n12659 = ~new_n12325 & new_n12658 ;
  assign new_n12660 = new_n12472 & new_n12659 ;
  assign new_n12661 = ~lo1292 & new_n12367 ;
  assign new_n12662 = ~lo1291 & ~new_n12661 ;
  assign new_n12663 = ~new_n12338 & ~new_n12662 ;
  assign new_n12664 = ~lo1293 & ~new_n12663 ;
  assign new_n12665 = ~new_n12659 & new_n12664 ;
  assign new_n12666 = new_n12358 & ~new_n12574 ;
  assign new_n12667 = ~new_n12665 & ~new_n12666 ;
  assign new_n12668 = ~lo1294 & ~new_n12667 ;
  assign new_n12669 = ~new_n12660 & ~new_n12668 ;
  assign new_n12670 = ~new_n2446 & ~new_n12669 ;
  assign new_n12671 = ~new_n12657 & ~new_n12670 ;
  assign new_n12672 = new_n12656 & ~new_n12671 ;
  assign new_n12673 = ~new_n12649 & new_n12672 ;
  assign new_n12674 = ~new_n12654 & ~new_n12673 ;
  assign new_n12675 = ~new_n12653 & new_n12674 ;
  assign new_n12676 = new_n2456 & new_n12368 ;
  assign new_n12677 = new_n12357 & ~new_n12676 ;
  assign new_n12678 = new_n12325 & ~new_n12677 ;
  assign new_n12679 = new_n12370 & new_n12376 ;
  assign new_n12680 = ~new_n12678 & ~new_n12679 ;
  assign new_n12681 = new_n2450 & ~new_n12680 ;
  assign new_n12682 = ~new_n12358 & ~new_n12395 ;
  assign new_n12683 = new_n12325 & ~new_n12682 ;
  assign new_n12684 = new_n2262 & new_n12339 ;
  assign new_n12685 = ~lo1292 & new_n12387 ;
  assign new_n12686 = ~lo1294 & ~new_n12685 ;
  assign new_n12687 = ~new_n12684 & new_n12686 ;
  assign new_n12688 = new_n12683 & new_n12687 ;
  assign new_n12689 = ~new_n12370 & ~new_n12682 ;
  assign new_n12690 = new_n2262 & ~new_n12663 ;
  assign new_n12691 = ~new_n12689 & new_n12690 ;
  assign new_n12692 = ~new_n12688 & ~new_n12691 ;
  assign new_n12693 = ~new_n2450 & ~new_n12692 ;
  assign new_n12694 = ~new_n12681 & ~new_n12693 ;
  assign new_n12695 = ~new_n12404 & ~new_n12405 ;
  assign new_n12696 = new_n12522 & new_n12695 ;
  assign new_n12697 = ~new_n12694 & new_n12696 ;
  assign new_n12698 = ~new_n2450 & new_n12329 ;
  assign new_n12699 = ~new_n2454 & new_n12509 ;
  assign new_n12700 = ~new_n12549 & new_n12699 ;
  assign new_n12701 = ~new_n12524 & ~new_n12550 ;
  assign new_n12702 = new_n12420 & ~new_n12701 ;
  assign new_n12703 = ~new_n12549 & ~new_n12702 ;
  assign new_n12704 = ~new_n12452 & ~new_n12703 ;
  assign new_n12705 = ~new_n12509 & ~new_n12704 ;
  assign new_n12706 = new_n2454 & ~new_n12705 ;
  assign new_n12707 = ~new_n12700 & ~new_n12706 ;
  assign new_n12708 = new_n12698 & ~new_n12707 ;
  assign new_n12709 = new_n2454 & ~new_n12329 ;
  assign new_n12710 = ~new_n12523 & new_n12605 ;
  assign new_n12711 = ~new_n12429 & ~new_n12602 ;
  assign new_n12712 = new_n12420 & ~new_n12711 ;
  assign new_n12713 = new_n12376 & new_n12443 ;
  assign new_n12714 = ~new_n12712 & ~new_n12713 ;
  assign new_n12715 = new_n12523 & ~new_n12714 ;
  assign new_n12716 = ~new_n12710 & ~new_n12715 ;
  assign new_n12717 = new_n2450 & new_n12452 ;
  assign new_n12718 = ~new_n12716 & new_n12717 ;
  assign new_n12719 = ~new_n12441 & new_n12509 ;
  assign new_n12720 = ~new_n12420 & ~new_n12452 ;
  assign new_n12721 = new_n12442 & new_n12553 ;
  assign new_n12722 = ~new_n12720 & ~new_n12721 ;
  assign new_n12723 = ~new_n12719 & new_n12722 ;
  assign new_n12724 = ~new_n2450 & ~new_n12723 ;
  assign new_n12725 = ~new_n12718 & ~new_n12724 ;
  assign new_n12726 = new_n12709 & ~new_n12725 ;
  assign new_n12727 = ~new_n12708 & ~new_n12726 ;
  assign new_n12728 = new_n2446 & ~new_n12727 ;
  assign new_n12729 = ~new_n12697 & ~new_n12728 ;
  assign new_n12730 = ~lo0875 & ~lo0876 ;
  assign new_n12731 = lo0872 & ~lo0873 ;
  assign new_n12732 = ~lo0874 & new_n12731 ;
  assign new_n12733 = new_n12730 & new_n12732 ;
  assign new_n12734 = new_n12729 & new_n12733 ;
  assign new_n12735 = ~new_n12675 & new_n12734 ;
  assign new_n12736 = new_n12589 & new_n12735 ;
  assign new_n12737 = ~new_n12420 & new_n12550 ;
  assign new_n12738 = ~new_n12569 & ~new_n12737 ;
  assign new_n12739 = new_n12698 & ~new_n12738 ;
  assign new_n12740 = new_n12452 & new_n12550 ;
  assign new_n12741 = ~new_n12429 & ~new_n12452 ;
  assign new_n12742 = new_n12420 & ~new_n12741 ;
  assign new_n12743 = ~new_n12740 & ~new_n12742 ;
  assign new_n12744 = new_n12511 & new_n12549 ;
  assign new_n12745 = new_n12442 & new_n12509 ;
  assign new_n12746 = new_n12334 & new_n12592 ;
  assign new_n12747 = new_n12745 & new_n12746 ;
  assign new_n12748 = ~new_n12598 & ~new_n12747 ;
  assign new_n12749 = ~new_n12744 & new_n12748 ;
  assign new_n12750 = new_n2450 & new_n12329 ;
  assign new_n12751 = ~new_n12749 & new_n12750 ;
  assign new_n12752 = ~new_n2450 & ~new_n12329 ;
  assign new_n12753 = new_n12460 & ~new_n12604 ;
  assign new_n12754 = new_n2263 & new_n12443 ;
  assign new_n12755 = ~new_n12712 & ~new_n12754 ;
  assign new_n12756 = new_n12523 & ~new_n12755 ;
  assign new_n12757 = ~new_n12753 & ~new_n12756 ;
  assign new_n12758 = new_n12452 & ~new_n12757 ;
  assign new_n12759 = ~new_n12460 & ~new_n12467 ;
  assign new_n12760 = new_n12452 & ~new_n12759 ;
  assign new_n12761 = new_n2264 & new_n12442 ;
  assign new_n12762 = new_n12420 & new_n12761 ;
  assign new_n12763 = ~new_n12550 & ~new_n12762 ;
  assign new_n12764 = ~new_n12760 & ~new_n12763 ;
  assign new_n12765 = ~new_n12460 & new_n12737 ;
  assign new_n12766 = ~new_n12764 & ~new_n12765 ;
  assign new_n12767 = ~new_n12758 & new_n12766 ;
  assign new_n12768 = new_n2450 & ~new_n12329 ;
  assign new_n12769 = ~new_n12767 & new_n12768 ;
  assign new_n12770 = ~new_n12752 & ~new_n12769 ;
  assign new_n12771 = ~new_n12751 & new_n12770 ;
  assign new_n12772 = new_n2450 & ~new_n12771 ;
  assign new_n12773 = ~new_n2450 & new_n12771 ;
  assign new_n12774 = ~new_n12772 & ~new_n12773 ;
  assign new_n12775 = ~new_n12743 & ~new_n12774 ;
  assign new_n12776 = new_n12743 & new_n12772 ;
  assign new_n12777 = new_n12509 & ~new_n12551 ;
  assign new_n12778 = ~new_n12420 & ~new_n12429 ;
  assign new_n12779 = new_n12420 & ~new_n12549 ;
  assign new_n12780 = ~new_n12778 & ~new_n12779 ;
  assign new_n12781 = ~new_n12452 & ~new_n12780 ;
  assign new_n12782 = ~new_n12777 & ~new_n12781 ;
  assign new_n12783 = ~new_n2450 & ~new_n12782 ;
  assign new_n12784 = ~new_n12771 & new_n12783 ;
  assign new_n12785 = ~new_n12776 & ~new_n12784 ;
  assign new_n12786 = ~new_n12775 & new_n12785 ;
  assign new_n12787 = new_n2446 & new_n2454 ;
  assign new_n12788 = ~new_n12786 & new_n12787 ;
  assign new_n12789 = ~new_n2446 & ~new_n2454 ;
  assign new_n12790 = ~lo1291 & lo1294 ;
  assign new_n12791 = ~lo1291 & ~new_n12790 ;
  assign new_n12792 = new_n12339 & new_n12387 ;
  assign new_n12793 = new_n12791 & ~new_n12792 ;
  assign new_n12794 = new_n12369 & new_n12793 ;
  assign new_n12795 = ~new_n12325 & ~new_n12376 ;
  assign new_n12796 = ~new_n12357 & ~new_n12795 ;
  assign new_n12797 = ~new_n2465 & new_n12367 ;
  assign new_n12798 = new_n12796 & new_n12797 ;
  assign new_n12799 = ~new_n12794 & ~new_n12798 ;
  assign new_n12800 = ~new_n2446 & new_n2454 ;
  assign new_n12801 = new_n12768 & new_n12800 ;
  assign new_n12802 = ~new_n12799 & new_n12801 ;
  assign new_n12803 = ~new_n12789 & ~new_n12802 ;
  assign new_n12804 = ~new_n12788 & new_n12803 ;
  assign new_n12805 = new_n2454 & ~new_n12804 ;
  assign new_n12806 = ~new_n2454 & new_n12804 ;
  assign new_n12807 = ~new_n12805 & ~new_n12806 ;
  assign new_n12808 = new_n12739 & ~new_n12807 ;
  assign new_n12809 = ~new_n12739 & new_n12805 ;
  assign new_n12810 = ~lo1291 & ~new_n12367 ;
  assign new_n12811 = ~lo1292 & ~lo1293 ;
  assign new_n12812 = ~new_n12810 & new_n12811 ;
  assign new_n12813 = ~new_n12339 & ~new_n12812 ;
  assign new_n12814 = ~lo1294 & ~new_n12813 ;
  assign new_n12815 = ~new_n12386 & new_n12814 ;
  assign new_n12816 = ~lo1291 & lo1293 ;
  assign new_n12817 = lo1292 & new_n12816 ;
  assign new_n12818 = ~lo1291 & ~new_n12817 ;
  assign new_n12819 = ~lo1294 & ~new_n12818 ;
  assign new_n12820 = new_n12325 & new_n12819 ;
  assign new_n12821 = ~lo1292 & new_n12816 ;
  assign new_n12822 = lo1291 & ~lo1293 ;
  assign new_n12823 = lo1292 & new_n12822 ;
  assign new_n12824 = ~new_n12821 & ~new_n12823 ;
  assign new_n12825 = ~lo1294 & ~new_n12824 ;
  assign new_n12826 = new_n12395 & new_n12825 ;
  assign new_n12827 = ~new_n12820 & ~new_n12826 ;
  assign new_n12828 = new_n12357 & ~new_n12827 ;
  assign new_n12829 = ~new_n12815 & ~new_n12828 ;
  assign new_n12830 = ~new_n2454 & new_n12752 ;
  assign new_n12831 = ~new_n12829 & new_n12830 ;
  assign new_n12832 = ~new_n12804 & new_n12831 ;
  assign new_n12833 = ~new_n12809 & ~new_n12832 ;
  assign new_n12834 = ~new_n12808 & new_n12833 ;
  assign new_n12835 = new_n12376 & ~new_n12467 ;
  assign new_n12836 = new_n2264 & new_n12467 ;
  assign new_n12837 = ~new_n12835 & ~new_n12836 ;
  assign new_n12838 = new_n12460 & ~new_n12837 ;
  assign new_n12839 = new_n12745 & new_n12838 ;
  assign new_n12840 = ~new_n12442 & ~new_n12452 ;
  assign new_n12841 = ~new_n12740 & ~new_n12840 ;
  assign new_n12842 = ~new_n12839 & new_n12841 ;
  assign new_n12843 = ~new_n12744 & new_n12842 ;
  assign new_n12844 = new_n12508 & ~new_n12843 ;
  assign new_n12845 = new_n12420 & new_n12429 ;
  assign new_n12846 = ~new_n12443 & ~new_n12845 ;
  assign new_n12847 = new_n12376 & ~new_n12420 ;
  assign new_n12848 = new_n12420 & new_n12441 ;
  assign new_n12849 = ~new_n12847 & ~new_n12848 ;
  assign new_n12850 = new_n12606 & ~new_n12849 ;
  assign new_n12851 = ~new_n12846 & new_n12850 ;
  assign new_n12852 = new_n12526 & new_n12851 ;
  assign new_n12853 = ~new_n12522 & ~new_n12852 ;
  assign new_n12854 = ~new_n12844 & new_n12853 ;
  assign new_n12855 = new_n2446 & ~new_n12854 ;
  assign new_n12856 = ~new_n2446 & new_n12854 ;
  assign new_n12857 = ~new_n12855 & ~new_n12856 ;
  assign new_n12858 = new_n12591 & ~new_n12857 ;
  assign new_n12859 = ~new_n12591 & new_n12855 ;
  assign new_n12860 = new_n12387 & new_n12391 ;
  assign new_n12861 = ~new_n12325 & new_n12860 ;
  assign new_n12862 = new_n12860 & ~new_n12861 ;
  assign new_n12863 = new_n12357 & ~new_n12368 ;
  assign new_n12864 = ~new_n12862 & new_n12863 ;
  assign new_n12865 = ~new_n12358 & ~new_n12370 ;
  assign new_n12866 = new_n12860 & ~new_n12865 ;
  assign new_n12867 = new_n12370 & ~new_n12860 ;
  assign new_n12868 = ~new_n12866 & ~new_n12867 ;
  assign new_n12869 = ~new_n12864 & new_n12868 ;
  assign new_n12870 = ~new_n12357 & new_n12368 ;
  assign new_n12871 = new_n12869 & new_n12870 ;
  assign new_n12872 = new_n12357 & ~new_n12869 ;
  assign new_n12873 = new_n12376 & new_n12870 ;
  assign new_n12874 = ~new_n12869 & new_n12873 ;
  assign new_n12875 = ~new_n12872 & ~new_n12874 ;
  assign new_n12876 = ~new_n12871 & new_n12875 ;
  assign new_n12877 = ~new_n2446 & ~new_n12876 ;
  assign new_n12878 = ~new_n12854 & new_n12877 ;
  assign new_n12879 = ~new_n12859 & ~new_n12878 ;
  assign new_n12880 = ~new_n12858 & new_n12879 ;
  assign new_n12881 = new_n2455 & ~new_n12880 ;
  assign new_n12882 = ~new_n12778 & ~new_n12845 ;
  assign new_n12883 = new_n12329 & ~new_n12882 ;
  assign new_n12884 = ~new_n12329 & new_n12845 ;
  assign new_n12885 = ~new_n12883 & ~new_n12884 ;
  assign new_n12886 = new_n12441 & ~new_n12885 ;
  assign new_n12887 = ~new_n12420 & new_n12429 ;
  assign new_n12888 = new_n12429 & ~new_n12887 ;
  assign new_n12889 = ~new_n12329 & ~new_n12441 ;
  assign new_n12890 = ~new_n12888 & new_n12889 ;
  assign new_n12891 = ~new_n12886 & ~new_n12890 ;
  assign new_n12892 = ~new_n12452 & ~new_n12891 ;
  assign new_n12893 = new_n12329 & new_n12443 ;
  assign new_n12894 = ~new_n12420 & ~new_n12524 ;
  assign new_n12895 = ~new_n12329 & ~new_n12894 ;
  assign new_n12896 = ~new_n12893 & ~new_n12895 ;
  assign new_n12897 = new_n12452 & ~new_n12896 ;
  assign new_n12898 = ~new_n12892 & ~new_n12897 ;
  assign new_n12899 = new_n2446 & ~new_n12898 ;
  assign new_n12900 = ~new_n12522 & ~new_n12899 ;
  assign new_n12901 = new_n12405 & ~new_n12900 ;
  assign new_n12902 = ~new_n12402 & ~new_n12901 ;
  assign new_n12903 = ~new_n12881 & new_n12902 ;
  assign new_n12904 = new_n2454 & ~new_n12903 ;
  assign new_n12905 = ~new_n2454 & new_n12903 ;
  assign new_n12906 = ~new_n12904 & ~new_n12905 ;
  assign new_n12907 = new_n2446 & ~new_n12906 ;
  assign new_n12908 = ~new_n2446 & new_n12904 ;
  assign new_n12909 = lo1292 & new_n12387 ;
  assign new_n12910 = ~lo1291 & new_n12909 ;
  assign new_n12911 = ~new_n12386 & new_n12910 ;
  assign new_n12912 = ~new_n12816 & ~new_n12822 ;
  assign new_n12913 = ~lo1292 & ~lo1294 ;
  assign new_n12914 = ~new_n12912 & new_n12913 ;
  assign new_n12915 = new_n12395 & new_n12914 ;
  assign new_n12916 = new_n12338 & new_n12387 ;
  assign new_n12917 = new_n12325 & new_n12916 ;
  assign new_n12918 = ~new_n12915 & ~new_n12917 ;
  assign new_n12919 = new_n12357 & ~new_n12918 ;
  assign new_n12920 = ~new_n12911 & ~new_n12919 ;
  assign new_n12921 = ~new_n2446 & ~new_n12920 ;
  assign new_n12922 = ~new_n12443 & ~new_n12569 ;
  assign new_n12923 = new_n2446 & ~new_n12922 ;
  assign new_n12924 = ~new_n12921 & ~new_n12923 ;
  assign new_n12925 = new_n12656 & ~new_n12924 ;
  assign new_n12926 = ~new_n12903 & new_n12925 ;
  assign new_n12927 = ~new_n12908 & ~new_n12926 ;
  assign new_n12928 = ~new_n12907 & new_n12927 ;
  assign new_n12929 = ~new_n12834 & ~new_n12928 ;
  assign new_n12930 = new_n12736 & new_n12929 ;
  assign new_n12931 = ~new_n12367 & ~new_n12441 ;
  assign new_n12932 = ~new_n2454 & new_n12778 ;
  assign new_n12933 = new_n12429 & new_n12452 ;
  assign new_n12934 = new_n2454 & new_n12933 ;
  assign new_n12935 = ~new_n12932 & ~new_n12934 ;
  assign new_n12936 = new_n12508 & new_n12695 ;
  assign new_n12937 = ~new_n12935 & new_n12936 ;
  assign new_n12938 = new_n12931 & new_n12937 ;
  assign new_n12939 = ~new_n12367 & ~new_n12442 ;
  assign new_n12940 = new_n2446 & ~new_n2450 ;
  assign new_n12941 = ~new_n2450 & ~new_n12940 ;
  assign new_n12942 = ~new_n12329 & new_n12940 ;
  assign new_n12943 = ~new_n12941 & ~new_n12942 ;
  assign new_n12944 = ~new_n12420 & new_n12943 ;
  assign new_n12945 = new_n12940 & ~new_n12944 ;
  assign new_n12946 = new_n12940 & ~new_n12943 ;
  assign new_n12947 = lo1292 & ~new_n12460 ;
  assign new_n12948 = ~lo1292 & ~new_n12367 ;
  assign new_n12949 = ~new_n12947 & ~new_n12948 ;
  assign new_n12950 = new_n2456 & ~new_n12949 ;
  assign new_n12951 = new_n12329 & ~new_n12452 ;
  assign new_n12952 = new_n2446 & ~new_n12951 ;
  assign new_n12953 = ~new_n12443 & ~new_n12952 ;
  assign new_n12954 = new_n12508 & ~new_n12953 ;
  assign new_n12955 = ~new_n12329 & new_n12369 ;
  assign new_n12956 = new_n2456 & new_n12955 ;
  assign new_n12957 = ~new_n12508 & ~new_n12952 ;
  assign new_n12958 = new_n12508 & new_n12952 ;
  assign new_n12959 = ~new_n12957 & ~new_n12958 ;
  assign new_n12960 = new_n12956 & ~new_n12959 ;
  assign new_n12961 = ~new_n12956 & new_n12958 ;
  assign new_n12962 = ~new_n12960 & ~new_n12961 ;
  assign new_n12963 = ~new_n12508 & new_n12952 ;
  assign new_n12964 = ~new_n2264 & ~new_n12429 ;
  assign new_n12965 = ~new_n12441 & ~new_n12964 ;
  assign new_n12966 = ~new_n12367 & new_n12965 ;
  assign new_n12967 = new_n12420 & ~new_n12460 ;
  assign new_n12968 = new_n2456 & ~new_n12441 ;
  assign new_n12969 = ~new_n12949 & new_n12968 ;
  assign new_n12970 = new_n12452 & new_n12467 ;
  assign new_n12971 = new_n12967 & ~new_n12970 ;
  assign new_n12972 = new_n12420 & ~new_n12971 ;
  assign new_n12973 = new_n12429 & ~new_n12972 ;
  assign new_n12974 = ~new_n12967 & ~new_n12973 ;
  assign new_n12975 = ~new_n12972 & new_n12974 ;
  assign new_n12976 = new_n12972 & ~new_n12974 ;
  assign new_n12977 = ~new_n12975 & ~new_n12976 ;
  assign new_n12978 = new_n12969 & ~new_n12977 ;
  assign new_n12979 = ~new_n12969 & new_n12976 ;
  assign new_n12980 = ~new_n12367 & new_n12429 ;
  assign new_n12981 = ~new_n12367 & new_n12602 ;
  assign new_n12982 = ~new_n12367 & new_n12441 ;
  assign new_n12983 = ~new_n12981 & ~new_n12982 ;
  assign new_n12984 = ~new_n12429 & ~new_n12983 ;
  assign new_n12985 = ~new_n12980 & ~new_n12984 ;
  assign new_n12986 = new_n12972 & new_n12974 ;
  assign new_n12987 = ~new_n12985 & new_n12986 ;
  assign new_n12988 = ~new_n12979 & ~new_n12987 ;
  assign new_n12989 = ~new_n12978 & new_n12988 ;
  assign new_n12990 = ~new_n12967 & ~new_n12989 ;
  assign new_n12991 = new_n12967 & new_n12989 ;
  assign new_n12992 = ~new_n12990 & ~new_n12991 ;
  assign new_n12993 = new_n12966 & ~new_n12992 ;
  assign new_n12994 = ~new_n12966 & new_n12990 ;
  assign new_n12995 = new_n12967 & new_n12981 ;
  assign new_n12996 = ~new_n12989 & new_n12995 ;
  assign new_n12997 = ~new_n12994 & ~new_n12996 ;
  assign new_n12998 = ~new_n12993 & new_n12997 ;
  assign new_n12999 = new_n12963 & ~new_n12998 ;
  assign new_n13000 = new_n12962 & ~new_n12999 ;
  assign new_n13001 = ~new_n12954 & ~new_n13000 ;
  assign new_n13002 = new_n12954 & new_n13000 ;
  assign new_n13003 = ~new_n13001 & ~new_n13002 ;
  assign new_n13004 = new_n12950 & ~new_n13003 ;
  assign new_n13005 = ~new_n12950 & new_n13001 ;
  assign new_n13006 = ~new_n12441 & new_n12592 ;
  assign new_n13007 = new_n12596 & new_n13006 ;
  assign new_n13008 = new_n12954 & new_n13007 ;
  assign new_n13009 = ~new_n13000 & new_n13008 ;
  assign new_n13010 = ~new_n13005 & ~new_n13009 ;
  assign new_n13011 = ~new_n13004 & new_n13010 ;
  assign new_n13012 = new_n12946 & new_n13011 ;
  assign new_n13013 = ~new_n12940 & new_n12943 ;
  assign new_n13014 = ~new_n12946 & ~new_n13013 ;
  assign new_n13015 = ~new_n13011 & ~new_n13014 ;
  assign new_n13016 = ~new_n12940 & ~new_n12943 ;
  assign new_n13017 = ~new_n12329 & ~new_n12367 ;
  assign new_n13018 = new_n13016 & new_n13017 ;
  assign new_n13019 = ~new_n13015 & ~new_n13018 ;
  assign new_n13020 = ~new_n13012 & new_n13019 ;
  assign new_n13021 = ~new_n12945 & ~new_n13020 ;
  assign new_n13022 = new_n12945 & new_n13020 ;
  assign new_n13023 = ~new_n13021 & ~new_n13022 ;
  assign new_n13024 = new_n12939 & ~new_n13023 ;
  assign new_n13025 = ~new_n12939 & new_n13021 ;
  assign new_n13026 = ~new_n12460 & new_n12945 ;
  assign new_n13027 = ~new_n13020 & new_n13026 ;
  assign new_n13028 = ~new_n13025 & ~new_n13027 ;
  assign new_n13029 = ~new_n13024 & new_n13028 ;
  assign new_n13030 = new_n12329 & new_n12720 ;
  assign new_n13031 = ~new_n12429 & new_n13030 ;
  assign new_n13032 = ~new_n2450 & ~new_n13031 ;
  assign new_n13033 = ~new_n12329 & ~new_n12420 ;
  assign new_n13034 = new_n12452 & new_n13033 ;
  assign new_n13035 = new_n2450 & ~new_n13034 ;
  assign new_n13036 = new_n2446 & ~new_n13035 ;
  assign new_n13037 = ~new_n13032 & new_n13036 ;
  assign new_n13038 = new_n2454 & ~new_n13037 ;
  assign new_n13039 = ~new_n12452 & new_n12940 ;
  assign new_n13040 = new_n12429 & new_n13039 ;
  assign new_n13041 = ~new_n2454 & ~new_n13040 ;
  assign new_n13042 = ~new_n13038 & ~new_n13041 ;
  assign new_n13043 = ~new_n12329 & new_n12523 ;
  assign new_n13044 = new_n12429 & new_n12517 ;
  assign new_n13045 = new_n13043 & new_n13044 ;
  assign new_n13046 = new_n12329 & new_n12509 ;
  assign new_n13047 = new_n12441 & ~new_n12467 ;
  assign new_n13048 = new_n13046 & new_n13047 ;
  assign new_n13049 = ~new_n13045 & ~new_n13048 ;
  assign new_n13050 = new_n2455 & ~new_n13049 ;
  assign new_n13051 = new_n12452 & ~new_n13033 ;
  assign new_n13052 = new_n12442 & new_n13051 ;
  assign new_n13053 = ~new_n12442 & new_n12553 ;
  assign new_n13054 = ~new_n13051 & ~new_n13053 ;
  assign new_n13055 = new_n2454 & ~new_n13054 ;
  assign new_n13056 = ~new_n13052 & new_n13055 ;
  assign new_n13057 = ~new_n12329 & ~new_n13056 ;
  assign new_n13058 = new_n2454 & ~new_n12477 ;
  assign new_n13059 = ~new_n12420 & ~new_n13058 ;
  assign new_n13060 = ~new_n13057 & ~new_n13059 ;
  assign new_n13061 = ~new_n2450 & ~new_n13060 ;
  assign new_n13062 = ~new_n13050 & ~new_n13061 ;
  assign new_n13063 = new_n2446 & ~new_n13062 ;
  assign new_n13064 = ~new_n13042 & ~new_n13063 ;
  assign new_n13065 = ~new_n2446 & ~new_n2450 ;
  assign new_n13066 = ~new_n2454 & new_n13064 ;
  assign new_n13067 = ~new_n13063 & ~new_n13066 ;
  assign new_n13068 = ~new_n13065 & ~new_n13067 ;
  assign new_n13069 = new_n13064 & ~new_n13068 ;
  assign new_n13070 = new_n12940 & new_n13051 ;
  assign new_n13071 = new_n13069 & ~new_n13070 ;
  assign new_n13072 = new_n12441 & new_n13067 ;
  assign new_n13073 = ~new_n12367 & ~new_n13064 ;
  assign new_n13074 = new_n13072 & new_n13073 ;
  assign new_n13075 = new_n13064 & new_n13067 ;
  assign new_n13076 = ~new_n13067 & new_n13073 ;
  assign new_n13077 = ~new_n13075 & ~new_n13076 ;
  assign new_n13078 = ~new_n13074 & new_n13077 ;
  assign new_n13079 = new_n13071 & ~new_n13078 ;
  assign new_n13080 = ~new_n13029 & new_n13079 ;
  assign new_n13081 = ~lo1293 & new_n12341 ;
  assign new_n13082 = ~new_n12386 & new_n13081 ;
  assign new_n13083 = new_n12573 & new_n12909 ;
  assign new_n13084 = ~new_n13082 & ~new_n13083 ;
  assign new_n13085 = ~new_n12329 & ~new_n13084 ;
  assign new_n13086 = ~new_n13069 & ~new_n13078 ;
  assign new_n13087 = new_n13069 & new_n13078 ;
  assign new_n13088 = ~new_n13086 & ~new_n13087 ;
  assign new_n13089 = new_n13085 & ~new_n13088 ;
  assign new_n13090 = ~new_n13085 & new_n13086 ;
  assign new_n13091 = ~new_n13089 & ~new_n13090 ;
  assign new_n13092 = ~new_n13080 & new_n13091 ;
  assign new_n13093 = ~new_n12937 & ~new_n13092 ;
  assign new_n13094 = ~new_n12938 & ~new_n13093 ;
  assign new_n13095 = ~lo0876 & ~new_n13094 ;
  assign new_n13096 = ~new_n12357 & ~new_n12441 ;
  assign new_n13097 = new_n12937 & new_n13096 ;
  assign new_n13098 = ~new_n12357 & ~new_n12442 ;
  assign new_n13099 = lo0877 & ~new_n2265 ;
  assign new_n13100 = ~new_n2335 & ~new_n2442 ;
  assign new_n13101 = lo0878 & new_n2442 ;
  assign new_n13102 = ~new_n13100 & ~new_n13101 ;
  assign new_n13103 = ~new_n12454 & ~new_n13102 ;
  assign new_n13104 = new_n2265 & new_n13103 ;
  assign new_n13105 = ~new_n13099 & ~new_n13104 ;
  assign new_n13106 = lo1292 & ~new_n13105 ;
  assign new_n13107 = ~lo1292 & ~new_n12357 ;
  assign new_n13108 = ~new_n13106 & ~new_n13107 ;
  assign new_n13109 = new_n2456 & ~new_n13108 ;
  assign new_n13110 = ~new_n12357 & new_n12965 ;
  assign new_n13111 = new_n12968 & ~new_n13108 ;
  assign new_n13112 = ~new_n12977 & new_n13111 ;
  assign new_n13113 = new_n12976 & ~new_n13111 ;
  assign new_n13114 = ~new_n12357 & new_n12429 ;
  assign new_n13115 = ~new_n12357 & new_n12602 ;
  assign new_n13116 = ~new_n12357 & new_n12441 ;
  assign new_n13117 = ~new_n13115 & ~new_n13116 ;
  assign new_n13118 = ~new_n12429 & ~new_n13117 ;
  assign new_n13119 = ~new_n13114 & ~new_n13118 ;
  assign new_n13120 = new_n12986 & ~new_n13119 ;
  assign new_n13121 = ~new_n13113 & ~new_n13120 ;
  assign new_n13122 = ~new_n13112 & new_n13121 ;
  assign new_n13123 = ~new_n12967 & ~new_n13122 ;
  assign new_n13124 = new_n12967 & new_n13122 ;
  assign new_n13125 = ~new_n13123 & ~new_n13124 ;
  assign new_n13126 = new_n13110 & ~new_n13125 ;
  assign new_n13127 = ~new_n13110 & new_n13123 ;
  assign new_n13128 = new_n12967 & new_n13115 ;
  assign new_n13129 = ~new_n13122 & new_n13128 ;
  assign new_n13130 = ~new_n13127 & ~new_n13129 ;
  assign new_n13131 = ~new_n13126 & new_n13130 ;
  assign new_n13132 = new_n12963 & ~new_n13131 ;
  assign new_n13133 = new_n12962 & ~new_n13132 ;
  assign new_n13134 = ~new_n12954 & ~new_n13133 ;
  assign new_n13135 = new_n12954 & new_n13133 ;
  assign new_n13136 = ~new_n13134 & ~new_n13135 ;
  assign new_n13137 = new_n13109 & ~new_n13136 ;
  assign new_n13138 = ~new_n13109 & new_n13134 ;
  assign new_n13139 = new_n13008 & ~new_n13133 ;
  assign new_n13140 = ~new_n13138 & ~new_n13139 ;
  assign new_n13141 = ~new_n13137 & new_n13140 ;
  assign new_n13142 = new_n12946 & new_n13141 ;
  assign new_n13143 = ~new_n13014 & ~new_n13141 ;
  assign new_n13144 = ~new_n12329 & ~new_n12357 ;
  assign new_n13145 = new_n13016 & new_n13144 ;
  assign new_n13146 = ~new_n13143 & ~new_n13145 ;
  assign new_n13147 = ~new_n13142 & new_n13146 ;
  assign new_n13148 = ~new_n12945 & ~new_n13147 ;
  assign new_n13149 = new_n12945 & new_n13147 ;
  assign new_n13150 = ~new_n13148 & ~new_n13149 ;
  assign new_n13151 = new_n13098 & ~new_n13150 ;
  assign new_n13152 = ~new_n13098 & new_n13148 ;
  assign new_n13153 = new_n12945 & ~new_n13105 ;
  assign new_n13154 = ~new_n13147 & new_n13153 ;
  assign new_n13155 = ~new_n13152 & ~new_n13154 ;
  assign new_n13156 = ~new_n13151 & new_n13155 ;
  assign new_n13157 = ~new_n12357 & ~new_n13064 ;
  assign new_n13158 = new_n13072 & new_n13157 ;
  assign new_n13159 = ~new_n13067 & new_n13157 ;
  assign new_n13160 = ~new_n13075 & ~new_n13159 ;
  assign new_n13161 = ~new_n13158 & new_n13160 ;
  assign new_n13162 = new_n13071 & ~new_n13161 ;
  assign new_n13163 = ~new_n13156 & new_n13162 ;
  assign new_n13164 = ~new_n13069 & ~new_n13161 ;
  assign new_n13165 = new_n13069 & new_n13161 ;
  assign new_n13166 = ~new_n13164 & ~new_n13165 ;
  assign new_n13167 = new_n13085 & ~new_n13166 ;
  assign new_n13168 = ~new_n13085 & new_n13164 ;
  assign new_n13169 = ~new_n13167 & ~new_n13168 ;
  assign new_n13170 = ~new_n13163 & new_n13169 ;
  assign new_n13171 = ~new_n12937 & ~new_n13170 ;
  assign new_n13172 = ~new_n13097 & ~new_n13171 ;
  assign new_n13173 = lo0873 & new_n13172 ;
  assign new_n13174 = ~lo0873 & ~new_n13172 ;
  assign new_n13175 = ~new_n13173 & ~new_n13174 ;
  assign new_n13176 = ~new_n13095 & new_n13175 ;
  assign new_n13177 = ~new_n2465 & ~new_n12441 ;
  assign new_n13178 = new_n12937 & new_n13177 ;
  assign new_n13179 = ~new_n2465 & ~new_n12442 ;
  assign new_n13180 = lo1292 & ~new_n12467 ;
  assign new_n13181 = ~lo1292 & ~new_n2465 ;
  assign new_n13182 = ~new_n13180 & ~new_n13181 ;
  assign new_n13183 = new_n2456 & ~new_n13182 ;
  assign new_n13184 = ~new_n2465 & new_n12965 ;
  assign new_n13185 = new_n12968 & ~new_n13182 ;
  assign new_n13186 = ~new_n12977 & new_n13185 ;
  assign new_n13187 = new_n12976 & ~new_n13185 ;
  assign new_n13188 = ~new_n2465 & new_n12429 ;
  assign new_n13189 = ~new_n2465 & new_n12602 ;
  assign new_n13190 = ~new_n2465 & new_n12441 ;
  assign new_n13191 = ~new_n13189 & ~new_n13190 ;
  assign new_n13192 = ~new_n12429 & ~new_n13191 ;
  assign new_n13193 = ~new_n13188 & ~new_n13192 ;
  assign new_n13194 = new_n12986 & ~new_n13193 ;
  assign new_n13195 = ~new_n13187 & ~new_n13194 ;
  assign new_n13196 = ~new_n13186 & new_n13195 ;
  assign new_n13197 = ~new_n12967 & ~new_n13196 ;
  assign new_n13198 = new_n12967 & new_n13196 ;
  assign new_n13199 = ~new_n13197 & ~new_n13198 ;
  assign new_n13200 = new_n13184 & ~new_n13199 ;
  assign new_n13201 = ~new_n13184 & new_n13197 ;
  assign new_n13202 = new_n12967 & new_n13189 ;
  assign new_n13203 = ~new_n13196 & new_n13202 ;
  assign new_n13204 = ~new_n13201 & ~new_n13203 ;
  assign new_n13205 = ~new_n13200 & new_n13204 ;
  assign new_n13206 = new_n12963 & ~new_n13205 ;
  assign new_n13207 = new_n12962 & ~new_n13206 ;
  assign new_n13208 = ~new_n12954 & ~new_n13207 ;
  assign new_n13209 = new_n12954 & new_n13207 ;
  assign new_n13210 = ~new_n13208 & ~new_n13209 ;
  assign new_n13211 = new_n13183 & ~new_n13210 ;
  assign new_n13212 = ~new_n13183 & new_n13208 ;
  assign new_n13213 = new_n13008 & ~new_n13207 ;
  assign new_n13214 = ~new_n13212 & ~new_n13213 ;
  assign new_n13215 = ~new_n13211 & new_n13214 ;
  assign new_n13216 = new_n12946 & new_n13215 ;
  assign new_n13217 = ~new_n13014 & ~new_n13215 ;
  assign new_n13218 = ~new_n2465 & ~new_n12329 ;
  assign new_n13219 = new_n13016 & new_n13218 ;
  assign new_n13220 = ~new_n13217 & ~new_n13219 ;
  assign new_n13221 = ~new_n13216 & new_n13220 ;
  assign new_n13222 = ~new_n12945 & ~new_n13221 ;
  assign new_n13223 = new_n12945 & new_n13221 ;
  assign new_n13224 = ~new_n13222 & ~new_n13223 ;
  assign new_n13225 = new_n13179 & ~new_n13224 ;
  assign new_n13226 = ~new_n13179 & new_n13222 ;
  assign new_n13227 = ~new_n12467 & new_n12945 ;
  assign new_n13228 = ~new_n13221 & new_n13227 ;
  assign new_n13229 = ~new_n13226 & ~new_n13228 ;
  assign new_n13230 = ~new_n13225 & new_n13229 ;
  assign new_n13231 = ~new_n2465 & ~new_n13064 ;
  assign new_n13232 = new_n13072 & new_n13231 ;
  assign new_n13233 = ~new_n13067 & new_n13231 ;
  assign new_n13234 = ~new_n13075 & ~new_n13233 ;
  assign new_n13235 = ~new_n13232 & new_n13234 ;
  assign new_n13236 = new_n13071 & ~new_n13235 ;
  assign new_n13237 = ~new_n13230 & new_n13236 ;
  assign new_n13238 = ~new_n13069 & ~new_n13235 ;
  assign new_n13239 = new_n13069 & new_n13235 ;
  assign new_n13240 = ~new_n13238 & ~new_n13239 ;
  assign new_n13241 = new_n13085 & ~new_n13240 ;
  assign new_n13242 = ~new_n13085 & new_n13238 ;
  assign new_n13243 = ~new_n13241 & ~new_n13242 ;
  assign new_n13244 = ~new_n13237 & new_n13243 ;
  assign new_n13245 = ~new_n12937 & ~new_n13244 ;
  assign new_n13246 = ~new_n13178 & ~new_n13245 ;
  assign new_n13247 = lo0875 & new_n13246 ;
  assign new_n13248 = ~new_n12452 & new_n12593 ;
  assign new_n13249 = new_n2456 & new_n12460 ;
  assign new_n13250 = ~new_n12441 & ~new_n13249 ;
  assign new_n13251 = ~new_n12467 & new_n12778 ;
  assign new_n13252 = ~new_n13250 & new_n13251 ;
  assign new_n13253 = ~new_n12550 & ~new_n13252 ;
  assign new_n13254 = new_n12452 & ~new_n13253 ;
  assign new_n13255 = ~new_n13248 & ~new_n13254 ;
  assign new_n13256 = new_n12508 & ~new_n13255 ;
  assign new_n13257 = ~new_n12467 & ~new_n12604 ;
  assign new_n13258 = new_n12467 & ~new_n12711 ;
  assign new_n13259 = ~new_n13257 & ~new_n13258 ;
  assign new_n13260 = new_n12420 & ~new_n13259 ;
  assign new_n13261 = ~new_n12512 & ~new_n13260 ;
  assign new_n13262 = new_n12452 & new_n12460 ;
  assign new_n13263 = lo0865 & new_n12964 ;
  assign new_n13264 = new_n12420 & ~new_n13263 ;
  assign new_n13265 = ~new_n12512 & ~new_n13264 ;
  assign new_n13266 = new_n13262 & ~new_n13265 ;
  assign new_n13267 = ~new_n12452 & ~new_n12460 ;
  assign new_n13268 = ~new_n12452 & new_n12460 ;
  assign new_n13269 = ~new_n12593 & ~new_n13264 ;
  assign new_n13270 = new_n13268 & ~new_n13269 ;
  assign new_n13271 = ~new_n13267 & ~new_n13270 ;
  assign new_n13272 = ~new_n13266 & new_n13271 ;
  assign new_n13273 = new_n12460 & ~new_n13272 ;
  assign new_n13274 = ~new_n12460 & new_n13272 ;
  assign new_n13275 = ~new_n13273 & ~new_n13274 ;
  assign new_n13276 = ~new_n13261 & ~new_n13275 ;
  assign new_n13277 = new_n13261 & new_n13273 ;
  assign new_n13278 = ~new_n12593 & ~new_n12605 ;
  assign new_n13279 = ~new_n12460 & ~new_n13278 ;
  assign new_n13280 = ~new_n13272 & new_n13279 ;
  assign new_n13281 = ~new_n13277 & ~new_n13280 ;
  assign new_n13282 = ~new_n13276 & new_n13281 ;
  assign new_n13283 = new_n2446 & ~new_n13282 ;
  assign new_n13284 = ~new_n2456 & new_n12325 ;
  assign new_n13285 = new_n12536 & ~new_n13284 ;
  assign new_n13286 = new_n2465 & new_n12367 ;
  assign new_n13287 = new_n12325 & ~new_n12357 ;
  assign new_n13288 = ~new_n13286 & new_n13287 ;
  assign new_n13289 = ~new_n13285 & ~new_n13288 ;
  assign new_n13290 = ~new_n2446 & ~new_n13289 ;
  assign new_n13291 = ~new_n13283 & ~new_n13290 ;
  assign new_n13292 = ~new_n12329 & ~new_n13291 ;
  assign new_n13293 = ~new_n13256 & ~new_n13292 ;
  assign new_n13294 = new_n2455 & ~new_n13293 ;
  assign new_n13295 = ~new_n12442 & new_n12517 ;
  assign new_n13296 = ~new_n12329 & ~new_n13295 ;
  assign new_n13297 = new_n12509 & ~new_n12524 ;
  assign new_n13298 = new_n12420 & ~new_n12442 ;
  assign new_n13299 = ~new_n12627 & ~new_n13298 ;
  assign new_n13300 = ~new_n12452 & ~new_n13299 ;
  assign new_n13301 = ~new_n13297 & ~new_n13300 ;
  assign new_n13302 = new_n12329 & ~new_n13301 ;
  assign new_n13303 = ~new_n13296 & ~new_n13302 ;
  assign new_n13304 = new_n2446 & ~new_n13303 ;
  assign new_n13305 = ~new_n12522 & ~new_n13304 ;
  assign new_n13306 = new_n2454 & ~new_n13305 ;
  assign new_n13307 = ~new_n2446 & new_n13085 ;
  assign new_n13308 = ~new_n12572 & ~new_n13307 ;
  assign new_n13309 = ~new_n2454 & ~new_n13308 ;
  assign new_n13310 = ~new_n13306 & ~new_n13309 ;
  assign new_n13311 = ~new_n2450 & ~new_n13310 ;
  assign new_n13312 = ~new_n13294 & ~new_n13311 ;
  assign new_n13313 = lo0872 & ~new_n13312 ;
  assign new_n13314 = ~new_n13247 & new_n13313 ;
  assign new_n13315 = ~new_n12325 & ~new_n12441 ;
  assign new_n13316 = new_n12937 & new_n13315 ;
  assign new_n13317 = ~new_n12325 & ~new_n12442 ;
  assign new_n13318 = lo0879 & ~new_n2265 ;
  assign new_n13319 = ~new_n2369 & ~new_n2442 ;
  assign new_n13320 = lo0880 & new_n2442 ;
  assign new_n13321 = ~new_n13319 & ~new_n13320 ;
  assign new_n13322 = ~new_n12454 & ~new_n13321 ;
  assign new_n13323 = new_n2265 & new_n13322 ;
  assign new_n13324 = ~new_n13318 & ~new_n13323 ;
  assign new_n13325 = lo1292 & ~new_n13324 ;
  assign new_n13326 = ~lo1292 & ~new_n12325 ;
  assign new_n13327 = ~new_n13325 & ~new_n13326 ;
  assign new_n13328 = new_n2456 & ~new_n13327 ;
  assign new_n13329 = ~new_n12325 & new_n12965 ;
  assign new_n13330 = new_n12968 & ~new_n13327 ;
  assign new_n13331 = ~new_n12977 & new_n13330 ;
  assign new_n13332 = new_n12976 & ~new_n13330 ;
  assign new_n13333 = ~new_n12325 & new_n12429 ;
  assign new_n13334 = ~new_n12325 & new_n12602 ;
  assign new_n13335 = ~new_n12325 & new_n12441 ;
  assign new_n13336 = ~new_n13334 & ~new_n13335 ;
  assign new_n13337 = ~new_n12429 & ~new_n13336 ;
  assign new_n13338 = ~new_n13333 & ~new_n13337 ;
  assign new_n13339 = new_n12986 & ~new_n13338 ;
  assign new_n13340 = ~new_n13332 & ~new_n13339 ;
  assign new_n13341 = ~new_n13331 & new_n13340 ;
  assign new_n13342 = ~new_n12967 & ~new_n13341 ;
  assign new_n13343 = new_n12967 & new_n13341 ;
  assign new_n13344 = ~new_n13342 & ~new_n13343 ;
  assign new_n13345 = new_n13329 & ~new_n13344 ;
  assign new_n13346 = ~new_n13329 & new_n13342 ;
  assign new_n13347 = new_n12967 & new_n13334 ;
  assign new_n13348 = ~new_n13341 & new_n13347 ;
  assign new_n13349 = ~new_n13346 & ~new_n13348 ;
  assign new_n13350 = ~new_n13345 & new_n13349 ;
  assign new_n13351 = new_n12963 & ~new_n13350 ;
  assign new_n13352 = new_n12962 & ~new_n13351 ;
  assign new_n13353 = ~new_n12954 & ~new_n13352 ;
  assign new_n13354 = new_n12954 & new_n13352 ;
  assign new_n13355 = ~new_n13353 & ~new_n13354 ;
  assign new_n13356 = new_n13328 & ~new_n13355 ;
  assign new_n13357 = ~new_n13328 & new_n13353 ;
  assign new_n13358 = new_n13008 & ~new_n13352 ;
  assign new_n13359 = ~new_n13357 & ~new_n13358 ;
  assign new_n13360 = ~new_n13356 & new_n13359 ;
  assign new_n13361 = new_n12946 & new_n13360 ;
  assign new_n13362 = ~new_n13014 & ~new_n13360 ;
  assign new_n13363 = new_n12337 & new_n13016 ;
  assign new_n13364 = ~new_n13362 & ~new_n13363 ;
  assign new_n13365 = ~new_n13361 & new_n13364 ;
  assign new_n13366 = ~new_n12945 & ~new_n13365 ;
  assign new_n13367 = new_n12945 & new_n13365 ;
  assign new_n13368 = ~new_n13366 & ~new_n13367 ;
  assign new_n13369 = new_n13317 & ~new_n13368 ;
  assign new_n13370 = ~new_n13317 & new_n13366 ;
  assign new_n13371 = new_n12945 & ~new_n13324 ;
  assign new_n13372 = ~new_n13365 & new_n13371 ;
  assign new_n13373 = ~new_n13370 & ~new_n13372 ;
  assign new_n13374 = ~new_n13369 & new_n13373 ;
  assign new_n13375 = ~new_n12325 & ~new_n13064 ;
  assign new_n13376 = new_n13072 & new_n13375 ;
  assign new_n13377 = ~new_n13067 & new_n13375 ;
  assign new_n13378 = ~new_n13075 & ~new_n13377 ;
  assign new_n13379 = ~new_n13376 & new_n13378 ;
  assign new_n13380 = new_n13071 & ~new_n13379 ;
  assign new_n13381 = ~new_n13374 & new_n13380 ;
  assign new_n13382 = ~new_n13069 & ~new_n13379 ;
  assign new_n13383 = new_n13069 & new_n13379 ;
  assign new_n13384 = ~new_n13382 & ~new_n13383 ;
  assign new_n13385 = new_n13085 & ~new_n13384 ;
  assign new_n13386 = ~new_n13085 & new_n13382 ;
  assign new_n13387 = ~new_n13385 & ~new_n13386 ;
  assign new_n13388 = ~new_n13381 & new_n13387 ;
  assign new_n13389 = ~new_n12937 & ~new_n13388 ;
  assign new_n13390 = ~new_n13316 & ~new_n13389 ;
  assign new_n13391 = lo0874 & new_n13390 ;
  assign new_n13392 = ~lo0874 & ~new_n13390 ;
  assign new_n13393 = ~new_n13391 & ~new_n13392 ;
  assign new_n13394 = lo0876 & new_n13094 ;
  assign new_n13395 = ~lo0875 & ~new_n13246 ;
  assign new_n13396 = ~new_n13394 & ~new_n13395 ;
  assign new_n13397 = new_n13393 & new_n13396 ;
  assign new_n13398 = new_n13314 & new_n13397 ;
  assign new_n13399 = new_n13176 & new_n13398 ;
  assign new_n13400 = new_n2450 & new_n13030 ;
  assign new_n13401 = new_n12553 & new_n12752 ;
  assign new_n13402 = ~new_n13400 & ~new_n13401 ;
  assign new_n13403 = new_n2446 & ~new_n12442 ;
  assign new_n13404 = new_n2454 & new_n13403 ;
  assign new_n13405 = ~new_n13402 & new_n13404 ;
  assign new_n13406 = ~new_n2454 & ~new_n12329 ;
  assign new_n13407 = new_n2446 & new_n13406 ;
  assign new_n13408 = new_n12590 & new_n12591 ;
  assign new_n13409 = new_n2454 & new_n13408 ;
  assign new_n13410 = ~new_n13407 & ~new_n13409 ;
  assign new_n13411 = new_n2450 & ~new_n13410 ;
  assign new_n13412 = ~new_n13405 & ~new_n13411 ;
  assign new_n13413 = ~new_n13324 & ~new_n13412 ;
  assign new_n13414 = new_n12329 & new_n12420 ;
  assign new_n13415 = new_n12951 & new_n13414 ;
  assign new_n13416 = ~new_n12329 & new_n12429 ;
  assign new_n13417 = ~new_n12460 & new_n13416 ;
  assign new_n13418 = new_n12510 & new_n13417 ;
  assign new_n13419 = ~new_n13415 & ~new_n13418 ;
  assign new_n13420 = new_n2450 & ~new_n13419 ;
  assign new_n13421 = new_n12452 & new_n12549 ;
  assign new_n13422 = new_n12698 & new_n13421 ;
  assign new_n13423 = ~new_n2454 & ~new_n13422 ;
  assign new_n13424 = new_n2454 & new_n12698 ;
  assign new_n13425 = ~new_n13423 & ~new_n13424 ;
  assign new_n13426 = ~new_n13420 & new_n13425 ;
  assign new_n13427 = new_n2446 & ~new_n13426 ;
  assign new_n13428 = ~new_n12325 & new_n13427 ;
  assign new_n13429 = new_n2446 & new_n2450 ;
  assign new_n13430 = lo1291 & lo1293 ;
  assign new_n13431 = lo1291 & ~new_n13430 ;
  assign new_n13432 = lo1292 & ~lo1294 ;
  assign new_n13433 = ~new_n13431 & new_n13432 ;
  assign new_n13434 = new_n12573 & new_n13433 ;
  assign new_n13435 = ~new_n13082 & ~new_n13434 ;
  assign new_n13436 = new_n13406 & ~new_n13435 ;
  assign new_n13437 = new_n2446 & new_n12951 ;
  assign new_n13438 = new_n2450 & ~new_n13437 ;
  assign new_n13439 = new_n2446 & new_n13438 ;
  assign new_n13440 = ~new_n13436 & new_n13439 ;
  assign new_n13441 = ~new_n2446 & ~new_n13438 ;
  assign new_n13442 = ~new_n13439 & ~new_n13441 ;
  assign new_n13443 = new_n13436 & ~new_n13442 ;
  assign new_n13444 = new_n12800 & new_n13438 ;
  assign new_n13445 = new_n12956 & new_n13444 ;
  assign new_n13446 = ~new_n13443 & ~new_n13445 ;
  assign new_n13447 = ~new_n13440 & new_n13446 ;
  assign new_n13448 = new_n13429 & ~new_n13447 ;
  assign new_n13449 = new_n12420 & ~new_n12467 ;
  assign new_n13450 = ~new_n12720 & ~new_n13449 ;
  assign new_n13451 = ~new_n12420 & ~new_n13450 ;
  assign new_n13452 = new_n12420 & new_n13450 ;
  assign new_n13453 = ~new_n13451 & ~new_n13452 ;
  assign new_n13454 = new_n13334 & ~new_n13453 ;
  assign new_n13455 = ~new_n13334 & new_n13451 ;
  assign new_n13456 = ~new_n12420 & new_n13334 ;
  assign new_n13457 = new_n13334 & ~new_n13456 ;
  assign new_n13458 = new_n13335 & new_n13450 ;
  assign new_n13459 = ~new_n13457 & new_n13458 ;
  assign new_n13460 = ~new_n13455 & ~new_n13459 ;
  assign new_n13461 = ~new_n13454 & new_n13460 ;
  assign new_n13462 = new_n13450 & ~new_n13461 ;
  assign new_n13463 = ~new_n13450 & new_n13461 ;
  assign new_n13464 = ~new_n13462 & ~new_n13463 ;
  assign new_n13465 = new_n13329 & ~new_n13464 ;
  assign new_n13466 = ~new_n13329 & new_n13462 ;
  assign new_n13467 = new_n13330 & ~new_n13450 ;
  assign new_n13468 = ~new_n13461 & new_n13467 ;
  assign new_n13469 = ~new_n13466 & ~new_n13468 ;
  assign new_n13470 = ~new_n13465 & new_n13469 ;
  assign new_n13471 = ~new_n12452 & new_n12523 ;
  assign new_n13472 = new_n12420 & ~new_n13471 ;
  assign new_n13473 = new_n12429 & ~new_n12509 ;
  assign new_n13474 = ~new_n13472 & new_n13473 ;
  assign new_n13475 = ~new_n12329 & ~new_n13474 ;
  assign new_n13476 = ~new_n12329 & ~new_n13475 ;
  assign new_n13477 = new_n12460 & ~new_n12720 ;
  assign new_n13478 = ~new_n12606 & ~new_n13477 ;
  assign new_n13479 = new_n13475 & ~new_n13478 ;
  assign new_n13480 = ~new_n13476 & ~new_n13479 ;
  assign new_n13481 = new_n13475 & ~new_n13480 ;
  assign new_n13482 = new_n12594 & ~new_n13475 ;
  assign new_n13483 = new_n13480 & new_n13482 ;
  assign new_n13484 = ~new_n13481 & ~new_n13483 ;
  assign new_n13485 = new_n13315 & ~new_n13475 ;
  assign new_n13486 = ~new_n13480 & new_n13485 ;
  assign new_n13487 = new_n13484 & ~new_n13486 ;
  assign new_n13488 = ~new_n13475 & ~new_n13487 ;
  assign new_n13489 = new_n13475 & new_n13487 ;
  assign new_n13490 = ~new_n13488 & ~new_n13489 ;
  assign new_n13491 = ~new_n13470 & ~new_n13490 ;
  assign new_n13492 = new_n13470 & new_n13488 ;
  assign new_n13493 = ~new_n13338 & new_n13475 ;
  assign new_n13494 = ~new_n13487 & new_n13493 ;
  assign new_n13495 = ~new_n13492 & ~new_n13494 ;
  assign new_n13496 = ~new_n13491 & new_n13495 ;
  assign new_n13497 = new_n13448 & ~new_n13496 ;
  assign new_n13498 = ~new_n13429 & ~new_n13447 ;
  assign new_n13499 = new_n13429 & new_n13447 ;
  assign new_n13500 = ~new_n13498 & ~new_n13499 ;
  assign new_n13501 = new_n13328 & ~new_n13500 ;
  assign new_n13502 = ~new_n13328 & new_n13498 ;
  assign new_n13503 = ~new_n13501 & ~new_n13502 ;
  assign new_n13504 = ~new_n13497 & new_n13503 ;
  assign new_n13505 = ~new_n13427 & ~new_n13504 ;
  assign new_n13506 = ~new_n13428 & ~new_n13505 ;
  assign new_n13507 = new_n13412 & ~new_n13506 ;
  assign new_n13508 = ~new_n13413 & ~new_n13507 ;
  assign new_n13509 = ~lo0874 & ~new_n13508 ;
  assign new_n13510 = ~new_n2454 & ~new_n13421 ;
  assign new_n13511 = new_n2454 & new_n13053 ;
  assign new_n13512 = ~new_n2454 & new_n12329 ;
  assign new_n13513 = ~new_n12709 & ~new_n13512 ;
  assign new_n13514 = ~new_n13511 & ~new_n13513 ;
  assign new_n13515 = ~new_n13510 & new_n13514 ;
  assign new_n13516 = new_n12467 & ~new_n13263 ;
  assign new_n13517 = ~new_n12420 & ~new_n12442 ;
  assign new_n13518 = ~new_n12605 & ~new_n13517 ;
  assign new_n13519 = ~new_n12467 & ~new_n13518 ;
  assign new_n13520 = ~new_n13516 & ~new_n13519 ;
  assign new_n13521 = ~new_n12429 & new_n12968 ;
  assign new_n13522 = ~new_n12550 & ~new_n13521 ;
  assign new_n13523 = ~new_n12420 & ~new_n13522 ;
  assign new_n13524 = ~new_n13264 & ~new_n13523 ;
  assign new_n13525 = new_n13268 & ~new_n13524 ;
  assign new_n13526 = new_n13262 & ~new_n13263 ;
  assign new_n13527 = ~new_n13267 & ~new_n13526 ;
  assign new_n13528 = ~new_n13525 & new_n13527 ;
  assign new_n13529 = new_n12460 & ~new_n13528 ;
  assign new_n13530 = ~new_n12460 & new_n13528 ;
  assign new_n13531 = ~new_n13529 & ~new_n13530 ;
  assign new_n13532 = ~new_n13520 & ~new_n13531 ;
  assign new_n13533 = new_n13520 & new_n13529 ;
  assign new_n13534 = ~new_n12420 & new_n12968 ;
  assign new_n13535 = ~new_n12467 & new_n12602 ;
  assign new_n13536 = lo0865 & ~new_n2264 ;
  assign new_n13537 = new_n12467 & ~new_n13536 ;
  assign new_n13538 = ~new_n13535 & ~new_n13537 ;
  assign new_n13539 = new_n12420 & ~new_n13538 ;
  assign new_n13540 = ~new_n13534 & ~new_n13539 ;
  assign new_n13541 = ~new_n12429 & ~new_n13540 ;
  assign new_n13542 = ~new_n12550 & ~new_n13541 ;
  assign new_n13543 = ~new_n12460 & ~new_n13542 ;
  assign new_n13544 = ~new_n13528 & new_n13543 ;
  assign new_n13545 = ~new_n13533 & ~new_n13544 ;
  assign new_n13546 = ~new_n13532 & new_n13545 ;
  assign new_n13547 = ~new_n12329 & ~new_n13546 ;
  assign new_n13548 = ~new_n2456 & new_n12443 ;
  assign new_n13549 = ~new_n12452 & ~new_n13548 ;
  assign new_n13550 = ~new_n12595 & ~new_n13549 ;
  assign new_n13551 = new_n12329 & ~new_n13550 ;
  assign new_n13552 = new_n2454 & ~new_n13551 ;
  assign new_n13553 = ~new_n13547 & new_n13552 ;
  assign new_n13554 = new_n13429 & ~new_n13553 ;
  assign new_n13555 = ~new_n12329 & new_n12678 ;
  assign new_n13556 = new_n12370 & new_n13286 ;
  assign new_n13557 = new_n2465 & new_n12373 ;
  assign new_n13558 = new_n2465 & new_n12329 ;
  assign new_n13559 = ~new_n13557 & new_n13558 ;
  assign new_n13560 = ~new_n13556 & new_n13559 ;
  assign new_n13561 = ~new_n13555 & ~new_n13560 ;
  assign new_n13562 = ~new_n2446 & new_n2455 ;
  assign new_n13563 = ~new_n13561 & new_n13562 ;
  assign new_n13564 = ~new_n13065 & ~new_n13563 ;
  assign new_n13565 = ~new_n13554 & new_n13564 ;
  assign new_n13566 = new_n2450 & ~new_n13565 ;
  assign new_n13567 = ~new_n2450 & new_n13565 ;
  assign new_n13568 = ~new_n13566 & ~new_n13567 ;
  assign new_n13569 = ~new_n13515 & ~new_n13568 ;
  assign new_n13570 = new_n13515 & new_n13566 ;
  assign new_n13571 = ~new_n2450 & new_n13436 ;
  assign new_n13572 = ~new_n13565 & new_n13571 ;
  assign new_n13573 = ~new_n13570 & ~new_n13572 ;
  assign new_n13574 = ~new_n13569 & new_n13573 ;
  assign new_n13575 = lo0872 & ~new_n13574 ;
  assign new_n13576 = ~new_n13509 & new_n13575 ;
  assign new_n13577 = lo0874 & new_n13508 ;
  assign new_n13578 = ~new_n12460 & ~new_n13412 ;
  assign new_n13579 = ~new_n12367 & new_n13427 ;
  assign new_n13580 = new_n12981 & ~new_n13453 ;
  assign new_n13581 = ~new_n12981 & new_n13451 ;
  assign new_n13582 = ~new_n12420 & new_n12981 ;
  assign new_n13583 = new_n12981 & ~new_n13582 ;
  assign new_n13584 = new_n12982 & new_n13450 ;
  assign new_n13585 = ~new_n13583 & new_n13584 ;
  assign new_n13586 = ~new_n13581 & ~new_n13585 ;
  assign new_n13587 = ~new_n13580 & new_n13586 ;
  assign new_n13588 = new_n13450 & ~new_n13587 ;
  assign new_n13589 = ~new_n13450 & new_n13587 ;
  assign new_n13590 = ~new_n13588 & ~new_n13589 ;
  assign new_n13591 = new_n12966 & ~new_n13590 ;
  assign new_n13592 = ~new_n12966 & new_n13588 ;
  assign new_n13593 = new_n12969 & ~new_n13450 ;
  assign new_n13594 = ~new_n13587 & new_n13593 ;
  assign new_n13595 = ~new_n13592 & ~new_n13594 ;
  assign new_n13596 = ~new_n13591 & new_n13595 ;
  assign new_n13597 = new_n12931 & ~new_n13475 ;
  assign new_n13598 = ~new_n13480 & new_n13597 ;
  assign new_n13599 = new_n13484 & ~new_n13598 ;
  assign new_n13600 = ~new_n13475 & ~new_n13599 ;
  assign new_n13601 = new_n13475 & new_n13599 ;
  assign new_n13602 = ~new_n13600 & ~new_n13601 ;
  assign new_n13603 = ~new_n13596 & ~new_n13602 ;
  assign new_n13604 = new_n13596 & new_n13600 ;
  assign new_n13605 = ~new_n12985 & new_n13475 ;
  assign new_n13606 = ~new_n13599 & new_n13605 ;
  assign new_n13607 = ~new_n13604 & ~new_n13606 ;
  assign new_n13608 = ~new_n13603 & new_n13607 ;
  assign new_n13609 = new_n13448 & ~new_n13608 ;
  assign new_n13610 = new_n12950 & ~new_n13500 ;
  assign new_n13611 = ~new_n12950 & new_n13498 ;
  assign new_n13612 = ~new_n13610 & ~new_n13611 ;
  assign new_n13613 = ~new_n13609 & new_n13612 ;
  assign new_n13614 = ~new_n13427 & ~new_n13613 ;
  assign new_n13615 = ~new_n13579 & ~new_n13614 ;
  assign new_n13616 = new_n13412 & ~new_n13615 ;
  assign new_n13617 = ~new_n13578 & ~new_n13616 ;
  assign new_n13618 = lo0876 & new_n13617 ;
  assign new_n13619 = ~lo0876 & ~new_n13617 ;
  assign new_n13620 = ~new_n13618 & ~new_n13619 ;
  assign new_n13621 = ~new_n13577 & new_n13620 ;
  assign new_n13622 = new_n13576 & new_n13621 ;
  assign new_n13623 = ~new_n12467 & ~new_n13412 ;
  assign new_n13624 = ~new_n2465 & new_n13427 ;
  assign new_n13625 = new_n13189 & ~new_n13453 ;
  assign new_n13626 = ~new_n13189 & new_n13451 ;
  assign new_n13627 = ~new_n12420 & new_n13189 ;
  assign new_n13628 = new_n13189 & ~new_n13627 ;
  assign new_n13629 = new_n13190 & new_n13450 ;
  assign new_n13630 = ~new_n13628 & new_n13629 ;
  assign new_n13631 = ~new_n13626 & ~new_n13630 ;
  assign new_n13632 = ~new_n13625 & new_n13631 ;
  assign new_n13633 = new_n13450 & ~new_n13632 ;
  assign new_n13634 = ~new_n13450 & new_n13632 ;
  assign new_n13635 = ~new_n13633 & ~new_n13634 ;
  assign new_n13636 = new_n13184 & ~new_n13635 ;
  assign new_n13637 = ~new_n13184 & new_n13633 ;
  assign new_n13638 = new_n13185 & ~new_n13450 ;
  assign new_n13639 = ~new_n13632 & new_n13638 ;
  assign new_n13640 = ~new_n13637 & ~new_n13639 ;
  assign new_n13641 = ~new_n13636 & new_n13640 ;
  assign new_n13642 = new_n13475 & new_n13480 ;
  assign new_n13643 = ~new_n13641 & new_n13642 ;
  assign new_n13644 = new_n13484 & ~new_n13643 ;
  assign new_n13645 = new_n13480 & ~new_n13644 ;
  assign new_n13646 = ~new_n13480 & new_n13644 ;
  assign new_n13647 = ~new_n13645 & ~new_n13646 ;
  assign new_n13648 = new_n13177 & ~new_n13647 ;
  assign new_n13649 = ~new_n13177 & new_n13645 ;
  assign new_n13650 = ~new_n13193 & ~new_n13480 ;
  assign new_n13651 = ~new_n13644 & new_n13650 ;
  assign new_n13652 = ~new_n13649 & ~new_n13651 ;
  assign new_n13653 = ~new_n13648 & new_n13652 ;
  assign new_n13654 = new_n13448 & ~new_n13653 ;
  assign new_n13655 = new_n13183 & ~new_n13500 ;
  assign new_n13656 = ~new_n13183 & new_n13498 ;
  assign new_n13657 = ~new_n13655 & ~new_n13656 ;
  assign new_n13658 = ~new_n13654 & new_n13657 ;
  assign new_n13659 = ~new_n13427 & ~new_n13658 ;
  assign new_n13660 = ~new_n13624 & ~new_n13659 ;
  assign new_n13661 = new_n13412 & ~new_n13660 ;
  assign new_n13662 = ~new_n13623 & ~new_n13661 ;
  assign new_n13663 = lo0875 & new_n13662 ;
  assign new_n13664 = ~new_n13105 & ~new_n13412 ;
  assign new_n13665 = ~new_n12357 & new_n13427 ;
  assign new_n13666 = new_n13115 & ~new_n13453 ;
  assign new_n13667 = ~new_n13115 & new_n13451 ;
  assign new_n13668 = ~new_n12420 & new_n13115 ;
  assign new_n13669 = new_n13115 & ~new_n13668 ;
  assign new_n13670 = new_n13116 & new_n13450 ;
  assign new_n13671 = ~new_n13669 & new_n13670 ;
  assign new_n13672 = ~new_n13667 & ~new_n13671 ;
  assign new_n13673 = ~new_n13666 & new_n13672 ;
  assign new_n13674 = new_n13450 & ~new_n13673 ;
  assign new_n13675 = ~new_n13450 & new_n13673 ;
  assign new_n13676 = ~new_n13674 & ~new_n13675 ;
  assign new_n13677 = new_n13110 & ~new_n13676 ;
  assign new_n13678 = ~new_n13110 & new_n13674 ;
  assign new_n13679 = new_n13111 & ~new_n13450 ;
  assign new_n13680 = ~new_n13673 & new_n13679 ;
  assign new_n13681 = ~new_n13678 & ~new_n13680 ;
  assign new_n13682 = ~new_n13677 & new_n13681 ;
  assign new_n13683 = new_n13642 & ~new_n13682 ;
  assign new_n13684 = new_n13484 & ~new_n13683 ;
  assign new_n13685 = new_n13480 & ~new_n13684 ;
  assign new_n13686 = ~new_n13480 & new_n13684 ;
  assign new_n13687 = ~new_n13685 & ~new_n13686 ;
  assign new_n13688 = new_n13096 & ~new_n13687 ;
  assign new_n13689 = ~new_n13096 & new_n13685 ;
  assign new_n13690 = ~new_n13119 & ~new_n13480 ;
  assign new_n13691 = ~new_n13684 & new_n13690 ;
  assign new_n13692 = ~new_n13689 & ~new_n13691 ;
  assign new_n13693 = ~new_n13688 & new_n13692 ;
  assign new_n13694 = new_n13448 & ~new_n13693 ;
  assign new_n13695 = new_n13109 & ~new_n13500 ;
  assign new_n13696 = ~new_n13109 & new_n13498 ;
  assign new_n13697 = ~new_n13695 & ~new_n13696 ;
  assign new_n13698 = ~new_n13694 & new_n13697 ;
  assign new_n13699 = ~new_n13427 & ~new_n13698 ;
  assign new_n13700 = ~new_n13665 & ~new_n13699 ;
  assign new_n13701 = new_n13412 & ~new_n13700 ;
  assign new_n13702 = ~new_n13664 & ~new_n13701 ;
  assign new_n13703 = ~lo0873 & ~new_n13702 ;
  assign new_n13704 = ~new_n13663 & ~new_n13703 ;
  assign new_n13705 = ~lo0875 & ~new_n13662 ;
  assign new_n13706 = lo0873 & new_n13702 ;
  assign new_n13707 = ~new_n13705 & ~new_n13706 ;
  assign new_n13708 = new_n13704 & new_n13707 ;
  assign new_n13709 = new_n13622 & new_n13708 ;
  assign new_n13710 = new_n12405 & ~new_n13053 ;
  assign new_n13711 = ~new_n2454 & new_n13421 ;
  assign new_n13712 = ~new_n2450 & ~new_n13711 ;
  assign new_n13713 = new_n2454 & new_n12553 ;
  assign new_n13714 = ~new_n12404 & ~new_n13713 ;
  assign new_n13715 = ~new_n13712 & new_n13714 ;
  assign new_n13716 = new_n12329 & ~new_n13715 ;
  assign new_n13717 = ~new_n13710 & ~new_n13716 ;
  assign new_n13718 = ~new_n13324 & ~new_n13717 ;
  assign new_n13719 = new_n2455 & new_n12603 ;
  assign new_n13720 = new_n13414 & new_n13719 ;
  assign new_n13721 = new_n13717 & new_n13720 ;
  assign new_n13722 = ~new_n12325 & new_n13721 ;
  assign new_n13723 = ~new_n13718 & ~new_n13722 ;
  assign new_n13724 = new_n2446 & ~new_n13723 ;
  assign new_n13725 = lo0874 & ~new_n13724 ;
  assign new_n13726 = ~lo0874 & new_n13724 ;
  assign new_n13727 = ~new_n13725 & ~new_n13726 ;
  assign new_n13728 = ~new_n12460 & ~new_n13717 ;
  assign new_n13729 = ~new_n12367 & new_n13721 ;
  assign new_n13730 = ~new_n13728 & ~new_n13729 ;
  assign new_n13731 = new_n2446 & ~new_n13730 ;
  assign new_n13732 = ~lo0876 & new_n13731 ;
  assign new_n13733 = ~new_n13105 & ~new_n13717 ;
  assign new_n13734 = ~new_n12357 & new_n13721 ;
  assign new_n13735 = ~new_n13733 & ~new_n13734 ;
  assign new_n13736 = new_n2446 & ~new_n13735 ;
  assign new_n13737 = ~lo0873 & new_n13736 ;
  assign new_n13738 = ~new_n13732 & ~new_n13737 ;
  assign new_n13739 = new_n13727 & new_n13738 ;
  assign new_n13740 = new_n12329 & ~new_n12467 ;
  assign new_n13741 = ~new_n12329 & ~new_n12467 ;
  assign new_n13742 = ~new_n13053 & new_n13741 ;
  assign new_n13743 = ~new_n13740 & ~new_n13742 ;
  assign new_n13744 = ~new_n12452 & ~new_n12467 ;
  assign new_n13745 = ~new_n2465 & new_n12452 ;
  assign new_n13746 = new_n12603 & new_n13745 ;
  assign new_n13747 = ~new_n13744 & ~new_n13746 ;
  assign new_n13748 = new_n2455 & new_n13414 ;
  assign new_n13749 = ~new_n13747 & new_n13748 ;
  assign new_n13750 = new_n12404 & new_n13740 ;
  assign new_n13751 = ~new_n12402 & ~new_n13750 ;
  assign new_n13752 = ~new_n13749 & new_n13751 ;
  assign new_n13753 = new_n2450 & ~new_n13752 ;
  assign new_n13754 = ~new_n2450 & new_n13752 ;
  assign new_n13755 = ~new_n13753 & ~new_n13754 ;
  assign new_n13756 = ~new_n13743 & ~new_n13755 ;
  assign new_n13757 = new_n13743 & new_n13753 ;
  assign new_n13758 = ~new_n2450 & new_n13740 ;
  assign new_n13759 = ~new_n13421 & new_n13758 ;
  assign new_n13760 = ~new_n13752 & new_n13759 ;
  assign new_n13761 = ~new_n13757 & ~new_n13760 ;
  assign new_n13762 = ~new_n13756 & new_n13761 ;
  assign new_n13763 = new_n2446 & ~new_n13762 ;
  assign new_n13764 = ~lo0875 & new_n13763 ;
  assign new_n13765 = lo0875 & ~new_n13763 ;
  assign new_n13766 = new_n12698 & ~new_n13421 ;
  assign new_n13767 = ~new_n2450 & ~new_n13053 ;
  assign new_n13768 = new_n12517 & new_n12761 ;
  assign new_n13769 = ~new_n12553 & ~new_n13768 ;
  assign new_n13770 = new_n12329 & ~new_n13769 ;
  assign new_n13771 = ~new_n13767 & ~new_n13770 ;
  assign new_n13772 = new_n2454 & ~new_n13771 ;
  assign new_n13773 = ~new_n13766 & ~new_n13772 ;
  assign new_n13774 = new_n2446 & ~new_n13773 ;
  assign new_n13775 = ~new_n2454 & new_n12508 ;
  assign new_n13776 = new_n2465 & new_n12358 ;
  assign new_n13777 = new_n12329 & new_n13776 ;
  assign new_n13778 = new_n12325 & ~new_n12368 ;
  assign new_n13779 = new_n2264 & ~new_n12325 ;
  assign new_n13780 = ~new_n13778 & ~new_n13779 ;
  assign new_n13781 = ~new_n12325 & new_n12357 ;
  assign new_n13782 = ~new_n13287 & ~new_n13781 ;
  assign new_n13783 = ~new_n12329 & new_n13782 ;
  assign new_n13784 = ~new_n13780 & new_n13783 ;
  assign new_n13785 = ~new_n13777 & ~new_n13784 ;
  assign new_n13786 = new_n12800 & ~new_n13785 ;
  assign new_n13787 = ~new_n13775 & ~new_n13786 ;
  assign new_n13788 = new_n2450 & ~new_n13787 ;
  assign new_n13789 = ~new_n13774 & ~new_n13788 ;
  assign new_n13790 = lo0872 & ~new_n13789 ;
  assign new_n13791 = ~new_n13765 & new_n13790 ;
  assign new_n13792 = ~new_n13764 & new_n13791 ;
  assign new_n13793 = lo0876 & ~new_n13731 ;
  assign new_n13794 = lo0873 & ~new_n13736 ;
  assign new_n13795 = ~new_n13793 & ~new_n13794 ;
  assign new_n13796 = new_n13792 & new_n13795 ;
  assign new_n13797 = new_n13739 & new_n13796 ;
  assign new_n13798 = new_n12517 & new_n12550 ;
  assign new_n13799 = new_n13741 & new_n13798 ;
  assign new_n13800 = new_n2264 & ~new_n12429 ;
  assign new_n13801 = new_n12468 & new_n13800 ;
  assign new_n13802 = new_n12429 & ~new_n12467 ;
  assign new_n13803 = ~new_n13801 & ~new_n13802 ;
  assign new_n13804 = ~new_n12441 & new_n13046 ;
  assign new_n13805 = ~new_n13803 & new_n13804 ;
  assign new_n13806 = ~new_n13799 & ~new_n13805 ;
  assign new_n13807 = new_n2446 & new_n2455 ;
  assign new_n13808 = ~new_n13806 & new_n13807 ;
  assign new_n13809 = ~new_n12329 & new_n13807 ;
  assign new_n13810 = new_n12509 & new_n12550 ;
  assign new_n13811 = ~new_n12467 & new_n13810 ;
  assign new_n13812 = new_n13809 & new_n13811 ;
  assign new_n13813 = ~new_n13808 & ~new_n13812 ;
  assign new_n13814 = lo0881 & ~new_n13813 ;
  assign new_n13815 = ~new_n13797 & ~new_n13814 ;
  assign new_n13816 = ~new_n13709 & new_n13815 ;
  assign new_n13817 = ~new_n13399 & new_n13816 ;
  assign new_n13818 = ~new_n12930 & new_n13817 ;
  assign new_n13819 = ~new_n12420 & ~new_n12441 ;
  assign new_n13820 = new_n2454 & new_n13819 ;
  assign new_n13821 = ~new_n2454 & new_n12549 ;
  assign new_n13822 = ~new_n13820 & ~new_n13821 ;
  assign new_n13823 = ~new_n2450 & ~new_n12452 ;
  assign new_n13824 = ~new_n13822 & new_n13823 ;
  assign new_n13825 = new_n12329 & new_n13824 ;
  assign new_n13826 = new_n12467 & new_n12550 ;
  assign new_n13827 = ~new_n12329 & ~new_n12720 ;
  assign new_n13828 = new_n13826 & new_n13827 ;
  assign new_n13829 = new_n12442 & ~new_n12452 ;
  assign new_n13830 = ~new_n12441 & new_n12467 ;
  assign new_n13831 = ~new_n13047 & ~new_n13830 ;
  assign new_n13832 = new_n12933 & ~new_n13831 ;
  assign new_n13833 = ~new_n13829 & ~new_n13832 ;
  assign new_n13834 = ~new_n12509 & ~new_n12553 ;
  assign new_n13835 = new_n12329 & ~new_n13834 ;
  assign new_n13836 = ~new_n13833 & new_n13835 ;
  assign new_n13837 = ~new_n13828 & ~new_n13836 ;
  assign new_n13838 = new_n2455 & ~new_n13837 ;
  assign new_n13839 = ~new_n13825 & ~new_n13838 ;
  assign new_n13840 = ~lo0888 & ~lo0889 ;
  assign new_n13841 = ~lo0887 & new_n13840 ;
  assign new_n13842 = new_n2020 & new_n13841 ;
  assign new_n13843 = ~lo0885 & ~lo0886 ;
  assign new_n13844 = ~lo0883 & ~lo0884 ;
  assign new_n13845 = ~lo0882 & new_n13844 ;
  assign new_n13846 = new_n13843 & new_n13845 ;
  assign new_n13847 = new_n13842 & new_n13846 ;
  assign new_n13848 = new_n2446 & ~new_n13847 ;
  assign new_n13849 = ~new_n13839 & new_n13848 ;
  assign new_n13850 = new_n13818 & ~new_n13849 ;
  assign new_n13851 = ~new_n12505 & new_n13850 ;
  assign new_n13852 = ~new_n2254 & new_n13851 ;
  assign new_n13853 = lo0118 & ~new_n2249 ;
  assign new_n13854 = lo0117 & lo0119 ;
  assign new_n13855 = ~new_n13853 & new_n13854 ;
  assign new_n13856 = ~lo0117 & ~lo0118 ;
  assign new_n13857 = new_n2249 & new_n13856 ;
  assign new_n13858 = ~new_n2257 & new_n13857 ;
  assign new_n13859 = ~new_n13855 & ~new_n13858 ;
  assign new_n13860 = ~new_n13852 & new_n13859 ;
  assign new_n13861 = new_n12383 & ~new_n12655 ;
  assign new_n13862 = ~new_n2446 & new_n12910 ;
  assign new_n13863 = new_n12420 & new_n12442 ;
  assign new_n13864 = ~new_n12778 & ~new_n13863 ;
  assign new_n13865 = new_n12383 & new_n12420 ;
  assign new_n13866 = new_n12383 & new_n12467 ;
  assign new_n13867 = ~new_n12467 & new_n12473 ;
  assign new_n13868 = ~new_n13866 & ~new_n13867 ;
  assign new_n13869 = ~new_n12441 & new_n12460 ;
  assign new_n13870 = ~new_n13868 & new_n13869 ;
  assign new_n13871 = ~new_n13865 & ~new_n13870 ;
  assign new_n13872 = ~new_n13864 & ~new_n13871 ;
  assign new_n13873 = new_n2446 & new_n13872 ;
  assign new_n13874 = ~new_n13862 & ~new_n13873 ;
  assign new_n13875 = new_n12655 & ~new_n13874 ;
  assign new_n13876 = ~new_n13861 & ~new_n13875 ;
  assign new_n13877 = new_n12443 & new_n12460 ;
  assign new_n13878 = ~new_n12329 & ~new_n13877 ;
  assign new_n13879 = new_n2446 & new_n12452 ;
  assign new_n13880 = ~new_n13878 & new_n13879 ;
  assign new_n13881 = ~new_n12374 & ~new_n12955 ;
  assign new_n13882 = ~new_n2446 & ~new_n13881 ;
  assign new_n13883 = ~new_n13880 & ~new_n13882 ;
  assign new_n13884 = new_n2455 & ~new_n13883 ;
  assign new_n13885 = ~new_n13876 & new_n13884 ;
  assign new_n13886 = ~new_n12386 & new_n12916 ;
  assign new_n13887 = new_n12395 & new_n12910 ;
  assign new_n13888 = lo1291 & new_n12909 ;
  assign new_n13889 = new_n12325 & new_n13888 ;
  assign new_n13890 = ~new_n13887 & ~new_n13889 ;
  assign new_n13891 = new_n12357 & ~new_n13890 ;
  assign new_n13892 = ~new_n13886 & ~new_n13891 ;
  assign new_n13893 = ~new_n12329 & ~new_n13892 ;
  assign new_n13894 = ~new_n12384 & ~new_n13893 ;
  assign new_n13895 = new_n12789 & ~new_n13894 ;
  assign new_n13896 = new_n12383 & new_n12590 ;
  assign new_n13897 = new_n2454 & new_n13896 ;
  assign new_n13898 = ~new_n13895 & ~new_n13897 ;
  assign new_n13899 = ~new_n2450 & ~new_n13898 ;
  assign new_n13900 = ~new_n13885 & ~new_n13899 ;
  assign new_n13901 = new_n13818 & ~new_n13900 ;
  assign new_n13902 = lo0954 & new_n11741 ;
  assign new_n13903 = new_n11741 & ~new_n13902 ;
  assign new_n13904 = ~new_n9180 & ~new_n13903 ;
  assign new_n13905 = ~lo0954 & new_n9180 ;
  assign new_n13906 = ~new_n11741 & new_n13905 ;
  assign new_n13907 = ~new_n13904 & ~new_n13906 ;
  assign new_n13908 = ~new_n13900 & ~new_n13907 ;
  assign new_n13909 = ~lo0803 & new_n13900 ;
  assign new_n13910 = ~new_n13908 & ~new_n13909 ;
  assign new_n13911 = ~new_n13901 & ~new_n13910 ;
  assign new_n13912 = ~lo0120 & new_n13851 ;
  assign new_n13913 = ~new_n13911 & new_n13912 ;
  assign new_n13914 = lo0119 & ~lo0893 ;
  assign new_n13915 = ~lo0037 & new_n13914 ;
  assign new_n13916 = new_n13856 & new_n13915 ;
  assign new_n13917 = ~lo0892 & ~new_n2249 ;
  assign new_n13918 = new_n13916 & new_n13917 ;
  assign new_n13919 = ~new_n13913 & new_n13918 ;
  assign new_n13920 = new_n2256 & new_n13911 ;
  assign new_n13921 = new_n2256 & ~new_n13851 ;
  assign new_n13922 = lo0118 & new_n2254 ;
  assign new_n13923 = ~new_n13921 & ~new_n13922 ;
  assign new_n13924 = ~new_n13920 & new_n13923 ;
  assign new_n13925 = ~new_n13919 & new_n13924 ;
  assign new_n13926 = ~new_n13860 & new_n13925 ;
  assign new_n13927 = new_n2261 & ~new_n13926 ;
  assign new_n13928 = ~new_n2252 & ~new_n13927 ;
  assign new_n13929 = ~new_n2253 & ~new_n13928 ;
  assign new_n13930 = lo0019 & ~new_n13928 ;
  assign new_n13931 = lo0954 & new_n11539 ;
  assign new_n13932 = new_n11539 & ~new_n13931 ;
  assign new_n13933 = ~new_n8324 & ~new_n13932 ;
  assign new_n13934 = ~lo0954 & new_n8324 ;
  assign new_n13935 = ~new_n11539 & new_n13934 ;
  assign new_n13936 = ~new_n13933 & ~new_n13935 ;
  assign new_n13937 = ~lo0895 & ~new_n2261 ;
  assign new_n13938 = lo0895 & ~new_n2261 ;
  assign new_n13939 = new_n2261 & ~new_n13900 ;
  assign new_n13940 = ~new_n13938 & ~new_n13939 ;
  assign new_n13941 = ~new_n13937 & ~new_n13940 ;
  assign new_n13942 = lo0248 & new_n13937 ;
  assign new_n13943 = ~new_n13941 & ~new_n13942 ;
  assign new_n13944 = lo0642 & lo0803 ;
  assign new_n13945 = lo0580 & new_n13944 ;
  assign new_n13946 = lo0226 & new_n13945 ;
  assign new_n13947 = lo0600 & new_n13946 ;
  assign new_n13948 = lo0516 & new_n13947 ;
  assign new_n13949 = lo0399 & new_n13948 ;
  assign new_n13950 = lo0111 & ~new_n13949 ;
  assign new_n13951 = ~lo0111 & new_n13949 ;
  assign new_n13952 = ~new_n13950 & ~new_n13951 ;
  assign new_n13953 = ~new_n13937 & ~new_n13952 ;
  assign new_n13954 = new_n13943 & new_n13953 ;
  assign new_n13955 = new_n13937 & ~new_n13943 ;
  assign new_n13956 = ~new_n5472 & new_n13937 ;
  assign new_n13957 = new_n13943 & new_n13956 ;
  assign new_n13958 = ~new_n13955 & ~new_n13957 ;
  assign new_n13959 = ~new_n13954 & new_n13958 ;
  assign new_n13960 = new_n13943 & ~new_n13959 ;
  assign new_n13961 = new_n13936 & new_n13960 ;
  assign new_n13962 = ~new_n13943 & new_n13959 ;
  assign new_n13963 = ~new_n13960 & ~new_n13962 ;
  assign new_n13964 = ~new_n13936 & ~new_n13963 ;
  assign new_n13965 = lo0763 & ~new_n13943 ;
  assign new_n13966 = ~new_n13959 & new_n13965 ;
  assign new_n13967 = ~new_n13964 & ~new_n13966 ;
  assign new_n13968 = ~new_n13961 & new_n13967 ;
  assign new_n13969 = new_n13928 & ~new_n13968 ;
  assign new_n13970 = ~new_n13930 & ~new_n13969 ;
  assign new_n13971 = lo0020 & ~new_n13928 ;
  assign new_n13972 = lo0954 & new_n11490 ;
  assign new_n13973 = new_n11490 & ~new_n13972 ;
  assign new_n13974 = ~new_n8192 & ~new_n13973 ;
  assign new_n13975 = ~lo0954 & new_n8192 ;
  assign new_n13976 = ~new_n11490 & new_n13975 ;
  assign new_n13977 = ~new_n13974 & ~new_n13976 ;
  assign new_n13978 = ~new_n13937 & ~new_n13943 ;
  assign new_n13979 = ~new_n13977 & new_n13978 ;
  assign new_n13980 = lo0111 & new_n13949 ;
  assign new_n13981 = lo0825 & ~new_n13980 ;
  assign new_n13982 = ~lo0825 & new_n13980 ;
  assign new_n13983 = ~new_n13981 & ~new_n13982 ;
  assign new_n13984 = ~new_n13937 & ~new_n13983 ;
  assign new_n13985 = new_n13943 & new_n13984 ;
  assign new_n13986 = ~new_n13955 & ~new_n13985 ;
  assign new_n13987 = ~new_n13979 & new_n13986 ;
  assign new_n13988 = ~new_n13937 & ~new_n13987 ;
  assign new_n13989 = new_n13937 & new_n13987 ;
  assign new_n13990 = ~new_n13988 & ~new_n13989 ;
  assign new_n13991 = ~new_n5187 & ~new_n13990 ;
  assign new_n13992 = new_n5187 & new_n13988 ;
  assign new_n13993 = lo0823 & new_n13937 ;
  assign new_n13994 = ~new_n13987 & new_n13993 ;
  assign new_n13995 = ~new_n13992 & ~new_n13994 ;
  assign new_n13996 = ~new_n13991 & new_n13995 ;
  assign new_n13997 = new_n13928 & ~new_n13996 ;
  assign new_n13998 = ~new_n13971 & ~new_n13997 ;
  assign new_n13999 = lo0021 & ~new_n13928 ;
  assign new_n14000 = lo0954 & new_n11298 ;
  assign new_n14001 = new_n11298 & ~new_n14000 ;
  assign new_n14002 = ~new_n7675 & ~new_n14001 ;
  assign new_n14003 = ~lo0954 & new_n7675 ;
  assign new_n14004 = ~new_n11298 & new_n14003 ;
  assign new_n14005 = ~new_n14002 & ~new_n14004 ;
  assign new_n14006 = lo0825 & new_n13980 ;
  assign new_n14007 = lo0699 & new_n14006 ;
  assign new_n14008 = lo0720 & new_n14007 ;
  assign new_n14009 = lo0357 & new_n14008 ;
  assign new_n14010 = lo0535 & ~new_n14009 ;
  assign new_n14011 = ~lo0535 & new_n14009 ;
  assign new_n14012 = ~new_n14010 & ~new_n14011 ;
  assign new_n14013 = ~new_n13937 & ~new_n14012 ;
  assign new_n14014 = new_n13943 & new_n14013 ;
  assign new_n14015 = ~new_n3734 & new_n13937 ;
  assign new_n14016 = new_n13943 & new_n14015 ;
  assign new_n14017 = ~new_n13955 & ~new_n14016 ;
  assign new_n14018 = ~new_n14014 & new_n14017 ;
  assign new_n14019 = new_n13943 & ~new_n14018 ;
  assign new_n14020 = new_n14005 & new_n14019 ;
  assign new_n14021 = ~new_n13943 & new_n14018 ;
  assign new_n14022 = ~new_n14019 & ~new_n14021 ;
  assign new_n14023 = ~new_n14005 & ~new_n14022 ;
  assign new_n14024 = lo0537 & ~new_n13943 ;
  assign new_n14025 = ~new_n14018 & new_n14024 ;
  assign new_n14026 = ~new_n14023 & ~new_n14025 ;
  assign new_n14027 = ~new_n14020 & new_n14026 ;
  assign new_n14028 = new_n13928 & ~new_n14027 ;
  assign new_n14029 = ~new_n13999 & ~new_n14028 ;
  assign new_n14030 = lo0022 & ~new_n13928 ;
  assign new_n14031 = lo0954 & new_n11181 ;
  assign new_n14032 = new_n11181 & ~new_n14031 ;
  assign new_n14033 = ~new_n7290 & ~new_n14032 ;
  assign new_n14034 = ~lo0954 & new_n7290 ;
  assign new_n14035 = ~new_n11181 & new_n14034 ;
  assign new_n14036 = ~new_n14033 & ~new_n14035 ;
  assign new_n14037 = ~new_n13940 & ~new_n14036 ;
  assign new_n14038 = lo0535 & new_n14009 ;
  assign new_n14039 = lo0437 & new_n14038 ;
  assign new_n14040 = lo0417 & new_n14039 ;
  assign new_n14041 = lo0556 & ~new_n14040 ;
  assign new_n14042 = ~lo0556 & new_n14040 ;
  assign new_n14043 = ~new_n14041 & ~new_n14042 ;
  assign new_n14044 = new_n2261 & ~new_n14043 ;
  assign new_n14045 = lo0248 & lo0558 ;
  assign new_n14046 = ~lo0248 & ~new_n5560 ;
  assign new_n14047 = ~new_n14045 & ~new_n14046 ;
  assign new_n14048 = ~new_n2261 & ~new_n14047 ;
  assign new_n14049 = ~new_n14044 & ~new_n14048 ;
  assign new_n14050 = new_n13940 & ~new_n14049 ;
  assign new_n14051 = ~new_n14037 & ~new_n14050 ;
  assign new_n14052 = new_n13928 & ~new_n14051 ;
  assign new_n14053 = ~new_n14030 & ~new_n14052 ;
  assign new_n14054 = lo0023 & ~new_n13928 ;
  assign new_n14055 = lo0954 & new_n10432 ;
  assign new_n14056 = new_n10432 & ~new_n14055 ;
  assign new_n14057 = ~new_n3098 & ~new_n14056 ;
  assign new_n14058 = ~lo0954 & new_n3098 ;
  assign new_n14059 = ~new_n10432 & new_n14058 ;
  assign new_n14060 = ~new_n14057 & ~new_n14059 ;
  assign new_n14061 = new_n13978 & ~new_n14060 ;
  assign new_n14062 = lo0556 & new_n14040 ;
  assign new_n14063 = lo0781 & new_n14062 ;
  assign new_n14064 = lo0339 & new_n14063 ;
  assign new_n14065 = lo0318 & new_n14064 ;
  assign new_n14066 = lo0245 & new_n14065 ;
  assign new_n14067 = lo0378 & new_n14066 ;
  assign new_n14068 = lo0275 & new_n14067 ;
  assign new_n14069 = lo0619 & new_n14068 ;
  assign new_n14070 = lo0739 & new_n14069 ;
  assign new_n14071 = lo0843 & new_n14070 ;
  assign new_n14072 = lo0680 & new_n14071 ;
  assign new_n14073 = lo0661 & new_n14072 ;
  assign new_n14074 = lo0294 & new_n14073 ;
  assign new_n14075 = lo0457 & new_n14074 ;
  assign new_n14076 = lo0495 & new_n14075 ;
  assign new_n14077 = lo0476 & ~new_n14076 ;
  assign new_n14078 = ~lo0476 & new_n14076 ;
  assign new_n14079 = ~new_n14077 & ~new_n14078 ;
  assign new_n14080 = ~new_n13937 & ~new_n14079 ;
  assign new_n14081 = new_n13943 & new_n14080 ;
  assign new_n14082 = ~new_n13955 & ~new_n14081 ;
  assign new_n14083 = ~new_n14061 & new_n14082 ;
  assign new_n14084 = ~new_n13937 & ~new_n14083 ;
  assign new_n14085 = new_n13937 & new_n14083 ;
  assign new_n14086 = ~new_n14084 & ~new_n14085 ;
  assign new_n14087 = ~new_n2739 & ~new_n14086 ;
  assign new_n14088 = new_n2739 & new_n14084 ;
  assign new_n14089 = lo0478 & new_n13937 ;
  assign new_n14090 = ~new_n14083 & new_n14089 ;
  assign new_n14091 = ~new_n14088 & ~new_n14090 ;
  assign new_n14092 = ~new_n14087 & new_n14091 ;
  assign new_n14093 = new_n13928 & ~new_n14092 ;
  assign new_n14094 = ~new_n14054 & ~new_n14093 ;
  assign new_n14095 = lo0024 & ~new_n13928 ;
  assign new_n14096 = lo0954 & new_n10482 ;
  assign new_n14097 = new_n10482 & ~new_n14096 ;
  assign new_n14098 = ~new_n3554 & ~new_n14097 ;
  assign new_n14099 = ~lo0954 & new_n3554 ;
  assign new_n14100 = ~new_n10482 & new_n14099 ;
  assign new_n14101 = ~new_n14098 & ~new_n14100 ;
  assign new_n14102 = lo0495 & ~new_n14075 ;
  assign new_n14103 = ~lo0495 & new_n14075 ;
  assign new_n14104 = ~new_n14102 & ~new_n14103 ;
  assign new_n14105 = ~new_n13937 & ~new_n14104 ;
  assign new_n14106 = new_n13943 & new_n14105 ;
  assign new_n14107 = ~new_n3092 & new_n13937 ;
  assign new_n14108 = new_n13943 & new_n14107 ;
  assign new_n14109 = ~new_n13955 & ~new_n14108 ;
  assign new_n14110 = ~new_n14106 & new_n14109 ;
  assign new_n14111 = new_n13943 & ~new_n14110 ;
  assign new_n14112 = new_n14101 & new_n14111 ;
  assign new_n14113 = ~new_n13943 & new_n14110 ;
  assign new_n14114 = ~new_n14111 & ~new_n14113 ;
  assign new_n14115 = ~new_n14101 & ~new_n14114 ;
  assign new_n14116 = lo0497 & ~new_n13943 ;
  assign new_n14117 = ~new_n14110 & new_n14116 ;
  assign new_n14118 = ~new_n14115 & ~new_n14117 ;
  assign new_n14119 = ~new_n14112 & new_n14118 ;
  assign new_n14120 = new_n13928 & ~new_n14119 ;
  assign new_n14121 = ~new_n14095 & ~new_n14120 ;
  assign new_n14122 = lo0025 & ~new_n13928 ;
  assign new_n14123 = lo0954 & new_n10529 ;
  assign new_n14124 = new_n10529 & ~new_n14123 ;
  assign new_n14125 = ~new_n3919 & ~new_n14124 ;
  assign new_n14126 = ~lo0954 & new_n3919 ;
  assign new_n14127 = ~new_n10529 & new_n14126 ;
  assign new_n14128 = ~new_n14125 & ~new_n14127 ;
  assign new_n14129 = new_n13978 & ~new_n14128 ;
  assign new_n14130 = lo0457 & ~new_n14074 ;
  assign new_n14131 = ~lo0457 & new_n14074 ;
  assign new_n14132 = ~new_n14130 & ~new_n14131 ;
  assign new_n14133 = ~new_n13937 & ~new_n14132 ;
  assign new_n14134 = new_n13943 & new_n14133 ;
  assign new_n14135 = ~new_n13955 & ~new_n14134 ;
  assign new_n14136 = ~new_n14129 & new_n14135 ;
  assign new_n14137 = ~new_n13937 & ~new_n14136 ;
  assign new_n14138 = new_n13937 & new_n14136 ;
  assign new_n14139 = ~new_n14137 & ~new_n14138 ;
  assign new_n14140 = ~new_n3001 & ~new_n14139 ;
  assign new_n14141 = new_n3001 & new_n14137 ;
  assign new_n14142 = lo0459 & new_n13937 ;
  assign new_n14143 = ~new_n14136 & new_n14142 ;
  assign new_n14144 = ~new_n14141 & ~new_n14143 ;
  assign new_n14145 = ~new_n14140 & new_n14144 ;
  assign new_n14146 = new_n13928 & ~new_n14145 ;
  assign new_n14147 = ~new_n14122 & ~new_n14146 ;
  assign new_n14148 = lo0026 & ~new_n13928 ;
  assign new_n14149 = lo0954 & new_n10575 ;
  assign new_n14150 = new_n10575 & ~new_n14149 ;
  assign new_n14151 = ~new_n4278 & ~new_n14150 ;
  assign new_n14152 = ~lo0954 & new_n4278 ;
  assign new_n14153 = ~new_n10575 & new_n14152 ;
  assign new_n14154 = ~new_n14151 & ~new_n14153 ;
  assign new_n14155 = lo0294 & ~new_n14073 ;
  assign new_n14156 = ~lo0294 & new_n14073 ;
  assign new_n14157 = ~new_n14155 & ~new_n14156 ;
  assign new_n14158 = ~new_n13937 & ~new_n14157 ;
  assign new_n14159 = new_n13943 & new_n14158 ;
  assign new_n14160 = ~new_n3464 & new_n13937 ;
  assign new_n14161 = new_n13943 & new_n14160 ;
  assign new_n14162 = ~new_n13955 & ~new_n14161 ;
  assign new_n14163 = ~new_n14159 & new_n14162 ;
  assign new_n14164 = new_n13943 & ~new_n14163 ;
  assign new_n14165 = new_n14154 & new_n14164 ;
  assign new_n14166 = ~new_n13943 & new_n14163 ;
  assign new_n14167 = ~new_n14164 & ~new_n14166 ;
  assign new_n14168 = ~new_n14154 & ~new_n14167 ;
  assign new_n14169 = lo0296 & ~new_n13943 ;
  assign new_n14170 = ~new_n14163 & new_n14169 ;
  assign new_n14171 = ~new_n14168 & ~new_n14170 ;
  assign new_n14172 = ~new_n14165 & new_n14171 ;
  assign new_n14173 = new_n13928 & ~new_n14172 ;
  assign new_n14174 = ~new_n14148 & ~new_n14173 ;
  assign new_n14175 = lo0027 & ~new_n13928 ;
  assign new_n14176 = lo0954 & new_n10622 ;
  assign new_n14177 = new_n10622 & ~new_n14176 ;
  assign new_n14178 = ~new_n4640 & ~new_n14177 ;
  assign new_n14179 = ~lo0954 & new_n4640 ;
  assign new_n14180 = ~new_n10622 & new_n14179 ;
  assign new_n14181 = ~new_n14178 & ~new_n14180 ;
  assign new_n14182 = new_n13978 & ~new_n14181 ;
  assign new_n14183 = lo0661 & ~new_n14072 ;
  assign new_n14184 = ~lo0661 & new_n14072 ;
  assign new_n14185 = ~new_n14183 & ~new_n14184 ;
  assign new_n14186 = ~new_n13937 & ~new_n14185 ;
  assign new_n14187 = new_n13943 & new_n14186 ;
  assign new_n14188 = ~new_n13955 & ~new_n14187 ;
  assign new_n14189 = ~new_n14182 & new_n14188 ;
  assign new_n14190 = ~new_n13937 & ~new_n14189 ;
  assign new_n14191 = new_n13937 & new_n14189 ;
  assign new_n14192 = ~new_n14190 & ~new_n14191 ;
  assign new_n14193 = ~new_n3817 & ~new_n14192 ;
  assign new_n14194 = new_n3817 & new_n14190 ;
  assign new_n14195 = lo0663 & new_n13937 ;
  assign new_n14196 = ~new_n14189 & new_n14195 ;
  assign new_n14197 = ~new_n14194 & ~new_n14196 ;
  assign new_n14198 = ~new_n14193 & new_n14197 ;
  assign new_n14199 = new_n13928 & ~new_n14198 ;
  assign new_n14200 = ~new_n14175 & ~new_n14199 ;
  assign new_n14201 = lo0028 & ~new_n13928 ;
  assign new_n14202 = lo0954 & new_n10667 ;
  assign new_n14203 = new_n10667 & ~new_n14202 ;
  assign new_n14204 = ~new_n5002 & ~new_n14203 ;
  assign new_n14205 = ~lo0954 & new_n5002 ;
  assign new_n14206 = ~new_n10667 & new_n14205 ;
  assign new_n14207 = ~new_n14204 & ~new_n14206 ;
  assign new_n14208 = lo0680 & ~new_n14071 ;
  assign new_n14209 = ~lo0680 & new_n14071 ;
  assign new_n14210 = ~new_n14208 & ~new_n14209 ;
  assign new_n14211 = ~new_n13937 & ~new_n14210 ;
  assign new_n14212 = new_n13943 & new_n14211 ;
  assign new_n14213 = ~new_n4097 & new_n13937 ;
  assign new_n14214 = new_n13943 & new_n14213 ;
  assign new_n14215 = ~new_n13955 & ~new_n14214 ;
  assign new_n14216 = ~new_n14212 & new_n14215 ;
  assign new_n14217 = new_n13943 & ~new_n14216 ;
  assign new_n14218 = new_n14207 & new_n14217 ;
  assign new_n14219 = ~new_n13943 & new_n14216 ;
  assign new_n14220 = ~new_n14217 & ~new_n14219 ;
  assign new_n14221 = ~new_n14207 & ~new_n14220 ;
  assign new_n14222 = lo0682 & ~new_n13943 ;
  assign new_n14223 = ~new_n14216 & new_n14222 ;
  assign new_n14224 = ~new_n14221 & ~new_n14223 ;
  assign new_n14225 = ~new_n14218 & new_n14224 ;
  assign new_n14226 = new_n13928 & ~new_n14225 ;
  assign new_n14227 = ~new_n14201 & ~new_n14226 ;
  assign new_n14228 = lo0029 & ~new_n13928 ;
  assign new_n14229 = lo0954 & new_n10714 ;
  assign new_n14230 = new_n10714 & ~new_n14229 ;
  assign new_n14231 = ~new_n5286 & ~new_n14230 ;
  assign new_n14232 = ~lo0954 & new_n5286 ;
  assign new_n14233 = ~new_n10714 & new_n14232 ;
  assign new_n14234 = ~new_n14231 & ~new_n14233 ;
  assign new_n14235 = new_n13978 & ~new_n14234 ;
  assign new_n14236 = lo0843 & ~new_n14070 ;
  assign new_n14237 = ~lo0843 & new_n14070 ;
  assign new_n14238 = ~new_n14236 & ~new_n14237 ;
  assign new_n14239 = ~new_n13937 & ~new_n14238 ;
  assign new_n14240 = new_n13943 & new_n14239 ;
  assign new_n14241 = ~new_n13955 & ~new_n14240 ;
  assign new_n14242 = ~new_n14235 & new_n14241 ;
  assign new_n14243 = ~new_n13937 & ~new_n14242 ;
  assign new_n14244 = new_n13937 & new_n14242 ;
  assign new_n14245 = ~new_n14243 & ~new_n14244 ;
  assign new_n14246 = ~new_n4541 & ~new_n14245 ;
  assign new_n14247 = new_n4541 & new_n14243 ;
  assign new_n14248 = lo0845 & new_n13937 ;
  assign new_n14249 = ~new_n14242 & new_n14248 ;
  assign new_n14250 = ~new_n14247 & ~new_n14249 ;
  assign new_n14251 = ~new_n14246 & new_n14250 ;
  assign new_n14252 = new_n13928 & ~new_n14251 ;
  assign new_n14253 = ~new_n14228 & ~new_n14252 ;
  assign new_n14254 = lo0030 & ~new_n13928 ;
  assign new_n14255 = lo0954 & new_n10759 ;
  assign new_n14256 = new_n10759 & ~new_n14255 ;
  assign new_n14257 = ~new_n5570 & ~new_n14256 ;
  assign new_n14258 = ~lo0954 & new_n5570 ;
  assign new_n14259 = ~new_n10759 & new_n14258 ;
  assign new_n14260 = ~new_n14257 & ~new_n14259 ;
  assign new_n14261 = lo0739 & ~new_n14069 ;
  assign new_n14262 = ~lo0739 & new_n14069 ;
  assign new_n14263 = ~new_n14261 & ~new_n14262 ;
  assign new_n14264 = ~new_n13937 & ~new_n14263 ;
  assign new_n14265 = new_n13943 & new_n14264 ;
  assign new_n14266 = ~new_n4818 & new_n13937 ;
  assign new_n14267 = new_n13943 & new_n14266 ;
  assign new_n14268 = ~new_n13955 & ~new_n14267 ;
  assign new_n14269 = ~new_n14265 & new_n14268 ;
  assign new_n14270 = new_n13943 & ~new_n14269 ;
  assign new_n14271 = new_n14260 & new_n14270 ;
  assign new_n14272 = ~new_n13943 & new_n14269 ;
  assign new_n14273 = ~new_n14270 & ~new_n14272 ;
  assign new_n14274 = ~new_n14260 & ~new_n14273 ;
  assign new_n14275 = lo0741 & ~new_n13943 ;
  assign new_n14276 = ~new_n14269 & new_n14275 ;
  assign new_n14277 = ~new_n14274 & ~new_n14276 ;
  assign new_n14278 = ~new_n14271 & new_n14277 ;
  assign new_n14279 = new_n13928 & ~new_n14278 ;
  assign new_n14280 = ~new_n14254 & ~new_n14279 ;
  assign new_n14281 = lo0031 & ~new_n13928 ;
  assign new_n14282 = lo0954 & new_n10806 ;
  assign new_n14283 = new_n10806 & ~new_n14282 ;
  assign new_n14284 = ~new_n5796 & ~new_n14283 ;
  assign new_n14285 = ~lo0954 & new_n5796 ;
  assign new_n14286 = ~new_n10806 & new_n14285 ;
  assign new_n14287 = ~new_n14284 & ~new_n14286 ;
  assign new_n14288 = new_n13978 & ~new_n14287 ;
  assign new_n14289 = lo0619 & ~new_n14068 ;
  assign new_n14290 = ~lo0619 & new_n14068 ;
  assign new_n14291 = ~new_n14289 & ~new_n14290 ;
  assign new_n14292 = ~new_n13937 & ~new_n14291 ;
  assign new_n14293 = new_n13943 & new_n14292 ;
  assign new_n14294 = ~new_n13955 & ~new_n14293 ;
  assign new_n14295 = ~new_n14288 & new_n14294 ;
  assign new_n14296 = ~new_n13937 & ~new_n14295 ;
  assign new_n14297 = new_n13937 & new_n14295 ;
  assign new_n14298 = ~new_n14296 & ~new_n14297 ;
  assign new_n14299 = ~new_n2824 & ~new_n14298 ;
  assign new_n14300 = new_n2824 & new_n14296 ;
  assign new_n14301 = lo0621 & new_n13937 ;
  assign new_n14302 = ~new_n14295 & new_n14301 ;
  assign new_n14303 = ~new_n14300 & ~new_n14302 ;
  assign new_n14304 = ~new_n14299 & new_n14303 ;
  assign new_n14305 = new_n13928 & ~new_n14304 ;
  assign new_n14306 = ~new_n14281 & ~new_n14305 ;
  assign new_n14307 = lo0032 & ~new_n13928 ;
  assign new_n14308 = lo0954 & new_n10851 ;
  assign new_n14309 = new_n10851 & ~new_n14308 ;
  assign new_n14310 = ~new_n6022 & ~new_n14309 ;
  assign new_n14311 = ~lo0954 & new_n6022 ;
  assign new_n14312 = ~new_n10851 & new_n14311 ;
  assign new_n14313 = ~new_n14310 & ~new_n14312 ;
  assign new_n14314 = lo0275 & ~new_n14067 ;
  assign new_n14315 = ~lo0275 & new_n14067 ;
  assign new_n14316 = ~new_n14314 & ~new_n14315 ;
  assign new_n14317 = ~new_n13937 & ~new_n14316 ;
  assign new_n14318 = new_n13943 & new_n14317 ;
  assign new_n14319 = ~new_n3549 & new_n13937 ;
  assign new_n14320 = new_n13943 & new_n14319 ;
  assign new_n14321 = ~new_n13955 & ~new_n14320 ;
  assign new_n14322 = ~new_n14318 & new_n14321 ;
  assign new_n14323 = new_n13943 & ~new_n14322 ;
  assign new_n14324 = new_n14313 & new_n14323 ;
  assign new_n14325 = ~new_n13943 & new_n14322 ;
  assign new_n14326 = ~new_n14323 & ~new_n14325 ;
  assign new_n14327 = ~new_n14313 & ~new_n14326 ;
  assign new_n14328 = lo0277 & ~new_n13943 ;
  assign new_n14329 = ~new_n14322 & new_n14328 ;
  assign new_n14330 = ~new_n14327 & ~new_n14329 ;
  assign new_n14331 = ~new_n14324 & new_n14330 ;
  assign new_n14332 = new_n13928 & ~new_n14331 ;
  assign new_n14333 = ~new_n14307 & ~new_n14332 ;
  assign new_n14334 = lo0033 & ~new_n13928 ;
  assign new_n14335 = lo0954 & new_n10898 ;
  assign new_n14336 = new_n10898 & ~new_n14335 ;
  assign new_n14337 = ~new_n6252 & ~new_n14336 ;
  assign new_n14338 = ~lo0954 & new_n6252 ;
  assign new_n14339 = ~new_n10898 & new_n14338 ;
  assign new_n14340 = ~new_n14337 & ~new_n14339 ;
  assign new_n14341 = new_n13978 & ~new_n14340 ;
  assign new_n14342 = lo0378 & ~new_n14066 ;
  assign new_n14343 = ~lo0378 & new_n14066 ;
  assign new_n14344 = ~new_n14342 & ~new_n14343 ;
  assign new_n14345 = ~new_n13937 & ~new_n14344 ;
  assign new_n14346 = new_n13943 & new_n14345 ;
  assign new_n14347 = ~new_n13955 & ~new_n14346 ;
  assign new_n14348 = ~new_n14341 & new_n14347 ;
  assign new_n14349 = ~new_n13937 & ~new_n14348 ;
  assign new_n14350 = new_n13937 & new_n14348 ;
  assign new_n14351 = ~new_n14349 & ~new_n14350 ;
  assign new_n14352 = ~new_n3908 & ~new_n14351 ;
  assign new_n14353 = new_n3908 & new_n14349 ;
  assign new_n14354 = lo0380 & new_n13937 ;
  assign new_n14355 = ~new_n14348 & new_n14354 ;
  assign new_n14356 = ~new_n14353 & ~new_n14355 ;
  assign new_n14357 = ~new_n14352 & new_n14356 ;
  assign new_n14358 = new_n13928 & ~new_n14357 ;
  assign new_n14359 = ~new_n14334 & ~new_n14358 ;
  assign new_n14360 = lo0034 & ~new_n13928 ;
  assign new_n14361 = lo0954 & new_n10943 ;
  assign new_n14362 = new_n10943 & ~new_n14361 ;
  assign new_n14363 = ~new_n6487 & ~new_n14362 ;
  assign new_n14364 = ~lo0954 & new_n6487 ;
  assign new_n14365 = ~new_n10943 & new_n14364 ;
  assign new_n14366 = ~new_n14363 & ~new_n14365 ;
  assign new_n14367 = lo0245 & ~new_n14065 ;
  assign new_n14368 = ~lo0245 & new_n14065 ;
  assign new_n14369 = ~new_n14367 & ~new_n14368 ;
  assign new_n14370 = ~new_n13937 & ~new_n14369 ;
  assign new_n14371 = new_n13943 & new_n14370 ;
  assign new_n14372 = ~new_n4268 & new_n13937 ;
  assign new_n14373 = new_n13943 & new_n14372 ;
  assign new_n14374 = ~new_n13955 & ~new_n14373 ;
  assign new_n14375 = ~new_n14371 & new_n14374 ;
  assign new_n14376 = new_n13943 & ~new_n14375 ;
  assign new_n14377 = new_n14366 & new_n14376 ;
  assign new_n14378 = ~new_n13943 & new_n14375 ;
  assign new_n14379 = ~new_n14376 & ~new_n14378 ;
  assign new_n14380 = ~new_n14366 & ~new_n14379 ;
  assign new_n14381 = lo0381 & ~new_n13943 ;
  assign new_n14382 = ~new_n14375 & new_n14381 ;
  assign new_n14383 = ~new_n14380 & ~new_n14382 ;
  assign new_n14384 = ~new_n14377 & new_n14383 ;
  assign new_n14385 = new_n13928 & ~new_n14384 ;
  assign new_n14386 = ~new_n14360 & ~new_n14385 ;
  assign new_n14387 = lo0035 & ~new_n13928 ;
  assign new_n14388 = lo0954 & new_n10990 ;
  assign new_n14389 = new_n10990 & ~new_n14388 ;
  assign new_n14390 = ~new_n6717 & ~new_n14389 ;
  assign new_n14391 = ~lo0954 & new_n6717 ;
  assign new_n14392 = ~new_n10990 & new_n14391 ;
  assign new_n14393 = ~new_n14390 & ~new_n14392 ;
  assign new_n14394 = new_n13978 & ~new_n14393 ;
  assign new_n14395 = lo0318 & ~new_n14064 ;
  assign new_n14396 = ~lo0318 & new_n14064 ;
  assign new_n14397 = ~new_n14395 & ~new_n14396 ;
  assign new_n14398 = ~new_n13937 & ~new_n14397 ;
  assign new_n14399 = new_n13943 & new_n14398 ;
  assign new_n14400 = ~new_n13955 & ~new_n14399 ;
  assign new_n14401 = ~new_n14394 & new_n14400 ;
  assign new_n14402 = ~new_n13937 & ~new_n14401 ;
  assign new_n14403 = new_n13937 & new_n14401 ;
  assign new_n14404 = ~new_n14402 & ~new_n14403 ;
  assign new_n14405 = ~new_n4630 & ~new_n14404 ;
  assign new_n14406 = new_n4630 & new_n14402 ;
  assign new_n14407 = lo0320 & new_n13937 ;
  assign new_n14408 = ~new_n14401 & new_n14407 ;
  assign new_n14409 = ~new_n14406 & ~new_n14408 ;
  assign new_n14410 = ~new_n14405 & new_n14409 ;
  assign new_n14411 = new_n13928 & ~new_n14410 ;
  assign new_n14412 = ~new_n14387 & ~new_n14411 ;
  assign new_n14413 = lo0036 & ~new_n13928 ;
  assign new_n14414 = lo0954 & new_n11035 ;
  assign new_n14415 = new_n11035 & ~new_n14414 ;
  assign new_n14416 = ~new_n6942 & ~new_n14415 ;
  assign new_n14417 = ~lo0954 & new_n6942 ;
  assign new_n14418 = ~new_n11035 & new_n14417 ;
  assign new_n14419 = ~new_n14416 & ~new_n14418 ;
  assign new_n14420 = lo0339 & ~new_n14063 ;
  assign new_n14421 = ~lo0339 & new_n14063 ;
  assign new_n14422 = ~new_n14420 & ~new_n14421 ;
  assign new_n14423 = ~new_n13937 & ~new_n14422 ;
  assign new_n14424 = new_n13943 & new_n14423 ;
  assign new_n14425 = ~new_n4992 & new_n13937 ;
  assign new_n14426 = new_n13943 & new_n14425 ;
  assign new_n14427 = ~new_n13955 & ~new_n14426 ;
  assign new_n14428 = ~new_n14424 & new_n14427 ;
  assign new_n14429 = new_n13943 & ~new_n14428 ;
  assign new_n14430 = new_n14419 & new_n14429 ;
  assign new_n14431 = ~new_n13943 & new_n14428 ;
  assign new_n14432 = ~new_n14429 & ~new_n14431 ;
  assign new_n14433 = ~new_n14419 & ~new_n14432 ;
  assign new_n14434 = lo0341 & ~new_n13943 ;
  assign new_n14435 = ~new_n14428 & new_n14434 ;
  assign new_n14436 = ~new_n14433 & ~new_n14435 ;
  assign new_n14437 = ~new_n14430 & new_n14436 ;
  assign new_n14438 = new_n13928 & ~new_n14437 ;
  assign new_n14439 = ~new_n14413 & ~new_n14438 ;
  assign new_n14440 = lo0037 & ~new_n13928 ;
  assign new_n14441 = lo0954 & new_n11082 ;
  assign new_n14442 = new_n11082 & ~new_n14441 ;
  assign new_n14443 = ~new_n7165 & ~new_n14442 ;
  assign new_n14444 = ~lo0954 & new_n7165 ;
  assign new_n14445 = ~new_n11082 & new_n14444 ;
  assign new_n14446 = ~new_n14443 & ~new_n14445 ;
  assign new_n14447 = new_n13978 & ~new_n14446 ;
  assign new_n14448 = lo0781 & ~new_n14062 ;
  assign new_n14449 = ~lo0781 & new_n14062 ;
  assign new_n14450 = ~new_n14448 & ~new_n14449 ;
  assign new_n14451 = ~new_n13937 & ~new_n14450 ;
  assign new_n14452 = new_n13943 & new_n14451 ;
  assign new_n14453 = ~new_n13955 & ~new_n14452 ;
  assign new_n14454 = ~new_n14447 & new_n14453 ;
  assign new_n14455 = ~new_n13937 & ~new_n14454 ;
  assign new_n14456 = new_n13937 & new_n14454 ;
  assign new_n14457 = ~new_n14455 & ~new_n14456 ;
  assign new_n14458 = ~new_n5276 & ~new_n14457 ;
  assign new_n14459 = new_n5276 & new_n14455 ;
  assign new_n14460 = lo0783 & new_n13937 ;
  assign new_n14461 = ~new_n14454 & new_n14460 ;
  assign new_n14462 = ~new_n14459 & ~new_n14461 ;
  assign new_n14463 = ~new_n14458 & new_n14462 ;
  assign new_n14464 = new_n13928 & ~new_n14463 ;
  assign new_n14465 = ~new_n14440 & ~new_n14464 ;
  assign new_n14466 = lo0038 & ~new_n13928 ;
  assign new_n14467 = lo0954 & new_n11136 ;
  assign new_n14468 = new_n11136 & ~new_n14467 ;
  assign new_n14469 = ~new_n7420 & ~new_n14468 ;
  assign new_n14470 = ~lo0954 & new_n7420 ;
  assign new_n14471 = ~new_n11136 & new_n14470 ;
  assign new_n14472 = ~new_n14469 & ~new_n14471 ;
  assign new_n14473 = lo0417 & ~new_n14039 ;
  assign new_n14474 = ~lo0417 & new_n14039 ;
  assign new_n14475 = ~new_n14473 & ~new_n14474 ;
  assign new_n14476 = ~new_n13937 & ~new_n14475 ;
  assign new_n14477 = new_n13943 & new_n14476 ;
  assign new_n14478 = ~new_n2910 & new_n13937 ;
  assign new_n14479 = new_n13943 & new_n14478 ;
  assign new_n14480 = ~new_n13955 & ~new_n14479 ;
  assign new_n14481 = ~new_n14477 & new_n14480 ;
  assign new_n14482 = new_n13943 & ~new_n14481 ;
  assign new_n14483 = new_n14472 & new_n14482 ;
  assign new_n14484 = ~new_n13943 & new_n14481 ;
  assign new_n14485 = ~new_n14482 & ~new_n14484 ;
  assign new_n14486 = ~new_n14472 & ~new_n14485 ;
  assign new_n14487 = lo0538 & ~new_n13943 ;
  assign new_n14488 = ~new_n14481 & new_n14487 ;
  assign new_n14489 = ~new_n14486 & ~new_n14488 ;
  assign new_n14490 = ~new_n14483 & new_n14489 ;
  assign new_n14491 = new_n13928 & ~new_n14490 ;
  assign new_n14492 = ~new_n14466 & ~new_n14491 ;
  assign new_n14493 = lo0039 & ~new_n13928 ;
  assign new_n14494 = lo0954 & new_n11250 ;
  assign new_n14495 = new_n11250 & ~new_n14494 ;
  assign new_n14496 = ~new_n7551 & ~new_n14495 ;
  assign new_n14497 = ~lo0954 & new_n7551 ;
  assign new_n14498 = ~new_n11250 & new_n14497 ;
  assign new_n14499 = ~new_n14496 & ~new_n14498 ;
  assign new_n14500 = new_n13978 & ~new_n14499 ;
  assign new_n14501 = lo0437 & ~new_n14038 ;
  assign new_n14502 = ~lo0437 & new_n14038 ;
  assign new_n14503 = ~new_n14501 & ~new_n14502 ;
  assign new_n14504 = ~new_n13937 & ~new_n14503 ;
  assign new_n14505 = new_n13943 & new_n14504 ;
  assign new_n14506 = ~new_n13955 & ~new_n14505 ;
  assign new_n14507 = ~new_n14500 & new_n14506 ;
  assign new_n14508 = ~new_n13937 & ~new_n14507 ;
  assign new_n14509 = new_n13937 & new_n14507 ;
  assign new_n14510 = ~new_n14508 & ~new_n14509 ;
  assign new_n14511 = ~new_n3383 & ~new_n14510 ;
  assign new_n14512 = new_n3383 & new_n14508 ;
  assign new_n14513 = lo0439 & new_n13937 ;
  assign new_n14514 = ~new_n14507 & new_n14513 ;
  assign new_n14515 = ~new_n14512 & ~new_n14514 ;
  assign new_n14516 = ~new_n14511 & new_n14515 ;
  assign new_n14517 = new_n13928 & ~new_n14516 ;
  assign new_n14518 = ~new_n14493 & ~new_n14517 ;
  assign new_n14519 = lo0040 & ~new_n13928 ;
  assign new_n14520 = lo0954 & new_n11443 ;
  assign new_n14521 = new_n11443 & ~new_n14520 ;
  assign new_n14522 = ~new_n8064 & ~new_n14521 ;
  assign new_n14523 = ~lo0954 & new_n8064 ;
  assign new_n14524 = ~new_n11443 & new_n14523 ;
  assign new_n14525 = ~new_n14522 & ~new_n14524 ;
  assign new_n14526 = lo0699 & ~new_n14006 ;
  assign new_n14527 = ~lo0699 & new_n14006 ;
  assign new_n14528 = ~new_n14526 & ~new_n14527 ;
  assign new_n14529 = ~new_n13937 & ~new_n14528 ;
  assign new_n14530 = new_n13943 & new_n14529 ;
  assign new_n14531 = ~new_n4904 & new_n13937 ;
  assign new_n14532 = new_n13943 & new_n14531 ;
  assign new_n14533 = ~new_n13955 & ~new_n14532 ;
  assign new_n14534 = ~new_n14530 & new_n14533 ;
  assign new_n14535 = new_n13943 & ~new_n14534 ;
  assign new_n14536 = new_n14525 & new_n14535 ;
  assign new_n14537 = ~new_n13943 & new_n14534 ;
  assign new_n14538 = ~new_n14535 & ~new_n14537 ;
  assign new_n14539 = ~new_n14525 & ~new_n14538 ;
  assign new_n14540 = lo0701 & ~new_n13943 ;
  assign new_n14541 = ~new_n14534 & new_n14540 ;
  assign new_n14542 = ~new_n14539 & ~new_n14541 ;
  assign new_n14543 = ~new_n14536 & new_n14542 ;
  assign new_n14544 = new_n13928 & ~new_n14543 ;
  assign new_n14545 = ~new_n14519 & ~new_n14544 ;
  assign new_n14546 = lo0041 & ~new_n13928 ;
  assign new_n14547 = lo0954 & new_n11347 ;
  assign new_n14548 = new_n11347 & ~new_n14547 ;
  assign new_n14549 = ~new_n7799 & ~new_n14548 ;
  assign new_n14550 = ~lo0954 & new_n7799 ;
  assign new_n14551 = ~new_n11347 & new_n14550 ;
  assign new_n14552 = ~new_n14549 & ~new_n14551 ;
  assign new_n14553 = new_n13978 & ~new_n14552 ;
  assign new_n14554 = lo0357 & ~new_n14008 ;
  assign new_n14555 = ~lo0357 & new_n14008 ;
  assign new_n14556 = ~new_n14554 & ~new_n14555 ;
  assign new_n14557 = ~new_n13937 & ~new_n14556 ;
  assign new_n14558 = new_n13943 & new_n14557 ;
  assign new_n14559 = ~new_n13955 & ~new_n14558 ;
  assign new_n14560 = ~new_n14553 & new_n14559 ;
  assign new_n14561 = ~new_n13937 & ~new_n14560 ;
  assign new_n14562 = new_n13937 & new_n14560 ;
  assign new_n14563 = ~new_n14561 & ~new_n14562 ;
  assign new_n14564 = ~new_n4179 & ~new_n14563 ;
  assign new_n14565 = new_n4179 & new_n14561 ;
  assign new_n14566 = lo0359 & new_n13937 ;
  assign new_n14567 = ~new_n14560 & new_n14566 ;
  assign new_n14568 = ~new_n14565 & ~new_n14567 ;
  assign new_n14569 = ~new_n14564 & new_n14568 ;
  assign new_n14570 = new_n13928 & ~new_n14569 ;
  assign new_n14571 = ~new_n14546 & ~new_n14570 ;
  assign new_n14572 = lo0042 & ~new_n13928 ;
  assign new_n14573 = lo0954 & new_n11394 ;
  assign new_n14574 = new_n11394 & ~new_n14573 ;
  assign new_n14575 = ~new_n7923 & ~new_n14574 ;
  assign new_n14576 = ~lo0954 & new_n7923 ;
  assign new_n14577 = ~new_n11394 & new_n14576 ;
  assign new_n14578 = ~new_n14575 & ~new_n14577 ;
  assign new_n14579 = lo0720 & ~new_n14007 ;
  assign new_n14580 = ~lo0720 & new_n14007 ;
  assign new_n14581 = ~new_n14579 & ~new_n14580 ;
  assign new_n14582 = ~new_n13937 & ~new_n14581 ;
  assign new_n14583 = new_n13943 & new_n14582 ;
  assign new_n14584 = ~new_n4461 & new_n13937 ;
  assign new_n14585 = new_n13943 & new_n14584 ;
  assign new_n14586 = ~new_n13955 & ~new_n14585 ;
  assign new_n14587 = ~new_n14583 & new_n14586 ;
  assign new_n14588 = new_n13943 & ~new_n14587 ;
  assign new_n14589 = new_n14578 & new_n14588 ;
  assign new_n14590 = ~new_n13943 & new_n14587 ;
  assign new_n14591 = ~new_n14588 & ~new_n14590 ;
  assign new_n14592 = ~new_n14578 & ~new_n14591 ;
  assign new_n14593 = lo0721 & ~new_n13943 ;
  assign new_n14594 = ~new_n14587 & new_n14593 ;
  assign new_n14595 = ~new_n14592 & ~new_n14594 ;
  assign new_n14596 = ~new_n14589 & new_n14595 ;
  assign new_n14597 = new_n13928 & ~new_n14596 ;
  assign new_n14598 = ~new_n14572 & ~new_n14597 ;
  assign new_n14599 = lo0043 & ~new_n13928 ;
  assign new_n14600 = new_n2261 & new_n13926 ;
  assign new_n14601 = ~lo0113 & ~lo0114 ;
  assign new_n14602 = lo0895 & ~new_n13907 ;
  assign new_n14603 = lo0248 & lo0804 ;
  assign new_n14604 = ~lo0248 & ~new_n7138 ;
  assign new_n14605 = ~new_n14603 & ~new_n14604 ;
  assign new_n14606 = ~lo0895 & ~new_n14605 ;
  assign new_n14607 = ~new_n14602 & ~new_n14606 ;
  assign new_n14608 = new_n14601 & new_n14607 ;
  assign new_n14609 = ~lo0113 & lo0114 ;
  assign new_n14610 = lo0113 & ~lo0114 ;
  assign new_n14611 = ~new_n14609 & ~new_n14610 ;
  assign new_n14612 = ~new_n14608 & new_n14611 ;
  assign new_n14613 = lo0895 & ~new_n10308 ;
  assign new_n14614 = lo0248 & lo0762 ;
  assign new_n14615 = ~lo0248 & ~new_n2619 ;
  assign new_n14616 = ~new_n14614 & ~new_n14615 ;
  assign new_n14617 = ~lo0895 & ~new_n14616 ;
  assign new_n14618 = ~new_n14613 & ~new_n14617 ;
  assign new_n14619 = new_n14601 & new_n14618 ;
  assign new_n14620 = ~new_n14607 & new_n14619 ;
  assign new_n14621 = new_n14612 & new_n14620 ;
  assign new_n14622 = ~new_n14607 & new_n14609 ;
  assign new_n14623 = ~new_n14610 & ~new_n14622 ;
  assign new_n14624 = ~new_n14612 & ~new_n14623 ;
  assign new_n14625 = ~new_n14621 & ~new_n14624 ;
  assign new_n14626 = ~new_n2261 & ~new_n14625 ;
  assign new_n14627 = ~new_n14600 & ~new_n14626 ;
  assign new_n14628 = new_n13928 & ~new_n14627 ;
  assign new_n14629 = ~new_n14599 & ~new_n14628 ;
  assign new_n14630 = lo0044 & new_n2252 ;
  assign new_n14631 = ~lo1290 & ~new_n2261 ;
  assign new_n14632 = ~new_n2252 & ~new_n14631 ;
  assign new_n14633 = ~new_n14600 & new_n14632 ;
  assign new_n14634 = ~new_n14630 & ~new_n14633 ;
  assign new_n14635 = lo0045 & ~new_n13928 ;
  assign new_n14636 = new_n14612 & ~new_n14620 ;
  assign new_n14637 = ~new_n14624 & ~new_n14636 ;
  assign new_n14638 = ~new_n2261 & ~new_n14637 ;
  assign new_n14639 = ~new_n14600 & ~new_n14638 ;
  assign new_n14640 = new_n13928 & ~new_n14639 ;
  assign new_n14641 = ~new_n14635 & ~new_n14640 ;
  assign new_n14642 = lo0046 & ~new_n13928 ;
  assign new_n14643 = new_n13910 & new_n14600 ;
  assign new_n14644 = new_n14601 & ~new_n14618 ;
  assign new_n14645 = ~new_n14609 & ~new_n14644 ;
  assign new_n14646 = new_n14607 & ~new_n14645 ;
  assign new_n14647 = ~new_n14610 & ~new_n14646 ;
  assign new_n14648 = ~new_n2261 & ~new_n14647 ;
  assign new_n14649 = ~new_n14643 & ~new_n14648 ;
  assign new_n14650 = new_n13928 & ~new_n14649 ;
  assign new_n14651 = ~new_n14642 & ~new_n14650 ;
  assign new_n14652 = lo0048 & lo0050 ;
  assign new_n14653 = lo0047 & ~new_n14652 ;
  assign new_n14654 = lo0896 & new_n14652 ;
  assign new_n14655 = ~new_n14653 & ~new_n14654 ;
  assign new_n14656 = lo0050 & lo0897 ;
  assign new_n14657 = ~new_n14655 & ~new_n14656 ;
  assign new_n14658 = lo1425 & lo1428 ;
  assign new_n14659 = ~lo1426 & ~lo1427 ;
  assign new_n14660 = new_n14658 & new_n14659 ;
  assign new_n14661 = ~lo0017 & ~lo0050 ;
  assign new_n14662 = ~lo0017 & lo0048 ;
  assign new_n14663 = ~new_n14661 & new_n14662 ;
  assign new_n14664 = lo0049 & new_n14661 ;
  assign new_n14665 = ~new_n14663 & ~new_n14664 ;
  assign new_n14666 = ~lo1429 & ~lo1430 ;
  assign new_n14667 = ~lo0898 & new_n14666 ;
  assign new_n14668 = lo0018 & new_n1968 ;
  assign new_n14669 = ~lo0044 & lo0045 ;
  assign new_n14670 = new_n14668 & new_n14669 ;
  assign new_n14671 = lo0899 & ~new_n14670 ;
  assign new_n14672 = lo0054 & new_n14671 ;
  assign new_n14673 = lo0051 & ~new_n14672 ;
  assign new_n14674 = ~lo0051 & new_n14672 ;
  assign new_n14675 = ~new_n14673 & ~new_n14674 ;
  assign new_n14676 = lo0900 & ~lo0901 ;
  assign new_n14677 = ~new_n2246 & new_n14676 ;
  assign new_n14678 = lo0052 & ~lo0053 ;
  assign new_n14679 = ~lo0052 & lo0053 ;
  assign new_n14680 = ~new_n14678 & ~new_n14679 ;
  assign new_n14681 = new_n14677 & ~new_n14680 ;
  assign new_n14682 = lo0052 & ~new_n14677 ;
  assign new_n14683 = ~new_n14681 & ~new_n14682 ;
  assign new_n14684 = lo0053 & ~new_n14677 ;
  assign new_n14685 = ~lo0053 & new_n14677 ;
  assign new_n14686 = ~new_n14684 & ~new_n14685 ;
  assign new_n14687 = lo0054 & ~new_n14671 ;
  assign new_n14688 = ~lo0054 & new_n14671 ;
  assign new_n14689 = ~new_n14687 & ~new_n14688 ;
  assign new_n14690 = lo0055 & new_n2252 ;
  assign new_n14691 = ~new_n2252 & ~new_n13789 ;
  assign new_n14692 = ~new_n14690 & ~new_n14691 ;
  assign new_n14693 = lo0056 & new_n2252 ;
  assign new_n14694 = ~new_n2252 & new_n13808 ;
  assign new_n14695 = ~new_n14693 & ~new_n14694 ;
  assign new_n14696 = lo0057 & new_n2252 ;
  assign new_n14697 = lo0902 & ~new_n2252 ;
  assign new_n14698 = ~new_n14696 & ~new_n14697 ;
  assign new_n14699 = ~lo0017 & ~new_n2252 ;
  assign new_n14700 = lo0058 & ~new_n14699 ;
  assign new_n14701 = lo0903 & new_n14699 ;
  assign new_n14702 = ~new_n14700 & ~new_n14701 ;
  assign new_n14703 = lo0059 & ~new_n14699 ;
  assign new_n14704 = new_n13724 & new_n14699 ;
  assign new_n14705 = ~new_n14703 & ~new_n14704 ;
  assign new_n14706 = lo0060 & ~new_n14699 ;
  assign new_n14707 = lo0904 & new_n14699 ;
  assign new_n14708 = ~new_n14706 & ~new_n14707 ;
  assign new_n14709 = lo0061 & ~new_n14699 ;
  assign new_n14710 = new_n13736 & new_n14699 ;
  assign new_n14711 = ~new_n14709 & ~new_n14710 ;
  assign new_n14712 = lo0062 & ~new_n14699 ;
  assign new_n14713 = lo0905 & new_n14699 ;
  assign new_n14714 = ~new_n14712 & ~new_n14713 ;
  assign new_n14715 = lo0063 & ~new_n14699 ;
  assign new_n14716 = new_n13731 & new_n14699 ;
  assign new_n14717 = ~new_n14715 & ~new_n14716 ;
  assign new_n14718 = lo0064 & ~new_n14699 ;
  assign new_n14719 = lo0906 & new_n14699 ;
  assign new_n14720 = ~new_n14718 & ~new_n14719 ;
  assign new_n14721 = lo0065 & ~new_n14699 ;
  assign new_n14722 = new_n13763 & new_n14699 ;
  assign new_n14723 = ~new_n14721 & ~new_n14722 ;
  assign new_n14724 = lo0066 & new_n2252 ;
  assign new_n14725 = lo0907 & ~new_n2252 ;
  assign new_n14726 = ~new_n14724 & ~new_n14725 ;
  assign new_n14727 = lo0067 & new_n2252 ;
  assign new_n14728 = new_n12329 & ~new_n13810 ;
  assign new_n14729 = ~new_n12329 & ~new_n13798 ;
  assign new_n14730 = new_n13807 & ~new_n14729 ;
  assign new_n14731 = ~new_n14728 & new_n14730 ;
  assign new_n14732 = ~new_n2252 & new_n12523 ;
  assign new_n14733 = new_n14731 & new_n14732 ;
  assign new_n14734 = ~new_n14727 & ~new_n14733 ;
  assign new_n14735 = lo0068 & new_n2252 ;
  assign new_n14736 = ~new_n2264 & ~new_n12367 ;
  assign new_n14737 = new_n2465 & new_n12325 ;
  assign new_n14738 = ~new_n14736 & new_n14737 ;
  assign new_n14739 = ~new_n12329 & ~new_n12795 ;
  assign new_n14740 = ~new_n14738 & ~new_n14739 ;
  assign new_n14741 = ~new_n12357 & ~new_n14740 ;
  assign new_n14742 = new_n12368 & new_n13781 ;
  assign new_n14743 = ~new_n12329 & new_n14742 ;
  assign new_n14744 = new_n12329 & new_n12507 ;
  assign new_n14745 = ~new_n14737 & new_n14744 ;
  assign new_n14746 = ~new_n14743 & ~new_n14745 ;
  assign new_n14747 = ~new_n14741 & new_n14746 ;
  assign new_n14748 = new_n13562 & ~new_n14747 ;
  assign new_n14749 = ~lo0191 & ~new_n2264 ;
  assign new_n14750 = new_n2454 & ~new_n14749 ;
  assign new_n14751 = new_n13065 & new_n14750 ;
  assign new_n14752 = ~new_n12402 & ~new_n14751 ;
  assign new_n14753 = ~new_n14748 & new_n14752 ;
  assign new_n14754 = new_n2454 & ~new_n14753 ;
  assign new_n14755 = ~new_n2454 & new_n14753 ;
  assign new_n14756 = ~new_n14754 & ~new_n14755 ;
  assign new_n14757 = ~new_n2446 & ~new_n14756 ;
  assign new_n14758 = new_n2446 & new_n14754 ;
  assign new_n14759 = new_n12325 & new_n12860 ;
  assign new_n14760 = ~new_n12377 & ~new_n14759 ;
  assign new_n14761 = new_n12386 & ~new_n14760 ;
  assign new_n14762 = ~new_n2446 & ~new_n14761 ;
  assign new_n14763 = ~new_n12329 & ~new_n14762 ;
  assign new_n14764 = ~new_n12548 & ~new_n14763 ;
  assign new_n14765 = ~new_n2454 & ~new_n14764 ;
  assign new_n14766 = ~new_n14753 & new_n14765 ;
  assign new_n14767 = ~new_n14758 & ~new_n14766 ;
  assign new_n14768 = ~new_n14757 & new_n14767 ;
  assign new_n14769 = ~new_n2252 & ~new_n14768 ;
  assign new_n14770 = ~new_n14735 & ~new_n14769 ;
  assign new_n14771 = lo0069 & new_n2252 ;
  assign new_n14772 = ~new_n2450 & new_n12376 ;
  assign new_n14773 = ~new_n12689 & new_n14772 ;
  assign new_n14774 = new_n2450 & new_n12383 ;
  assign new_n14775 = new_n12536 & new_n14774 ;
  assign new_n14776 = ~new_n2450 & new_n12472 ;
  assign new_n14777 = ~new_n12682 & new_n14776 ;
  assign new_n14778 = ~new_n14775 & ~new_n14777 ;
  assign new_n14779 = new_n12325 & ~new_n14778 ;
  assign new_n14780 = ~new_n14773 & ~new_n14779 ;
  assign new_n14781 = ~new_n2252 & new_n12696 ;
  assign new_n14782 = ~new_n14780 & new_n14781 ;
  assign new_n14783 = ~new_n14771 & ~new_n14782 ;
  assign new_n14784 = lo0070 & new_n2252 ;
  assign new_n14785 = ~new_n12329 & ~new_n13768 ;
  assign new_n14786 = new_n12329 & ~new_n13798 ;
  assign new_n14787 = new_n13807 & ~new_n14786 ;
  assign new_n14788 = ~new_n14785 & new_n14787 ;
  assign new_n14789 = new_n12468 & new_n14788 ;
  assign new_n14790 = ~new_n2446 & new_n12695 ;
  assign new_n14791 = new_n2450 & new_n12955 ;
  assign new_n14792 = new_n2264 & new_n14791 ;
  assign new_n14793 = new_n12376 & new_n12683 ;
  assign new_n14794 = new_n12383 & ~new_n12689 ;
  assign new_n14795 = ~new_n14793 & ~new_n14794 ;
  assign new_n14796 = new_n12752 & ~new_n14795 ;
  assign new_n14797 = ~new_n14792 & ~new_n14796 ;
  assign new_n14798 = new_n14790 & ~new_n14797 ;
  assign new_n14799 = ~new_n14789 & ~new_n14798 ;
  assign new_n14800 = ~new_n2252 & ~new_n14799 ;
  assign new_n14801 = ~new_n14784 & ~new_n14800 ;
  assign new_n14802 = lo0071 & new_n2252 ;
  assign new_n14803 = new_n14732 & new_n14788 ;
  assign new_n14804 = ~new_n14802 & ~new_n14803 ;
  assign new_n14805 = lo0072 & new_n2252 ;
  assign new_n14806 = ~new_n2252 & new_n12468 ;
  assign new_n14807 = new_n14731 & new_n14806 ;
  assign new_n14808 = ~new_n14805 & ~new_n14807 ;
  assign new_n14809 = lo0073 & new_n2252 ;
  assign new_n14810 = new_n12580 & new_n12752 ;
  assign new_n14811 = new_n12376 & new_n14791 ;
  assign new_n14812 = ~new_n14810 & ~new_n14811 ;
  assign new_n14813 = new_n14790 & ~new_n14812 ;
  assign new_n14814 = ~new_n12467 & new_n14788 ;
  assign new_n14815 = ~new_n14813 & ~new_n14814 ;
  assign new_n14816 = ~new_n2252 & ~new_n14815 ;
  assign new_n14817 = ~new_n14809 & ~new_n14816 ;
  assign new_n14818 = lo0057 & ~lo0908 ;
  assign new_n14819 = lo0909 & ~lo0910 ;
  assign new_n14820 = lo0911 & new_n14819 ;
  assign new_n14821 = ~lo0912 & new_n14820 ;
  assign new_n14822 = lo0062 & ~lo0064 ;
  assign new_n14823 = lo0058 & new_n14822 ;
  assign new_n14824 = ~lo0060 & new_n14823 ;
  assign new_n14825 = ~lo0064 & lo0910 ;
  assign new_n14826 = lo0058 & ~lo0911 ;
  assign new_n14827 = ~new_n14825 & ~new_n14826 ;
  assign new_n14828 = ~lo0060 & lo0912 ;
  assign new_n14829 = lo0064 & ~lo0910 ;
  assign new_n14830 = ~new_n14828 & ~new_n14829 ;
  assign new_n14831 = new_n14827 & new_n14830 ;
  assign new_n14832 = lo0060 & ~lo0912 ;
  assign new_n14833 = ~lo0062 & lo0909 ;
  assign new_n14834 = ~new_n14832 & ~new_n14833 ;
  assign new_n14835 = ~lo0058 & lo0911 ;
  assign new_n14836 = lo0062 & ~lo0909 ;
  assign new_n14837 = ~new_n14835 & ~new_n14836 ;
  assign new_n14838 = new_n14834 & new_n14837 ;
  assign new_n14839 = new_n14831 & new_n14838 ;
  assign new_n14840 = ~lo0057 & lo0908 ;
  assign new_n14841 = ~new_n14839 & ~new_n14840 ;
  assign new_n14842 = new_n14824 & new_n14841 ;
  assign new_n14843 = ~new_n14821 & ~new_n14842 ;
  assign new_n14844 = lo0908 & ~new_n14843 ;
  assign new_n14845 = ~new_n14818 & ~new_n14844 ;
  assign new_n14846 = new_n14818 & ~new_n14824 ;
  assign new_n14847 = ~new_n2252 & ~new_n14846 ;
  assign new_n14848 = ~new_n14845 & new_n14847 ;
  assign new_n14849 = lo0074 & ~new_n14848 ;
  assign new_n14850 = lo0057 & lo0908 ;
  assign new_n14851 = ~new_n14839 & new_n14850 ;
  assign new_n14852 = ~new_n14821 & new_n14851 ;
  assign new_n14853 = ~new_n14818 & ~new_n14852 ;
  assign new_n14854 = ~new_n5455 & ~new_n14853 ;
  assign new_n14855 = ~new_n13936 & new_n14853 ;
  assign new_n14856 = ~new_n14854 & ~new_n14855 ;
  assign new_n14857 = new_n14848 & ~new_n14856 ;
  assign new_n14858 = ~new_n14849 & ~new_n14857 ;
  assign new_n14859 = ~lo0911 & new_n14819 ;
  assign new_n14860 = lo0912 & new_n14859 ;
  assign new_n14861 = ~lo0058 & new_n14822 ;
  assign new_n14862 = lo0060 & new_n14861 ;
  assign new_n14863 = new_n14841 & new_n14862 ;
  assign new_n14864 = ~new_n14860 & ~new_n14863 ;
  assign new_n14865 = lo0908 & ~new_n14864 ;
  assign new_n14866 = ~new_n14818 & ~new_n14865 ;
  assign new_n14867 = new_n14818 & ~new_n14862 ;
  assign new_n14868 = ~new_n2252 & ~new_n14867 ;
  assign new_n14869 = ~new_n14866 & new_n14868 ;
  assign new_n14870 = lo0075 & ~new_n14869 ;
  assign new_n14871 = new_n14851 & ~new_n14860 ;
  assign new_n14872 = ~new_n14818 & ~new_n14871 ;
  assign new_n14873 = ~new_n5455 & ~new_n14872 ;
  assign new_n14874 = ~new_n13936 & new_n14872 ;
  assign new_n14875 = ~new_n14873 & ~new_n14874 ;
  assign new_n14876 = new_n14869 & ~new_n14875 ;
  assign new_n14877 = ~new_n14870 & ~new_n14876 ;
  assign new_n14878 = ~lo0912 & new_n14859 ;
  assign new_n14879 = ~lo0060 & new_n14861 ;
  assign new_n14880 = new_n14841 & new_n14879 ;
  assign new_n14881 = ~new_n14878 & ~new_n14880 ;
  assign new_n14882 = lo0908 & ~new_n14881 ;
  assign new_n14883 = ~new_n14818 & ~new_n14882 ;
  assign new_n14884 = new_n14818 & ~new_n14879 ;
  assign new_n14885 = ~new_n2252 & ~new_n14884 ;
  assign new_n14886 = ~new_n14883 & new_n14885 ;
  assign new_n14887 = lo0076 & ~new_n14886 ;
  assign new_n14888 = new_n14851 & ~new_n14878 ;
  assign new_n14889 = ~new_n14818 & ~new_n14888 ;
  assign new_n14890 = ~new_n5455 & ~new_n14889 ;
  assign new_n14891 = ~new_n13936 & new_n14889 ;
  assign new_n14892 = ~new_n14890 & ~new_n14891 ;
  assign new_n14893 = new_n14886 & ~new_n14892 ;
  assign new_n14894 = ~new_n14887 & ~new_n14893 ;
  assign new_n14895 = lo0912 & new_n14820 ;
  assign new_n14896 = lo0060 & new_n14823 ;
  assign new_n14897 = new_n14841 & new_n14896 ;
  assign new_n14898 = ~new_n14895 & ~new_n14897 ;
  assign new_n14899 = lo0908 & ~new_n14898 ;
  assign new_n14900 = ~new_n14818 & ~new_n14899 ;
  assign new_n14901 = new_n14818 & ~new_n14896 ;
  assign new_n14902 = ~new_n2252 & ~new_n14901 ;
  assign new_n14903 = ~new_n14900 & new_n14902 ;
  assign new_n14904 = lo0077 & ~new_n14903 ;
  assign new_n14905 = new_n14851 & ~new_n14895 ;
  assign new_n14906 = ~new_n14818 & ~new_n14905 ;
  assign new_n14907 = ~new_n5455 & ~new_n14906 ;
  assign new_n14908 = ~new_n13936 & new_n14906 ;
  assign new_n14909 = ~new_n14907 & ~new_n14908 ;
  assign new_n14910 = new_n14903 & ~new_n14909 ;
  assign new_n14911 = ~new_n14904 & ~new_n14910 ;
  assign new_n14912 = ~lo0909 & lo0910 ;
  assign new_n14913 = ~lo0911 & new_n14912 ;
  assign new_n14914 = lo0912 & new_n14913 ;
  assign new_n14915 = ~lo0062 & lo0064 ;
  assign new_n14916 = ~lo0058 & new_n14915 ;
  assign new_n14917 = lo0060 & new_n14916 ;
  assign new_n14918 = new_n14841 & new_n14917 ;
  assign new_n14919 = ~new_n14914 & ~new_n14918 ;
  assign new_n14920 = lo0908 & ~new_n14919 ;
  assign new_n14921 = ~new_n14818 & ~new_n14920 ;
  assign new_n14922 = new_n14818 & ~new_n14917 ;
  assign new_n14923 = ~new_n2252 & ~new_n14922 ;
  assign new_n14924 = ~new_n14921 & new_n14923 ;
  assign new_n14925 = lo0078 & ~new_n14924 ;
  assign new_n14926 = new_n14851 & ~new_n14914 ;
  assign new_n14927 = ~new_n14818 & ~new_n14926 ;
  assign new_n14928 = ~new_n5455 & ~new_n14927 ;
  assign new_n14929 = ~new_n13936 & new_n14927 ;
  assign new_n14930 = ~new_n14928 & ~new_n14929 ;
  assign new_n14931 = new_n14924 & ~new_n14930 ;
  assign new_n14932 = ~new_n14925 & ~new_n14931 ;
  assign new_n14933 = lo0911 & new_n14912 ;
  assign new_n14934 = ~lo0912 & new_n14933 ;
  assign new_n14935 = lo0058 & new_n14915 ;
  assign new_n14936 = ~lo0060 & new_n14935 ;
  assign new_n14937 = new_n14841 & new_n14936 ;
  assign new_n14938 = ~new_n14934 & ~new_n14937 ;
  assign new_n14939 = lo0908 & ~new_n14938 ;
  assign new_n14940 = ~new_n14818 & ~new_n14939 ;
  assign new_n14941 = new_n14818 & ~new_n14936 ;
  assign new_n14942 = ~new_n2252 & ~new_n14941 ;
  assign new_n14943 = ~new_n14940 & new_n14942 ;
  assign new_n14944 = lo0079 & ~new_n14943 ;
  assign new_n14945 = new_n14851 & ~new_n14934 ;
  assign new_n14946 = ~new_n14818 & ~new_n14945 ;
  assign new_n14947 = ~new_n5455 & ~new_n14946 ;
  assign new_n14948 = ~new_n13936 & new_n14946 ;
  assign new_n14949 = ~new_n14947 & ~new_n14948 ;
  assign new_n14950 = new_n14943 & ~new_n14949 ;
  assign new_n14951 = ~new_n14944 & ~new_n14950 ;
  assign new_n14952 = ~lo0912 & new_n14913 ;
  assign new_n14953 = ~lo0060 & new_n14916 ;
  assign new_n14954 = new_n14841 & new_n14953 ;
  assign new_n14955 = ~new_n14952 & ~new_n14954 ;
  assign new_n14956 = lo0908 & ~new_n14955 ;
  assign new_n14957 = ~new_n14818 & ~new_n14956 ;
  assign new_n14958 = new_n14818 & ~new_n14953 ;
  assign new_n14959 = ~new_n2252 & ~new_n14958 ;
  assign new_n14960 = ~new_n14957 & new_n14959 ;
  assign new_n14961 = lo0080 & ~new_n14960 ;
  assign new_n14962 = new_n14851 & ~new_n14952 ;
  assign new_n14963 = ~new_n14818 & ~new_n14962 ;
  assign new_n14964 = ~new_n5455 & ~new_n14963 ;
  assign new_n14965 = ~new_n13936 & new_n14963 ;
  assign new_n14966 = ~new_n14964 & ~new_n14965 ;
  assign new_n14967 = new_n14960 & ~new_n14966 ;
  assign new_n14968 = ~new_n14961 & ~new_n14967 ;
  assign new_n14969 = lo0912 & new_n14933 ;
  assign new_n14970 = lo0060 & new_n14935 ;
  assign new_n14971 = new_n14841 & new_n14970 ;
  assign new_n14972 = ~new_n14969 & ~new_n14971 ;
  assign new_n14973 = lo0908 & ~new_n14972 ;
  assign new_n14974 = ~new_n14818 & ~new_n14973 ;
  assign new_n14975 = new_n14818 & ~new_n14970 ;
  assign new_n14976 = ~new_n2252 & ~new_n14975 ;
  assign new_n14977 = ~new_n14974 & new_n14976 ;
  assign new_n14978 = lo0081 & ~new_n14977 ;
  assign new_n14979 = new_n14851 & ~new_n14969 ;
  assign new_n14980 = ~new_n14818 & ~new_n14979 ;
  assign new_n14981 = ~new_n5455 & ~new_n14980 ;
  assign new_n14982 = ~new_n13936 & new_n14980 ;
  assign new_n14983 = ~new_n14981 & ~new_n14982 ;
  assign new_n14984 = new_n14977 & ~new_n14983 ;
  assign new_n14985 = ~new_n14978 & ~new_n14984 ;
  assign new_n14986 = ~lo0909 & ~lo0910 ;
  assign new_n14987 = lo0911 & new_n14986 ;
  assign new_n14988 = ~lo0912 & new_n14987 ;
  assign new_n14989 = lo0058 & new_n3122 ;
  assign new_n14990 = ~lo0060 & new_n14989 ;
  assign new_n14991 = new_n14841 & new_n14990 ;
  assign new_n14992 = ~new_n14988 & ~new_n14991 ;
  assign new_n14993 = lo0908 & ~new_n14992 ;
  assign new_n14994 = ~new_n14818 & ~new_n14993 ;
  assign new_n14995 = new_n14818 & ~new_n14990 ;
  assign new_n14996 = ~new_n2252 & ~new_n14995 ;
  assign new_n14997 = ~new_n14994 & new_n14996 ;
  assign new_n14998 = lo0082 & ~new_n14997 ;
  assign new_n14999 = new_n14851 & ~new_n14988 ;
  assign new_n15000 = ~new_n14818 & ~new_n14999 ;
  assign new_n15001 = ~new_n5455 & ~new_n15000 ;
  assign new_n15002 = ~new_n13936 & new_n15000 ;
  assign new_n15003 = ~new_n15001 & ~new_n15002 ;
  assign new_n15004 = new_n14997 & ~new_n15003 ;
  assign new_n15005 = ~new_n14998 & ~new_n15004 ;
  assign new_n15006 = ~lo0911 & new_n14986 ;
  assign new_n15007 = lo0912 & new_n15006 ;
  assign new_n15008 = ~lo0058 & new_n3122 ;
  assign new_n15009 = lo0060 & new_n15008 ;
  assign new_n15010 = new_n14841 & new_n15009 ;
  assign new_n15011 = ~new_n15007 & ~new_n15010 ;
  assign new_n15012 = lo0908 & ~new_n15011 ;
  assign new_n15013 = ~new_n14818 & ~new_n15012 ;
  assign new_n15014 = new_n14818 & ~new_n15009 ;
  assign new_n15015 = ~new_n2252 & ~new_n15014 ;
  assign new_n15016 = ~new_n15013 & new_n15015 ;
  assign new_n15017 = lo0083 & ~new_n15016 ;
  assign new_n15018 = new_n14851 & ~new_n15007 ;
  assign new_n15019 = ~new_n14818 & ~new_n15018 ;
  assign new_n15020 = ~new_n5455 & ~new_n15019 ;
  assign new_n15021 = ~new_n13936 & new_n15019 ;
  assign new_n15022 = ~new_n15020 & ~new_n15021 ;
  assign new_n15023 = new_n15016 & ~new_n15022 ;
  assign new_n15024 = ~new_n15017 & ~new_n15023 ;
  assign new_n15025 = ~lo0912 & new_n15006 ;
  assign new_n15026 = ~lo0060 & new_n15008 ;
  assign new_n15027 = new_n14841 & new_n15026 ;
  assign new_n15028 = ~new_n15025 & ~new_n15027 ;
  assign new_n15029 = lo0908 & ~new_n15028 ;
  assign new_n15030 = ~new_n14818 & ~new_n15029 ;
  assign new_n15031 = new_n14818 & ~new_n15026 ;
  assign new_n15032 = ~new_n2252 & ~new_n15031 ;
  assign new_n15033 = ~new_n15030 & new_n15032 ;
  assign new_n15034 = lo0084 & ~new_n15033 ;
  assign new_n15035 = new_n14851 & ~new_n15025 ;
  assign new_n15036 = ~new_n14818 & ~new_n15035 ;
  assign new_n15037 = ~new_n5455 & ~new_n15036 ;
  assign new_n15038 = ~new_n13936 & new_n15036 ;
  assign new_n15039 = ~new_n15037 & ~new_n15038 ;
  assign new_n15040 = new_n15033 & ~new_n15039 ;
  assign new_n15041 = ~new_n15034 & ~new_n15040 ;
  assign new_n15042 = lo0912 & new_n14987 ;
  assign new_n15043 = lo0060 & new_n14989 ;
  assign new_n15044 = new_n14841 & new_n15043 ;
  assign new_n15045 = ~new_n15042 & ~new_n15044 ;
  assign new_n15046 = lo0908 & ~new_n15045 ;
  assign new_n15047 = ~new_n14818 & ~new_n15046 ;
  assign new_n15048 = new_n14818 & ~new_n15043 ;
  assign new_n15049 = ~new_n2252 & ~new_n15048 ;
  assign new_n15050 = ~new_n15047 & new_n15049 ;
  assign new_n15051 = lo0085 & ~new_n15050 ;
  assign new_n15052 = new_n14851 & ~new_n15042 ;
  assign new_n15053 = ~new_n14818 & ~new_n15052 ;
  assign new_n15054 = ~new_n5455 & ~new_n15053 ;
  assign new_n15055 = ~new_n13936 & new_n15053 ;
  assign new_n15056 = ~new_n15054 & ~new_n15055 ;
  assign new_n15057 = new_n15050 & ~new_n15056 ;
  assign new_n15058 = ~new_n15051 & ~new_n15057 ;
  assign new_n15059 = lo0909 & lo0910 ;
  assign new_n15060 = ~lo0911 & new_n15059 ;
  assign new_n15061 = lo0912 & new_n15060 ;
  assign new_n15062 = lo0062 & lo0064 ;
  assign new_n15063 = ~lo0058 & new_n15062 ;
  assign new_n15064 = lo0060 & new_n15063 ;
  assign new_n15065 = new_n14841 & new_n15064 ;
  assign new_n15066 = ~new_n15061 & ~new_n15065 ;
  assign new_n15067 = lo0908 & ~new_n15066 ;
  assign new_n15068 = ~new_n14818 & ~new_n15067 ;
  assign new_n15069 = new_n14818 & ~new_n15064 ;
  assign new_n15070 = ~new_n2252 & ~new_n15069 ;
  assign new_n15071 = ~new_n15068 & new_n15070 ;
  assign new_n15072 = lo0086 & ~new_n15071 ;
  assign new_n15073 = new_n14851 & ~new_n15061 ;
  assign new_n15074 = ~new_n14818 & ~new_n15073 ;
  assign new_n15075 = ~new_n5455 & ~new_n15074 ;
  assign new_n15076 = ~new_n13936 & new_n15074 ;
  assign new_n15077 = ~new_n15075 & ~new_n15076 ;
  assign new_n15078 = new_n15071 & ~new_n15077 ;
  assign new_n15079 = ~new_n15072 & ~new_n15078 ;
  assign new_n15080 = lo0911 & new_n15059 ;
  assign new_n15081 = ~lo0912 & new_n15080 ;
  assign new_n15082 = lo0058 & new_n15062 ;
  assign new_n15083 = ~lo0060 & new_n15082 ;
  assign new_n15084 = new_n14841 & new_n15083 ;
  assign new_n15085 = ~new_n15081 & ~new_n15084 ;
  assign new_n15086 = lo0908 & ~new_n15085 ;
  assign new_n15087 = ~new_n14818 & ~new_n15086 ;
  assign new_n15088 = new_n14818 & ~new_n15083 ;
  assign new_n15089 = ~new_n2252 & ~new_n15088 ;
  assign new_n15090 = ~new_n15087 & new_n15089 ;
  assign new_n15091 = lo0087 & ~new_n15090 ;
  assign new_n15092 = new_n14851 & ~new_n15081 ;
  assign new_n15093 = ~new_n14818 & ~new_n15092 ;
  assign new_n15094 = ~new_n5455 & ~new_n15093 ;
  assign new_n15095 = ~new_n13936 & new_n15093 ;
  assign new_n15096 = ~new_n15094 & ~new_n15095 ;
  assign new_n15097 = new_n15090 & ~new_n15096 ;
  assign new_n15098 = ~new_n15091 & ~new_n15097 ;
  assign new_n15099 = ~lo0912 & new_n15060 ;
  assign new_n15100 = ~lo0060 & new_n15063 ;
  assign new_n15101 = new_n14841 & new_n15100 ;
  assign new_n15102 = ~new_n15099 & ~new_n15101 ;
  assign new_n15103 = lo0908 & ~new_n15102 ;
  assign new_n15104 = ~new_n14818 & ~new_n15103 ;
  assign new_n15105 = new_n14818 & ~new_n15100 ;
  assign new_n15106 = ~new_n2252 & ~new_n15105 ;
  assign new_n15107 = ~new_n15104 & new_n15106 ;
  assign new_n15108 = lo0088 & ~new_n15107 ;
  assign new_n15109 = new_n14851 & ~new_n15099 ;
  assign new_n15110 = ~new_n14818 & ~new_n15109 ;
  assign new_n15111 = ~new_n5455 & ~new_n15110 ;
  assign new_n15112 = ~new_n13936 & new_n15110 ;
  assign new_n15113 = ~new_n15111 & ~new_n15112 ;
  assign new_n15114 = new_n15107 & ~new_n15113 ;
  assign new_n15115 = ~new_n15108 & ~new_n15114 ;
  assign new_n15116 = lo0912 & new_n15080 ;
  assign new_n15117 = lo0060 & new_n15082 ;
  assign new_n15118 = new_n14841 & new_n15117 ;
  assign new_n15119 = ~new_n15116 & ~new_n15118 ;
  assign new_n15120 = lo0908 & ~new_n15119 ;
  assign new_n15121 = ~new_n14818 & ~new_n15120 ;
  assign new_n15122 = new_n14818 & ~new_n15117 ;
  assign new_n15123 = ~new_n2252 & ~new_n15122 ;
  assign new_n15124 = ~new_n15121 & new_n15123 ;
  assign new_n15125 = lo0089 & ~new_n15124 ;
  assign new_n15126 = new_n14851 & ~new_n15116 ;
  assign new_n15127 = ~new_n14818 & ~new_n15126 ;
  assign new_n15128 = ~new_n5455 & ~new_n15127 ;
  assign new_n15129 = ~new_n13936 & new_n15127 ;
  assign new_n15130 = ~new_n15128 & ~new_n15129 ;
  assign new_n15131 = new_n15124 & ~new_n15130 ;
  assign new_n15132 = ~new_n15125 & ~new_n15131 ;
  assign new_n15133 = lo0090 & new_n2252 ;
  assign new_n15134 = lo0913 & ~new_n2252 ;
  assign new_n15135 = ~new_n15133 & ~new_n15134 ;
  assign new_n15136 = ~lo0044 & lo0117 ;
  assign new_n15137 = ~new_n2249 & new_n15136 ;
  assign new_n15138 = lo0091 & ~new_n15137 ;
  assign new_n15139 = lo0914 & new_n15137 ;
  assign new_n15140 = ~new_n15138 & ~new_n15139 ;
  assign new_n15141 = lo0092 & ~new_n15137 ;
  assign new_n15142 = lo0893 & new_n15137 ;
  assign new_n15143 = ~new_n15141 & ~new_n15142 ;
  assign new_n15144 = lo0093 & ~new_n15137 ;
  assign new_n15145 = lo0915 & new_n15137 ;
  assign new_n15146 = ~new_n15144 & ~new_n15145 ;
  assign new_n15147 = lo0094 & ~new_n15137 ;
  assign new_n15148 = pi020 & new_n1982 ;
  assign new_n15149 = pi017 & new_n1973 ;
  assign new_n15150 = pi018 & new_n1976 ;
  assign new_n15151 = ~new_n15149 & ~new_n15150 ;
  assign new_n15152 = ~new_n15148 & new_n15151 ;
  assign new_n15153 = pi024 & new_n1991 ;
  assign new_n15154 = new_n1965 & new_n1970 ;
  assign new_n15155 = lo0917 & lo0918 ;
  assign new_n15156 = lo0182 & ~lo0917 ;
  assign new_n15157 = ~new_n15155 & ~new_n15156 ;
  assign new_n15158 = new_n15154 & ~new_n15157 ;
  assign new_n15159 = lo0916 & new_n14668 ;
  assign new_n15160 = ~new_n15158 & ~new_n15159 ;
  assign new_n15161 = ~new_n15153 & new_n15160 ;
  assign new_n15162 = pi021 & new_n1985 ;
  assign new_n15163 = pi022 & new_n1987 ;
  assign new_n15164 = ~new_n15162 & ~new_n15163 ;
  assign new_n15165 = pi019 & new_n1979 ;
  assign new_n15166 = pi023 & new_n1989 ;
  assign new_n15167 = ~new_n15165 & ~new_n15166 ;
  assign new_n15168 = new_n15164 & new_n15167 ;
  assign new_n15169 = new_n15161 & new_n15168 ;
  assign new_n15170 = new_n15152 & new_n15169 ;
  assign new_n15171 = new_n15137 & ~new_n15170 ;
  assign new_n15172 = ~new_n15147 & ~new_n15171 ;
  assign new_n15173 = lo0095 & ~new_n15137 ;
  assign new_n15174 = lo0892 & new_n15137 ;
  assign new_n15175 = ~new_n15173 & ~new_n15174 ;
  assign new_n15176 = lo0096 & ~new_n15137 ;
  assign new_n15177 = pi028 & new_n1989 ;
  assign new_n15178 = pi026 & new_n1979 ;
  assign new_n15179 = pi027 & new_n1987 ;
  assign new_n15180 = ~new_n15178 & ~new_n15179 ;
  assign new_n15181 = ~new_n15177 & new_n15180 ;
  assign new_n15182 = lo0917 & lo0919 ;
  assign new_n15183 = lo0860 & ~lo0917 ;
  assign new_n15184 = ~new_n15182 & ~new_n15183 ;
  assign new_n15185 = new_n15154 & ~new_n15184 ;
  assign new_n15186 = pi032 & new_n1991 ;
  assign new_n15187 = ~new_n15185 & ~new_n15186 ;
  assign new_n15188 = pi030 & new_n1976 ;
  assign new_n15189 = pi031 & new_n1982 ;
  assign new_n15190 = ~new_n15188 & ~new_n15189 ;
  assign new_n15191 = pi025 & new_n1973 ;
  assign new_n15192 = pi029 & new_n1985 ;
  assign new_n15193 = ~new_n15191 & ~new_n15192 ;
  assign new_n15194 = new_n15190 & new_n15193 ;
  assign new_n15195 = new_n15187 & new_n15194 ;
  assign new_n15196 = new_n15181 & new_n15195 ;
  assign new_n15197 = new_n15137 & ~new_n15196 ;
  assign new_n15198 = ~new_n15176 & ~new_n15197 ;
  assign new_n15199 = lo0097 & ~new_n15137 ;
  assign new_n15200 = pi037 & new_n1982 ;
  assign new_n15201 = pi033 & new_n1987 ;
  assign new_n15202 = pi034 & new_n1989 ;
  assign new_n15203 = ~new_n15201 & ~new_n15202 ;
  assign new_n15204 = ~new_n15200 & new_n15203 ;
  assign new_n15205 = pi040 & new_n1991 ;
  assign new_n15206 = lo0920 & new_n14668 ;
  assign new_n15207 = lo0917 & new_n15154 ;
  assign new_n15208 = lo0921 & new_n15207 ;
  assign new_n15209 = ~new_n15206 & ~new_n15208 ;
  assign new_n15210 = ~new_n15205 & new_n15209 ;
  assign new_n15211 = pi038 & new_n1985 ;
  assign new_n15212 = pi039 & new_n1973 ;
  assign new_n15213 = ~new_n15211 & ~new_n15212 ;
  assign new_n15214 = pi035 & new_n1976 ;
  assign new_n15215 = pi036 & new_n1979 ;
  assign new_n15216 = ~new_n15214 & ~new_n15215 ;
  assign new_n15217 = new_n15213 & new_n15216 ;
  assign new_n15218 = new_n15210 & new_n15217 ;
  assign new_n15219 = new_n15204 & new_n15218 ;
  assign new_n15220 = new_n15137 & ~new_n15219 ;
  assign new_n15221 = ~new_n15199 & ~new_n15220 ;
  assign new_n15222 = lo0098 & ~new_n15137 ;
  assign new_n15223 = pi041 & new_n1987 ;
  assign new_n15224 = pi042 & new_n1991 ;
  assign new_n15225 = pi048 & new_n1985 ;
  assign new_n15226 = ~new_n15224 & ~new_n15225 ;
  assign new_n15227 = ~new_n15223 & new_n15226 ;
  assign new_n15228 = pi047 & new_n1982 ;
  assign new_n15229 = lo0917 & lo0922 ;
  assign new_n15230 = ~lo0917 & ~lo1431 ;
  assign new_n15231 = ~new_n15229 & ~new_n15230 ;
  assign new_n15232 = new_n15154 & ~new_n15231 ;
  assign new_n15233 = pi001 & new_n2187 ;
  assign new_n15234 = ~lo0054 & lo0925 ;
  assign new_n15235 = ~lo0051 & new_n15234 ;
  assign new_n15236 = lo0051 & lo0054 ;
  assign new_n15237 = ~lo0054 & lo0924 ;
  assign new_n15238 = lo0051 & new_n15237 ;
  assign new_n15239 = ~new_n15236 & ~new_n15238 ;
  assign new_n15240 = ~new_n15235 & new_n15239 ;
  assign new_n15241 = ~lo0054 & ~new_n15240 ;
  assign new_n15242 = lo0054 & new_n15240 ;
  assign new_n15243 = ~new_n15241 & ~new_n15242 ;
  assign new_n15244 = lo0923 & ~new_n15243 ;
  assign new_n15245 = ~lo0923 & new_n15241 ;
  assign new_n15246 = lo0054 & lo0926 ;
  assign new_n15247 = ~new_n15240 & new_n15246 ;
  assign new_n15248 = ~new_n15245 & ~new_n15247 ;
  assign new_n15249 = ~new_n15244 & new_n15248 ;
  assign new_n15250 = new_n14668 & ~new_n15249 ;
  assign new_n15251 = ~new_n15233 & ~new_n15250 ;
  assign new_n15252 = ~new_n15232 & new_n15251 ;
  assign new_n15253 = ~new_n15228 & new_n15252 ;
  assign new_n15254 = pi044 & new_n1973 ;
  assign new_n15255 = pi045 & new_n1976 ;
  assign new_n15256 = ~new_n15254 & ~new_n15255 ;
  assign new_n15257 = pi043 & new_n1989 ;
  assign new_n15258 = pi046 & new_n1979 ;
  assign new_n15259 = ~new_n15257 & ~new_n15258 ;
  assign new_n15260 = new_n15256 & new_n15259 ;
  assign new_n15261 = new_n15253 & new_n15260 ;
  assign new_n15262 = new_n15227 & new_n15261 ;
  assign new_n15263 = new_n15137 & ~new_n15262 ;
  assign new_n15264 = ~new_n15222 & ~new_n15263 ;
  assign new_n15265 = lo0099 & ~new_n15137 ;
  assign new_n15266 = pi052 & new_n1989 ;
  assign new_n15267 = pi049 & new_n1982 ;
  assign new_n15268 = pi050 & new_n1985 ;
  assign new_n15269 = ~new_n15267 & ~new_n15268 ;
  assign new_n15270 = ~new_n15266 & new_n15269 ;
  assign new_n15271 = pi056 & new_n1991 ;
  assign new_n15272 = lo0917 & lo0927 ;
  assign new_n15273 = ~lo0917 & ~lo1432 ;
  assign new_n15274 = ~new_n15272 & ~new_n15273 ;
  assign new_n15275 = new_n15154 & ~new_n15274 ;
  assign new_n15276 = ~lo1285 & new_n2245 ;
  assign new_n15277 = new_n14668 & new_n15276 ;
  assign new_n15278 = ~new_n15275 & ~new_n15277 ;
  assign new_n15279 = ~new_n15271 & new_n15278 ;
  assign new_n15280 = pi053 & new_n1976 ;
  assign new_n15281 = pi054 & new_n1973 ;
  assign new_n15282 = ~new_n15280 & ~new_n15281 ;
  assign new_n15283 = pi051 & new_n1987 ;
  assign new_n15284 = pi055 & new_n1979 ;
  assign new_n15285 = ~new_n15283 & ~new_n15284 ;
  assign new_n15286 = new_n15282 & new_n15285 ;
  assign new_n15287 = new_n15279 & new_n15286 ;
  assign new_n15288 = new_n15270 & new_n15287 ;
  assign new_n15289 = new_n15137 & ~new_n15288 ;
  assign new_n15290 = ~new_n15265 & ~new_n15289 ;
  assign new_n15291 = lo0100 & ~new_n15137 ;
  assign new_n15292 = pi060 & new_n1982 ;
  assign new_n15293 = pi057 & new_n1973 ;
  assign new_n15294 = pi058 & new_n1976 ;
  assign new_n15295 = ~new_n15293 & ~new_n15294 ;
  assign new_n15296 = ~new_n15292 & new_n15295 ;
  assign new_n15297 = pi064 & new_n1991 ;
  assign new_n15298 = lo0917 & lo0929 ;
  assign new_n15299 = ~lo0917 & lo0930 ;
  assign new_n15300 = ~new_n15298 & ~new_n15299 ;
  assign new_n15301 = new_n15154 & ~new_n15300 ;
  assign new_n15302 = lo0928 & new_n14668 ;
  assign new_n15303 = ~new_n15301 & ~new_n15302 ;
  assign new_n15304 = ~new_n15297 & new_n15303 ;
  assign new_n15305 = pi061 & new_n1985 ;
  assign new_n15306 = pi062 & new_n1987 ;
  assign new_n15307 = ~new_n15305 & ~new_n15306 ;
  assign new_n15308 = pi059 & new_n1979 ;
  assign new_n15309 = pi063 & new_n1989 ;
  assign new_n15310 = ~new_n15308 & ~new_n15309 ;
  assign new_n15311 = new_n15307 & new_n15310 ;
  assign new_n15312 = new_n15304 & new_n15311 ;
  assign new_n15313 = new_n15296 & new_n15312 ;
  assign new_n15314 = new_n15137 & ~new_n15313 ;
  assign new_n15315 = ~new_n15291 & ~new_n15314 ;
  assign new_n15316 = lo0101 & new_n2252 ;
  assign new_n15317 = ~new_n2252 & ~new_n13324 ;
  assign new_n15318 = ~new_n15316 & ~new_n15317 ;
  assign new_n15319 = lo0102 & new_n2252 ;
  assign new_n15320 = new_n12325 & new_n12368 ;
  assign new_n15321 = new_n12376 & new_n15320 ;
  assign new_n15322 = ~new_n2465 & ~new_n15320 ;
  assign new_n15323 = ~new_n15321 & ~new_n15322 ;
  assign new_n15324 = new_n2455 & new_n12357 ;
  assign new_n15325 = ~new_n15323 & new_n15324 ;
  assign new_n15326 = ~new_n12580 & ~new_n14761 ;
  assign new_n15327 = new_n12402 & ~new_n15326 ;
  assign new_n15328 = ~new_n12404 & ~new_n15327 ;
  assign new_n15329 = ~new_n15325 & new_n15328 ;
  assign new_n15330 = ~new_n2252 & new_n12522 ;
  assign new_n15331 = ~new_n15329 & new_n15330 ;
  assign new_n15332 = ~new_n15319 & ~new_n15331 ;
  assign new_n15333 = lo0103 & new_n2252 ;
  assign new_n15334 = ~new_n12367 & new_n12591 ;
  assign new_n15335 = ~new_n12329 & ~new_n15334 ;
  assign new_n15336 = ~new_n2446 & new_n2450 ;
  assign new_n15337 = ~new_n2252 & new_n15336 ;
  assign new_n15338 = ~new_n13513 & new_n15337 ;
  assign new_n15339 = ~new_n15335 & new_n15338 ;
  assign new_n15340 = ~new_n15333 & ~new_n15339 ;
  assign new_n15341 = lo0104 & new_n2252 ;
  assign new_n15342 = ~new_n2252 & ~new_n13105 ;
  assign new_n15343 = ~new_n15341 & ~new_n15342 ;
  assign new_n15344 = lo0105 & new_n2252 ;
  assign new_n15345 = new_n12357 & new_n13286 ;
  assign new_n15346 = ~new_n12796 & ~new_n15345 ;
  assign new_n15347 = new_n2455 & new_n12522 ;
  assign new_n15348 = ~new_n2252 & new_n15347 ;
  assign new_n15349 = ~new_n15346 & new_n15348 ;
  assign new_n15350 = ~new_n15344 & ~new_n15349 ;
  assign new_n15351 = lo0106 & new_n2252 ;
  assign new_n15352 = new_n2455 & new_n13408 ;
  assign new_n15353 = ~new_n2252 & new_n12367 ;
  assign new_n15354 = new_n15352 & new_n15353 ;
  assign new_n15355 = ~new_n15351 & ~new_n15354 ;
  assign new_n15356 = lo0107 & new_n2252 ;
  assign new_n15357 = ~new_n2252 & ~new_n12367 ;
  assign new_n15358 = new_n15352 & new_n15357 ;
  assign new_n15359 = ~new_n15356 & ~new_n15358 ;
  assign new_n15360 = lo0108 & new_n2252 ;
  assign new_n15361 = ~new_n2252 & ~new_n2454 ;
  assign new_n15362 = new_n13429 & new_n15361 ;
  assign new_n15363 = ~new_n15360 & ~new_n15362 ;
  assign new_n15364 = ~lo0952 & ~lo0953 ;
  assign new_n15365 = ~new_n2252 & ~new_n15364 ;
  assign new_n15366 = lo0109 & ~new_n15365 ;
  assign new_n15367 = lo0952 & ~new_n13936 ;
  assign new_n15368 = ~lo0952 & ~new_n5455 ;
  assign new_n15369 = ~new_n15367 & ~new_n15368 ;
  assign new_n15370 = new_n15365 & ~new_n15369 ;
  assign new_n15371 = ~new_n15366 & ~new_n15370 ;
  assign new_n15372 = new_n12402 & new_n12522 ;
  assign new_n15373 = new_n12357 & new_n15372 ;
  assign new_n15374 = new_n12383 & new_n12395 ;
  assign new_n15375 = new_n15373 & new_n15374 ;
  assign new_n15376 = ~new_n2252 & ~new_n15375 ;
  assign new_n15377 = lo0110 & ~new_n15376 ;
  assign new_n15378 = lo0854 & ~new_n10220 ;
  assign new_n15379 = lo0855 & ~new_n2739 ;
  assign new_n15380 = ~lo0855 & ~lo0957 ;
  assign new_n15381 = lo0858 & ~new_n5455 ;
  assign new_n15382 = lo0859 & ~new_n13936 ;
  assign new_n15383 = lo0110 & ~lo0859 ;
  assign new_n15384 = ~new_n15382 & ~new_n15383 ;
  assign new_n15385 = ~lo0858 & ~new_n15384 ;
  assign new_n15386 = ~new_n15381 & ~new_n15385 ;
  assign new_n15387 = new_n15380 & ~new_n15386 ;
  assign new_n15388 = ~new_n15379 & ~new_n15387 ;
  assign new_n15389 = ~lo0854 & ~new_n15388 ;
  assign new_n15390 = ~new_n15378 & ~new_n15389 ;
  assign new_n15391 = new_n15376 & ~new_n15390 ;
  assign new_n15392 = ~new_n15377 & ~new_n15391 ;
  assign new_n15393 = lo0958 & ~new_n2252 ;
  assign new_n15394 = new_n12460 & ~new_n13536 ;
  assign new_n15395 = ~new_n12460 & ~new_n12482 ;
  assign new_n15396 = ~new_n15394 & ~new_n15395 ;
  assign new_n15397 = ~new_n12420 & ~new_n15396 ;
  assign new_n15398 = new_n12460 & new_n13864 ;
  assign new_n15399 = ~new_n12442 & ~new_n12460 ;
  assign new_n15400 = ~new_n13865 & ~new_n15399 ;
  assign new_n15401 = ~new_n15398 & new_n15400 ;
  assign new_n15402 = ~new_n15397 & new_n15401 ;
  assign new_n15403 = new_n12486 & ~new_n15402 ;
  assign new_n15404 = ~new_n12420 & ~new_n12592 ;
  assign new_n15405 = new_n2264 & ~new_n15404 ;
  assign new_n15406 = ~new_n12460 & new_n12473 ;
  assign new_n15407 = new_n12442 & ~new_n15406 ;
  assign new_n15408 = ~new_n15405 & new_n15407 ;
  assign new_n15409 = new_n12477 & ~new_n15408 ;
  assign new_n15410 = ~new_n12479 & ~new_n15409 ;
  assign new_n15411 = ~new_n15403 & new_n15410 ;
  assign new_n15412 = new_n12452 & ~new_n15411 ;
  assign new_n15413 = ~new_n12452 & new_n15411 ;
  assign new_n15414 = ~new_n15412 & ~new_n15413 ;
  assign new_n15415 = ~new_n12444 & ~new_n15414 ;
  assign new_n15416 = new_n12444 & new_n15412 ;
  assign new_n15417 = new_n12499 & ~new_n15411 ;
  assign new_n15418 = new_n2450 & ~new_n15417 ;
  assign new_n15419 = ~new_n15416 & new_n15418 ;
  assign new_n15420 = ~new_n15415 & new_n15419 ;
  assign new_n15421 = new_n2446 & ~new_n15420 ;
  assign new_n15422 = ~new_n12386 & new_n13888 ;
  assign new_n15423 = new_n12325 & new_n12392 ;
  assign new_n15424 = new_n12395 & new_n12916 ;
  assign new_n15425 = ~new_n15423 & ~new_n15424 ;
  assign new_n15426 = new_n12357 & ~new_n15425 ;
  assign new_n15427 = ~new_n15422 & ~new_n15426 ;
  assign new_n15428 = ~new_n12329 & ~new_n15427 ;
  assign new_n15429 = ~new_n2450 & ~new_n12547 ;
  assign new_n15430 = ~new_n15428 & new_n15429 ;
  assign new_n15431 = ~new_n2454 & ~new_n15430 ;
  assign new_n15432 = ~new_n2263 & ~new_n12357 ;
  assign new_n15433 = new_n12325 & ~new_n15432 ;
  assign new_n15434 = ~lo0192 & ~new_n12325 ;
  assign new_n15435 = ~new_n12367 & ~new_n15434 ;
  assign new_n15436 = ~new_n15433 & new_n15435 ;
  assign new_n15437 = new_n12329 & ~new_n15436 ;
  assign new_n15438 = new_n12620 & ~new_n12917 ;
  assign new_n15439 = ~new_n12329 & ~new_n15438 ;
  assign new_n15440 = ~new_n15437 & ~new_n15439 ;
  assign new_n15441 = new_n15336 & ~new_n15440 ;
  assign new_n15442 = new_n2264 & new_n12590 ;
  assign new_n15443 = ~new_n12325 & new_n15442 ;
  assign new_n15444 = ~new_n2450 & ~new_n14749 ;
  assign new_n15445 = ~new_n15443 & ~new_n15444 ;
  assign new_n15446 = new_n2454 & ~new_n15445 ;
  assign new_n15447 = ~new_n15441 & ~new_n15446 ;
  assign new_n15448 = ~new_n15431 & new_n15447 ;
  assign new_n15449 = ~new_n15421 & new_n15448 ;
  assign new_n15450 = ~new_n2261 & new_n13926 ;
  assign new_n15451 = new_n13850 & ~new_n15450 ;
  assign new_n15452 = ~new_n2252 & new_n15451 ;
  assign new_n15453 = ~new_n15449 & new_n15452 ;
  assign new_n15454 = ~new_n15393 & ~new_n15453 ;
  assign new_n15455 = lo0111 & new_n15454 ;
  assign new_n15456 = lo0958 & ~new_n13936 ;
  assign new_n15457 = ~lo0958 & ~new_n13952 ;
  assign new_n15458 = ~new_n15456 & ~new_n15457 ;
  assign new_n15459 = ~new_n15454 & ~new_n15458 ;
  assign new_n15460 = ~new_n15455 & ~new_n15459 ;
  assign new_n15461 = lo0112 & new_n2252 ;
  assign new_n15462 = new_n2454 & new_n13414 ;
  assign new_n15463 = ~new_n13829 & new_n15462 ;
  assign new_n15464 = new_n12471 & new_n12573 ;
  assign new_n15465 = ~new_n13082 & ~new_n15464 ;
  assign new_n15466 = new_n13406 & ~new_n15465 ;
  assign new_n15467 = ~new_n15463 & ~new_n15466 ;
  assign new_n15468 = new_n2446 & ~new_n2454 ;
  assign new_n15469 = ~new_n12800 & ~new_n15468 ;
  assign new_n15470 = ~new_n2450 & new_n15469 ;
  assign new_n15471 = ~new_n15467 & new_n15470 ;
  assign new_n15472 = new_n12508 & new_n13053 ;
  assign new_n15473 = ~new_n12522 & ~new_n15472 ;
  assign new_n15474 = new_n12527 & ~new_n12604 ;
  assign new_n15475 = new_n15473 & ~new_n15474 ;
  assign new_n15476 = new_n2446 & ~new_n15475 ;
  assign new_n15477 = ~new_n2446 & new_n15475 ;
  assign new_n15478 = ~new_n15476 & ~new_n15477 ;
  assign new_n15479 = new_n13776 & ~new_n15478 ;
  assign new_n15480 = ~new_n13776 & new_n15476 ;
  assign new_n15481 = ~new_n2456 & new_n12368 ;
  assign new_n15482 = ~new_n2446 & new_n12358 ;
  assign new_n15483 = ~new_n15481 & new_n15482 ;
  assign new_n15484 = ~new_n15475 & new_n15483 ;
  assign new_n15485 = ~new_n15480 & ~new_n15484 ;
  assign new_n15486 = ~new_n15479 & new_n15485 ;
  assign new_n15487 = new_n2454 & ~new_n15486 ;
  assign new_n15488 = ~new_n13775 & ~new_n15487 ;
  assign new_n15489 = new_n2450 & ~new_n15488 ;
  assign new_n15490 = ~new_n15471 & ~new_n15489 ;
  assign new_n15491 = ~new_n2252 & ~new_n15490 ;
  assign new_n15492 = new_n15451 & new_n15491 ;
  assign new_n15493 = ~new_n15461 & ~new_n15492 ;
  assign new_n15494 = lo0113 & new_n2252 ;
  assign new_n15495 = ~new_n12441 & ~new_n12442 ;
  assign new_n15496 = ~new_n12593 & ~new_n15495 ;
  assign new_n15497 = ~new_n12452 & ~new_n15496 ;
  assign new_n15498 = ~new_n12595 & ~new_n15497 ;
  assign new_n15499 = new_n12508 & ~new_n15498 ;
  assign new_n15500 = new_n2446 & new_n12605 ;
  assign new_n15501 = new_n12367 & new_n12395 ;
  assign new_n15502 = new_n12334 & new_n12368 ;
  assign new_n15503 = ~new_n2465 & ~new_n12368 ;
  assign new_n15504 = ~new_n15502 & ~new_n15503 ;
  assign new_n15505 = new_n12325 & ~new_n15504 ;
  assign new_n15506 = ~new_n15501 & ~new_n15505 ;
  assign new_n15507 = ~new_n2446 & new_n12357 ;
  assign new_n15508 = ~new_n15506 & new_n15507 ;
  assign new_n15509 = ~new_n15500 & ~new_n15508 ;
  assign new_n15510 = ~new_n12329 & ~new_n15509 ;
  assign new_n15511 = ~new_n15499 & ~new_n15510 ;
  assign new_n15512 = new_n2455 & ~new_n15511 ;
  assign new_n15513 = new_n12442 & ~new_n12477 ;
  assign new_n15514 = new_n2446 & new_n12420 ;
  assign new_n15515 = ~new_n15513 & new_n15514 ;
  assign new_n15516 = new_n12405 & ~new_n12441 ;
  assign new_n15517 = new_n15515 & new_n15516 ;
  assign new_n15518 = ~new_n12402 & ~new_n15517 ;
  assign new_n15519 = ~new_n15512 & new_n15518 ;
  assign new_n15520 = new_n2454 & ~new_n15519 ;
  assign new_n15521 = ~new_n2454 & new_n15519 ;
  assign new_n15522 = ~new_n15520 & ~new_n15521 ;
  assign new_n15523 = ~new_n12590 & ~new_n15522 ;
  assign new_n15524 = new_n12590 & new_n15520 ;
  assign new_n15525 = ~lo1292 & ~new_n12338 ;
  assign new_n15526 = new_n2262 & ~new_n15525 ;
  assign new_n15527 = ~new_n12689 & new_n15526 ;
  assign new_n15528 = ~lo1292 & ~new_n12912 ;
  assign new_n15529 = ~new_n12823 & ~new_n15528 ;
  assign new_n15530 = ~lo1294 & ~new_n15529 ;
  assign new_n15531 = new_n12325 & new_n15530 ;
  assign new_n15532 = new_n12471 & new_n13781 ;
  assign new_n15533 = ~new_n15531 & ~new_n15532 ;
  assign new_n15534 = ~new_n12682 & ~new_n15533 ;
  assign new_n15535 = ~new_n15527 & ~new_n15534 ;
  assign new_n15536 = new_n12522 & ~new_n15535 ;
  assign new_n15537 = ~new_n2454 & new_n15536 ;
  assign new_n15538 = ~new_n15519 & new_n15537 ;
  assign new_n15539 = ~new_n15524 & ~new_n15538 ;
  assign new_n15540 = ~new_n15523 & new_n15539 ;
  assign new_n15541 = ~new_n2252 & ~new_n15540 ;
  assign new_n15542 = ~new_n15494 & ~new_n15541 ;
  assign new_n15543 = lo0114 & new_n2252 ;
  assign new_n15544 = new_n12329 & ~new_n13829 ;
  assign new_n15545 = ~new_n12329 & ~new_n12442 ;
  assign new_n15546 = ~new_n15544 & ~new_n15545 ;
  assign new_n15547 = new_n12420 & ~new_n12429 ;
  assign new_n15548 = new_n12646 & new_n15547 ;
  assign new_n15549 = ~new_n15546 & new_n15548 ;
  assign new_n15550 = ~new_n12429 & new_n12508 ;
  assign new_n15551 = new_n12840 & new_n15550 ;
  assign new_n15552 = new_n12526 & new_n12596 ;
  assign new_n15553 = new_n13829 & new_n15552 ;
  assign new_n15554 = ~new_n12522 & ~new_n15553 ;
  assign new_n15555 = ~new_n15551 & new_n15554 ;
  assign new_n15556 = ~new_n2446 & ~new_n12367 ;
  assign new_n15557 = new_n12591 & new_n15556 ;
  assign new_n15558 = ~new_n2446 & ~new_n15557 ;
  assign new_n15559 = ~new_n15555 & ~new_n15558 ;
  assign new_n15560 = ~new_n2446 & new_n15334 ;
  assign new_n15561 = new_n15555 & new_n15560 ;
  assign new_n15562 = ~new_n15559 & ~new_n15561 ;
  assign new_n15563 = new_n2454 & ~new_n15562 ;
  assign new_n15564 = ~new_n2454 & new_n12590 ;
  assign new_n15565 = ~new_n15563 & ~new_n15564 ;
  assign new_n15566 = new_n2450 & ~new_n15565 ;
  assign new_n15567 = ~new_n15549 & ~new_n15566 ;
  assign new_n15568 = ~new_n2252 & ~new_n15567 ;
  assign new_n15569 = ~new_n15543 & ~new_n15568 ;
  assign new_n15570 = lo0115 & ~lo0116 ;
  assign new_n15571 = ~lo0115 & lo0116 ;
  assign new_n15572 = ~new_n15570 & ~new_n15571 ;
  assign new_n15573 = lo0018 & lo0022 ;
  assign new_n15574 = ~lo0115 & ~new_n15573 ;
  assign new_n15575 = ~lo0116 & ~new_n15574 ;
  assign new_n15576 = lo0120 & new_n2252 ;
  assign new_n15577 = new_n2263 & new_n12442 ;
  assign new_n15578 = new_n12606 & new_n15577 ;
  assign new_n15579 = new_n2456 & new_n13829 ;
  assign new_n15580 = ~new_n15578 & ~new_n15579 ;
  assign new_n15581 = ~new_n12420 & ~new_n15580 ;
  assign new_n15582 = ~new_n12605 & ~new_n15581 ;
  assign new_n15583 = new_n12526 & ~new_n15582 ;
  assign new_n15584 = new_n12601 & ~new_n15583 ;
  assign new_n15585 = new_n2446 & ~new_n15584 ;
  assign new_n15586 = ~new_n2446 & new_n15584 ;
  assign new_n15587 = ~new_n15585 & ~new_n15586 ;
  assign new_n15588 = new_n12591 & ~new_n15587 ;
  assign new_n15589 = ~new_n12591 & new_n15585 ;
  assign new_n15590 = ~new_n12334 & new_n12368 ;
  assign new_n15591 = new_n12358 & ~new_n15590 ;
  assign new_n15592 = lo1291 & new_n13286 ;
  assign new_n15593 = new_n2263 & ~new_n12357 ;
  assign new_n15594 = ~new_n15592 & new_n15593 ;
  assign new_n15595 = ~new_n12863 & ~new_n15594 ;
  assign new_n15596 = ~new_n12325 & ~new_n15595 ;
  assign new_n15597 = ~new_n15591 & ~new_n15596 ;
  assign new_n15598 = ~new_n2446 & ~new_n15597 ;
  assign new_n15599 = ~new_n15584 & new_n15598 ;
  assign new_n15600 = ~new_n15589 & ~new_n15599 ;
  assign new_n15601 = ~new_n15588 & new_n15600 ;
  assign new_n15602 = new_n2450 & ~new_n15601 ;
  assign new_n15603 = ~new_n2450 & ~new_n15536 ;
  assign new_n15604 = ~new_n2454 & ~new_n15603 ;
  assign new_n15605 = new_n12405 & new_n15515 ;
  assign new_n15606 = ~new_n15604 & ~new_n15605 ;
  assign new_n15607 = ~new_n15602 & new_n15606 ;
  assign new_n15608 = ~new_n2252 & ~new_n15607 ;
  assign new_n15609 = new_n15451 & new_n15608 ;
  assign new_n15610 = ~new_n15576 & ~new_n15609 ;
  assign new_n15611 = ~new_n2252 & new_n2264 ;
  assign new_n15612 = ~lo0122 & new_n15611 ;
  assign new_n15613 = lo0121 & ~new_n15612 ;
  assign new_n15614 = ~new_n2444 & new_n15612 ;
  assign new_n15615 = ~new_n15613 & ~new_n15614 ;
  assign new_n15616 = lo0122 & new_n2252 ;
  assign new_n15617 = ~new_n2252 & ~new_n15451 ;
  assign new_n15618 = ~new_n15616 & ~new_n15617 ;
  assign new_n15619 = lo0117 & ~lo0118 ;
  assign new_n15620 = lo0119 & ~new_n15619 ;
  assign new_n15621 = ~new_n2252 & new_n15620 ;
  assign new_n15622 = lo0123 & ~new_n15621 ;
  assign new_n15623 = lo0963 & new_n15621 ;
  assign new_n15624 = ~new_n15622 & ~new_n15623 ;
  assign new_n15625 = lo0124 & ~new_n15621 ;
  assign new_n15626 = lo0118 & new_n15621 ;
  assign new_n15627 = ~new_n15625 & ~new_n15626 ;
  assign new_n15628 = lo0125 & ~new_n15621 ;
  assign new_n15629 = lo0117 & new_n15621 ;
  assign new_n15630 = ~new_n15628 & ~new_n15629 ;
  assign new_n15631 = lo0126 & ~new_n15621 ;
  assign new_n15632 = lo0893 & new_n15621 ;
  assign new_n15633 = ~new_n15631 & ~new_n15632 ;
  assign new_n15634 = lo0127 & ~new_n15621 ;
  assign new_n15635 = ~new_n15196 & new_n15621 ;
  assign new_n15636 = ~new_n15634 & ~new_n15635 ;
  assign new_n15637 = lo0128 & ~new_n15621 ;
  assign new_n15638 = ~new_n15219 & new_n15621 ;
  assign new_n15639 = ~new_n15637 & ~new_n15638 ;
  assign new_n15640 = ~new_n2450 & new_n13896 ;
  assign new_n15641 = new_n12383 & ~new_n12508 ;
  assign new_n15642 = new_n12508 & new_n13872 ;
  assign new_n15643 = ~new_n15641 & ~new_n15642 ;
  assign new_n15644 = ~new_n12357 & new_n12590 ;
  assign new_n15645 = ~new_n12325 & ~new_n12367 ;
  assign new_n15646 = new_n15644 & new_n15645 ;
  assign new_n15647 = ~new_n13880 & ~new_n15646 ;
  assign new_n15648 = new_n2455 & ~new_n15647 ;
  assign new_n15649 = ~new_n15643 & new_n15648 ;
  assign new_n15650 = ~new_n15640 & ~new_n15649 ;
  assign new_n15651 = new_n15452 & ~new_n15650 ;
  assign new_n15652 = lo0129 & ~new_n15452 ;
  assign new_n15653 = ~new_n15651 & ~new_n15652 ;
  assign new_n15654 = lo0130 & ~new_n15621 ;
  assign new_n15655 = lo0964 & new_n15621 ;
  assign new_n15656 = ~new_n15654 & ~new_n15655 ;
  assign new_n15657 = lo0131 & ~new_n15621 ;
  assign new_n15658 = pi065 & new_n1987 ;
  assign new_n15659 = pi066 & new_n1991 ;
  assign new_n15660 = pi072 & new_n1985 ;
  assign new_n15661 = ~new_n15659 & ~new_n15660 ;
  assign new_n15662 = ~new_n15658 & new_n15661 ;
  assign new_n15663 = pi071 & new_n1982 ;
  assign new_n15664 = lo0917 & lo0965 ;
  assign new_n15665 = ~lo0917 & ~lo1433 ;
  assign new_n15666 = ~new_n15664 & ~new_n15665 ;
  assign new_n15667 = new_n15154 & ~new_n15666 ;
  assign new_n15668 = pi002 & new_n2187 ;
  assign new_n15669 = ~lo0054 & lo0968 ;
  assign new_n15670 = ~lo0051 & new_n15669 ;
  assign new_n15671 = ~lo0054 & lo0967 ;
  assign new_n15672 = lo0051 & new_n15671 ;
  assign new_n15673 = ~new_n15236 & ~new_n15672 ;
  assign new_n15674 = ~new_n15670 & new_n15673 ;
  assign new_n15675 = ~lo0054 & ~new_n15674 ;
  assign new_n15676 = lo0054 & new_n15674 ;
  assign new_n15677 = ~new_n15675 & ~new_n15676 ;
  assign new_n15678 = lo0966 & ~new_n15677 ;
  assign new_n15679 = ~lo0966 & new_n15675 ;
  assign new_n15680 = lo0054 & lo0969 ;
  assign new_n15681 = ~new_n15674 & new_n15680 ;
  assign new_n15682 = ~new_n15679 & ~new_n15681 ;
  assign new_n15683 = ~new_n15678 & new_n15682 ;
  assign new_n15684 = new_n14668 & ~new_n15683 ;
  assign new_n15685 = ~new_n15668 & ~new_n15684 ;
  assign new_n15686 = ~new_n15667 & new_n15685 ;
  assign new_n15687 = ~new_n15663 & new_n15686 ;
  assign new_n15688 = pi068 & new_n1973 ;
  assign new_n15689 = pi069 & new_n1976 ;
  assign new_n15690 = ~new_n15688 & ~new_n15689 ;
  assign new_n15691 = pi067 & new_n1989 ;
  assign new_n15692 = pi070 & new_n1979 ;
  assign new_n15693 = ~new_n15691 & ~new_n15692 ;
  assign new_n15694 = new_n15690 & new_n15693 ;
  assign new_n15695 = new_n15687 & new_n15694 ;
  assign new_n15696 = new_n15662 & new_n15695 ;
  assign new_n15697 = new_n15621 & ~new_n15696 ;
  assign new_n15698 = ~new_n15657 & ~new_n15697 ;
  assign new_n15699 = lo0132 & ~new_n15621 ;
  assign new_n15700 = pi073 & new_n1987 ;
  assign new_n15701 = pi074 & new_n1991 ;
  assign new_n15702 = pi080 & new_n1985 ;
  assign new_n15703 = ~new_n15701 & ~new_n15702 ;
  assign new_n15704 = ~new_n15700 & new_n15703 ;
  assign new_n15705 = pi079 & new_n1982 ;
  assign new_n15706 = lo0917 & lo0970 ;
  assign new_n15707 = lo0878 & ~lo0917 ;
  assign new_n15708 = ~new_n15706 & ~new_n15707 ;
  assign new_n15709 = new_n15154 & ~new_n15708 ;
  assign new_n15710 = pi003 & new_n2187 ;
  assign new_n15711 = lo0971 & new_n14668 ;
  assign new_n15712 = ~new_n15710 & ~new_n15711 ;
  assign new_n15713 = ~new_n15709 & new_n15712 ;
  assign new_n15714 = ~new_n15705 & new_n15713 ;
  assign new_n15715 = pi076 & new_n1973 ;
  assign new_n15716 = pi077 & new_n1976 ;
  assign new_n15717 = ~new_n15715 & ~new_n15716 ;
  assign new_n15718 = pi075 & new_n1989 ;
  assign new_n15719 = pi078 & new_n1979 ;
  assign new_n15720 = ~new_n15718 & ~new_n15719 ;
  assign new_n15721 = new_n15717 & new_n15720 ;
  assign new_n15722 = new_n15714 & new_n15721 ;
  assign new_n15723 = new_n15704 & new_n15722 ;
  assign new_n15724 = new_n15621 & ~new_n15723 ;
  assign new_n15725 = ~new_n15699 & ~new_n15724 ;
  assign new_n15726 = lo0133 & ~new_n15621 ;
  assign new_n15727 = lo0972 & new_n15621 ;
  assign new_n15728 = ~new_n15726 & ~new_n15727 ;
  assign new_n15729 = lo0134 & ~new_n15621 ;
  assign new_n15730 = pi084 & new_n1989 ;
  assign new_n15731 = pi082 & new_n1979 ;
  assign new_n15732 = pi083 & new_n1987 ;
  assign new_n15733 = ~new_n15731 & ~new_n15732 ;
  assign new_n15734 = ~new_n15730 & new_n15733 ;
  assign new_n15735 = lo0917 & lo0973 ;
  assign new_n15736 = lo0866 & ~lo0917 ;
  assign new_n15737 = ~new_n15735 & ~new_n15736 ;
  assign new_n15738 = new_n15154 & ~new_n15737 ;
  assign new_n15739 = pi088 & new_n1991 ;
  assign new_n15740 = ~new_n15738 & ~new_n15739 ;
  assign new_n15741 = pi086 & new_n1976 ;
  assign new_n15742 = pi087 & new_n1982 ;
  assign new_n15743 = ~new_n15741 & ~new_n15742 ;
  assign new_n15744 = pi081 & new_n1973 ;
  assign new_n15745 = pi085 & new_n1985 ;
  assign new_n15746 = ~new_n15744 & ~new_n15745 ;
  assign new_n15747 = new_n15743 & new_n15746 ;
  assign new_n15748 = new_n15740 & new_n15747 ;
  assign new_n15749 = new_n15734 & new_n15748 ;
  assign new_n15750 = new_n15621 & ~new_n15749 ;
  assign new_n15751 = ~new_n15729 & ~new_n15750 ;
  assign new_n15752 = lo0135 & ~new_n15621 ;
  assign new_n15753 = pi093 & new_n1982 ;
  assign new_n15754 = pi089 & new_n1987 ;
  assign new_n15755 = pi090 & new_n1989 ;
  assign new_n15756 = ~new_n15754 & ~new_n15755 ;
  assign new_n15757 = ~new_n15753 & new_n15756 ;
  assign new_n15758 = pi096 & new_n1991 ;
  assign new_n15759 = lo0974 & new_n14668 ;
  assign new_n15760 = lo0975 & new_n15207 ;
  assign new_n15761 = ~new_n15759 & ~new_n15760 ;
  assign new_n15762 = ~new_n15758 & new_n15761 ;
  assign new_n15763 = pi094 & new_n1985 ;
  assign new_n15764 = pi095 & new_n1973 ;
  assign new_n15765 = ~new_n15763 & ~new_n15764 ;
  assign new_n15766 = pi091 & new_n1976 ;
  assign new_n15767 = pi092 & new_n1979 ;
  assign new_n15768 = ~new_n15766 & ~new_n15767 ;
  assign new_n15769 = new_n15765 & new_n15768 ;
  assign new_n15770 = new_n15762 & new_n15769 ;
  assign new_n15771 = new_n15757 & new_n15770 ;
  assign new_n15772 = new_n15621 & ~new_n15771 ;
  assign new_n15773 = ~new_n15752 & ~new_n15772 ;
  assign new_n15774 = lo0136 & ~new_n15621 ;
  assign new_n15775 = lo0976 & new_n15621 ;
  assign new_n15776 = ~new_n15774 & ~new_n15775 ;
  assign new_n15777 = lo0137 & ~new_n15621 ;
  assign new_n15778 = pi100 & new_n1982 ;
  assign new_n15779 = pi097 & new_n1973 ;
  assign new_n15780 = pi098 & new_n1976 ;
  assign new_n15781 = ~new_n15779 & ~new_n15780 ;
  assign new_n15782 = ~new_n15778 & new_n15781 ;
  assign new_n15783 = pi104 & new_n1991 ;
  assign new_n15784 = lo0917 & lo0981 ;
  assign new_n15785 = ~lo0917 & ~lo1435 ;
  assign new_n15786 = ~new_n15784 & ~new_n15785 ;
  assign new_n15787 = new_n15154 & ~new_n15786 ;
  assign new_n15788 = lo0977 & ~lo0978 ;
  assign new_n15789 = ~lo0977 & lo0978 ;
  assign new_n15790 = ~new_n15788 & ~new_n15789 ;
  assign new_n15791 = lo0979 & ~lo0980 ;
  assign new_n15792 = ~lo0979 & lo0980 ;
  assign new_n15793 = ~new_n15791 & ~new_n15792 ;
  assign new_n15794 = lo1434 & new_n15793 ;
  assign new_n15795 = new_n15790 & new_n15794 ;
  assign new_n15796 = new_n14668 & new_n15795 ;
  assign new_n15797 = ~new_n15787 & ~new_n15796 ;
  assign new_n15798 = ~new_n15783 & new_n15797 ;
  assign new_n15799 = pi101 & new_n1985 ;
  assign new_n15800 = pi102 & new_n1987 ;
  assign new_n15801 = ~new_n15799 & ~new_n15800 ;
  assign new_n15802 = pi099 & new_n1979 ;
  assign new_n15803 = pi103 & new_n1989 ;
  assign new_n15804 = ~new_n15802 & ~new_n15803 ;
  assign new_n15805 = new_n15801 & new_n15804 ;
  assign new_n15806 = new_n15798 & new_n15805 ;
  assign new_n15807 = new_n15782 & new_n15806 ;
  assign new_n15808 = new_n15621 & ~new_n15807 ;
  assign new_n15809 = ~new_n15777 & ~new_n15808 ;
  assign new_n15810 = lo0138 & ~new_n15621 ;
  assign new_n15811 = pi108 & new_n1982 ;
  assign new_n15812 = pi105 & new_n1973 ;
  assign new_n15813 = pi106 & new_n1976 ;
  assign new_n15814 = ~new_n15812 & ~new_n15813 ;
  assign new_n15815 = ~new_n15811 & new_n15814 ;
  assign new_n15816 = pi112 & new_n1991 ;
  assign new_n15817 = lo0917 & lo0983 ;
  assign new_n15818 = ~lo0917 & lo0984 ;
  assign new_n15819 = ~new_n15817 & ~new_n15818 ;
  assign new_n15820 = new_n15154 & ~new_n15819 ;
  assign new_n15821 = lo0982 & new_n14668 ;
  assign new_n15822 = ~new_n15820 & ~new_n15821 ;
  assign new_n15823 = ~new_n15816 & new_n15822 ;
  assign new_n15824 = pi109 & new_n1985 ;
  assign new_n15825 = pi110 & new_n1987 ;
  assign new_n15826 = ~new_n15824 & ~new_n15825 ;
  assign new_n15827 = pi107 & new_n1979 ;
  assign new_n15828 = pi111 & new_n1989 ;
  assign new_n15829 = ~new_n15827 & ~new_n15828 ;
  assign new_n15830 = new_n15826 & new_n15829 ;
  assign new_n15831 = new_n15823 & new_n15830 ;
  assign new_n15832 = new_n15815 & new_n15831 ;
  assign new_n15833 = new_n15621 & ~new_n15832 ;
  assign new_n15834 = ~new_n15810 & ~new_n15833 ;
  assign new_n15835 = lo0139 & ~new_n15621 ;
  assign new_n15836 = lo0985 & new_n15621 ;
  assign new_n15837 = ~new_n15835 & ~new_n15836 ;
  assign new_n15838 = lo0140 & ~new_n15621 ;
  assign new_n15839 = pi116 & new_n1989 ;
  assign new_n15840 = pi114 & new_n1979 ;
  assign new_n15841 = pi115 & new_n1987 ;
  assign new_n15842 = ~new_n15840 & ~new_n15841 ;
  assign new_n15843 = ~new_n15839 & new_n15842 ;
  assign new_n15844 = lo0917 & lo0986 ;
  assign new_n15845 = ~lo0917 & ~lo1436 ;
  assign new_n15846 = ~new_n15844 & ~new_n15845 ;
  assign new_n15847 = new_n15154 & ~new_n15846 ;
  assign new_n15848 = pi120 & new_n1991 ;
  assign new_n15849 = ~new_n15847 & ~new_n15848 ;
  assign new_n15850 = pi118 & new_n1976 ;
  assign new_n15851 = pi119 & new_n1982 ;
  assign new_n15852 = ~new_n15850 & ~new_n15851 ;
  assign new_n15853 = pi113 & new_n1973 ;
  assign new_n15854 = pi117 & new_n1985 ;
  assign new_n15855 = ~new_n15853 & ~new_n15854 ;
  assign new_n15856 = new_n15852 & new_n15855 ;
  assign new_n15857 = new_n15849 & new_n15856 ;
  assign new_n15858 = new_n15843 & new_n15857 ;
  assign new_n15859 = new_n15621 & ~new_n15858 ;
  assign new_n15860 = ~new_n15838 & ~new_n15859 ;
  assign new_n15861 = lo0141 & ~new_n15621 ;
  assign new_n15862 = pi125 & new_n1982 ;
  assign new_n15863 = pi121 & new_n1987 ;
  assign new_n15864 = pi122 & new_n1989 ;
  assign new_n15865 = ~new_n15863 & ~new_n15864 ;
  assign new_n15866 = ~new_n15862 & new_n15865 ;
  assign new_n15867 = pi128 & new_n1991 ;
  assign new_n15868 = lo0987 & new_n14668 ;
  assign new_n15869 = lo0988 & new_n15207 ;
  assign new_n15870 = ~new_n15868 & ~new_n15869 ;
  assign new_n15871 = ~new_n15867 & new_n15870 ;
  assign new_n15872 = pi126 & new_n1985 ;
  assign new_n15873 = pi127 & new_n1973 ;
  assign new_n15874 = ~new_n15872 & ~new_n15873 ;
  assign new_n15875 = pi123 & new_n1976 ;
  assign new_n15876 = pi124 & new_n1979 ;
  assign new_n15877 = ~new_n15875 & ~new_n15876 ;
  assign new_n15878 = new_n15874 & new_n15877 ;
  assign new_n15879 = new_n15871 & new_n15878 ;
  assign new_n15880 = new_n15866 & new_n15879 ;
  assign new_n15881 = new_n15621 & ~new_n15880 ;
  assign new_n15882 = ~new_n15861 & ~new_n15881 ;
  assign new_n15883 = lo0142 & ~new_n15621 ;
  assign new_n15884 = lo0989 & new_n15621 ;
  assign new_n15885 = ~new_n15883 & ~new_n15884 ;
  assign new_n15886 = lo0143 & ~new_n15621 ;
  assign new_n15887 = pi132 & new_n1989 ;
  assign new_n15888 = pi130 & new_n1979 ;
  assign new_n15889 = pi131 & new_n1987 ;
  assign new_n15890 = ~new_n15888 & ~new_n15889 ;
  assign new_n15891 = ~new_n15887 & new_n15890 ;
  assign new_n15892 = lo0917 & lo0990 ;
  assign new_n15893 = ~lo0917 & ~lo1437 ;
  assign new_n15894 = ~new_n15892 & ~new_n15893 ;
  assign new_n15895 = new_n15154 & ~new_n15894 ;
  assign new_n15896 = pi136 & new_n1991 ;
  assign new_n15897 = ~new_n15895 & ~new_n15896 ;
  assign new_n15898 = pi134 & new_n1976 ;
  assign new_n15899 = pi135 & new_n1982 ;
  assign new_n15900 = ~new_n15898 & ~new_n15899 ;
  assign new_n15901 = pi129 & new_n1973 ;
  assign new_n15902 = pi133 & new_n1985 ;
  assign new_n15903 = ~new_n15901 & ~new_n15902 ;
  assign new_n15904 = new_n15900 & new_n15903 ;
  assign new_n15905 = new_n15897 & new_n15904 ;
  assign new_n15906 = new_n15891 & new_n15905 ;
  assign new_n15907 = new_n15621 & ~new_n15906 ;
  assign new_n15908 = ~new_n15886 & ~new_n15907 ;
  assign new_n15909 = lo0144 & ~new_n15621 ;
  assign new_n15910 = pi141 & new_n1982 ;
  assign new_n15911 = pi137 & new_n1987 ;
  assign new_n15912 = pi138 & new_n1989 ;
  assign new_n15913 = ~new_n15911 & ~new_n15912 ;
  assign new_n15914 = ~new_n15910 & new_n15913 ;
  assign new_n15915 = pi144 & new_n1991 ;
  assign new_n15916 = lo0991 & new_n14668 ;
  assign new_n15917 = lo0992 & new_n15207 ;
  assign new_n15918 = ~new_n15916 & ~new_n15917 ;
  assign new_n15919 = ~new_n15915 & new_n15918 ;
  assign new_n15920 = pi142 & new_n1985 ;
  assign new_n15921 = pi143 & new_n1973 ;
  assign new_n15922 = ~new_n15920 & ~new_n15921 ;
  assign new_n15923 = pi139 & new_n1976 ;
  assign new_n15924 = pi140 & new_n1979 ;
  assign new_n15925 = ~new_n15923 & ~new_n15924 ;
  assign new_n15926 = new_n15922 & new_n15925 ;
  assign new_n15927 = new_n15919 & new_n15926 ;
  assign new_n15928 = new_n15914 & new_n15927 ;
  assign new_n15929 = new_n15621 & ~new_n15928 ;
  assign new_n15930 = ~new_n15909 & ~new_n15929 ;
  assign new_n15931 = lo0145 & ~new_n15621 ;
  assign new_n15932 = lo0993 & new_n15621 ;
  assign new_n15933 = ~new_n15931 & ~new_n15932 ;
  assign new_n15934 = lo0146 & ~new_n15621 ;
  assign new_n15935 = pi145 & new_n1987 ;
  assign new_n15936 = pi146 & new_n1991 ;
  assign new_n15937 = pi152 & new_n1985 ;
  assign new_n15938 = ~new_n15936 & ~new_n15937 ;
  assign new_n15939 = ~new_n15935 & new_n15938 ;
  assign new_n15940 = pi151 & new_n1982 ;
  assign new_n15941 = lo0917 & lo0994 ;
  assign new_n15942 = ~lo0917 & ~lo1438 ;
  assign new_n15943 = ~new_n15941 & ~new_n15942 ;
  assign new_n15944 = new_n15154 & ~new_n15943 ;
  assign new_n15945 = pi004 & new_n2187 ;
  assign new_n15946 = ~lo0051 & lo0997 ;
  assign new_n15947 = ~lo0054 & new_n15946 ;
  assign new_n15948 = ~lo0051 & lo0996 ;
  assign new_n15949 = lo0054 & new_n15948 ;
  assign new_n15950 = ~new_n15236 & ~new_n15949 ;
  assign new_n15951 = ~new_n15947 & new_n15950 ;
  assign new_n15952 = ~lo0051 & ~new_n15951 ;
  assign new_n15953 = lo0051 & new_n15951 ;
  assign new_n15954 = ~new_n15952 & ~new_n15953 ;
  assign new_n15955 = lo0995 & ~new_n15954 ;
  assign new_n15956 = ~lo0995 & new_n15952 ;
  assign new_n15957 = lo0051 & lo0998 ;
  assign new_n15958 = ~new_n15951 & new_n15957 ;
  assign new_n15959 = ~new_n15956 & ~new_n15958 ;
  assign new_n15960 = ~new_n15955 & new_n15959 ;
  assign new_n15961 = new_n14668 & ~new_n15960 ;
  assign new_n15962 = ~new_n15945 & ~new_n15961 ;
  assign new_n15963 = ~new_n15944 & new_n15962 ;
  assign new_n15964 = ~new_n15940 & new_n15963 ;
  assign new_n15965 = pi148 & new_n1973 ;
  assign new_n15966 = pi149 & new_n1976 ;
  assign new_n15967 = ~new_n15965 & ~new_n15966 ;
  assign new_n15968 = pi147 & new_n1989 ;
  assign new_n15969 = pi150 & new_n1979 ;
  assign new_n15970 = ~new_n15968 & ~new_n15969 ;
  assign new_n15971 = new_n15967 & new_n15970 ;
  assign new_n15972 = new_n15964 & new_n15971 ;
  assign new_n15973 = new_n15939 & new_n15972 ;
  assign new_n15974 = new_n15621 & ~new_n15973 ;
  assign new_n15975 = ~new_n15934 & ~new_n15974 ;
  assign new_n15976 = lo0147 & ~new_n15621 ;
  assign new_n15977 = pi156 & new_n1982 ;
  assign new_n15978 = pi153 & new_n1973 ;
  assign new_n15979 = pi154 & new_n1976 ;
  assign new_n15980 = ~new_n15978 & ~new_n15979 ;
  assign new_n15981 = ~new_n15977 & new_n15980 ;
  assign new_n15982 = pi160 & new_n1991 ;
  assign new_n15983 = lo0917 & lo1000 ;
  assign new_n15984 = lo0186 & ~lo0917 ;
  assign new_n15985 = ~new_n15983 & ~new_n15984 ;
  assign new_n15986 = new_n15154 & ~new_n15985 ;
  assign new_n15987 = lo0999 & new_n14668 ;
  assign new_n15988 = ~new_n15986 & ~new_n15987 ;
  assign new_n15989 = ~new_n15982 & new_n15988 ;
  assign new_n15990 = pi157 & new_n1985 ;
  assign new_n15991 = pi158 & new_n1987 ;
  assign new_n15992 = ~new_n15990 & ~new_n15991 ;
  assign new_n15993 = pi155 & new_n1979 ;
  assign new_n15994 = pi159 & new_n1989 ;
  assign new_n15995 = ~new_n15993 & ~new_n15994 ;
  assign new_n15996 = new_n15992 & new_n15995 ;
  assign new_n15997 = new_n15989 & new_n15996 ;
  assign new_n15998 = new_n15981 & new_n15997 ;
  assign new_n15999 = new_n15621 & ~new_n15998 ;
  assign new_n16000 = ~new_n15976 & ~new_n15999 ;
  assign new_n16001 = lo0148 & ~new_n15621 ;
  assign new_n16002 = lo1001 & new_n15621 ;
  assign new_n16003 = ~new_n16001 & ~new_n16002 ;
  assign new_n16004 = lo0149 & ~new_n15621 ;
  assign new_n16005 = ~new_n15288 & new_n15621 ;
  assign new_n16006 = ~new_n16004 & ~new_n16005 ;
  assign new_n16007 = lo0150 & ~new_n15621 ;
  assign new_n16008 = ~new_n15313 & new_n15621 ;
  assign new_n16009 = ~new_n16007 & ~new_n16008 ;
  assign new_n16010 = lo0151 & ~new_n15621 ;
  assign new_n16011 = lo1002 & new_n15621 ;
  assign new_n16012 = ~new_n16010 & ~new_n16011 ;
  assign new_n16013 = lo0152 & ~new_n15621 ;
  assign new_n16014 = pi161 & new_n1987 ;
  assign new_n16015 = pi162 & new_n1991 ;
  assign new_n16016 = pi168 & new_n1985 ;
  assign new_n16017 = ~new_n16015 & ~new_n16016 ;
  assign new_n16018 = ~new_n16014 & new_n16017 ;
  assign new_n16019 = pi167 & new_n1982 ;
  assign new_n16020 = lo0917 & lo1003 ;
  assign new_n16021 = ~lo0917 & ~lo1439 ;
  assign new_n16022 = ~new_n16020 & ~new_n16021 ;
  assign new_n16023 = new_n15154 & ~new_n16022 ;
  assign new_n16024 = pi005 & new_n2187 ;
  assign new_n16025 = ~lo0054 & lo1006 ;
  assign new_n16026 = ~lo0051 & new_n16025 ;
  assign new_n16027 = ~lo0054 & lo1005 ;
  assign new_n16028 = lo0051 & new_n16027 ;
  assign new_n16029 = ~new_n15236 & ~new_n16028 ;
  assign new_n16030 = ~new_n16026 & new_n16029 ;
  assign new_n16031 = ~lo0054 & ~new_n16030 ;
  assign new_n16032 = lo0054 & new_n16030 ;
  assign new_n16033 = ~new_n16031 & ~new_n16032 ;
  assign new_n16034 = lo1004 & ~new_n16033 ;
  assign new_n16035 = ~lo1004 & new_n16031 ;
  assign new_n16036 = lo0054 & lo1007 ;
  assign new_n16037 = ~new_n16030 & new_n16036 ;
  assign new_n16038 = ~new_n16035 & ~new_n16037 ;
  assign new_n16039 = ~new_n16034 & new_n16038 ;
  assign new_n16040 = new_n14668 & ~new_n16039 ;
  assign new_n16041 = ~new_n16024 & ~new_n16040 ;
  assign new_n16042 = ~new_n16023 & new_n16041 ;
  assign new_n16043 = ~new_n16019 & new_n16042 ;
  assign new_n16044 = pi164 & new_n1973 ;
  assign new_n16045 = pi165 & new_n1976 ;
  assign new_n16046 = ~new_n16044 & ~new_n16045 ;
  assign new_n16047 = pi163 & new_n1989 ;
  assign new_n16048 = pi166 & new_n1979 ;
  assign new_n16049 = ~new_n16047 & ~new_n16048 ;
  assign new_n16050 = new_n16046 & new_n16049 ;
  assign new_n16051 = new_n16043 & new_n16050 ;
  assign new_n16052 = new_n16018 & new_n16051 ;
  assign new_n16053 = new_n15621 & ~new_n16052 ;
  assign new_n16054 = ~new_n16013 & ~new_n16053 ;
  assign new_n16055 = lo0153 & ~new_n15621 ;
  assign new_n16056 = pi169 & new_n1987 ;
  assign new_n16057 = pi170 & new_n1991 ;
  assign new_n16058 = pi176 & new_n1985 ;
  assign new_n16059 = ~new_n16057 & ~new_n16058 ;
  assign new_n16060 = ~new_n16056 & new_n16059 ;
  assign new_n16061 = pi175 & new_n1982 ;
  assign new_n16062 = lo0917 & lo1008 ;
  assign new_n16063 = lo0880 & ~lo0917 ;
  assign new_n16064 = ~new_n16062 & ~new_n16063 ;
  assign new_n16065 = new_n15154 & ~new_n16064 ;
  assign new_n16066 = pi006 & new_n2187 ;
  assign new_n16067 = lo1009 & new_n14668 ;
  assign new_n16068 = ~new_n16066 & ~new_n16067 ;
  assign new_n16069 = ~new_n16065 & new_n16068 ;
  assign new_n16070 = ~new_n16061 & new_n16069 ;
  assign new_n16071 = pi172 & new_n1973 ;
  assign new_n16072 = pi173 & new_n1976 ;
  assign new_n16073 = ~new_n16071 & ~new_n16072 ;
  assign new_n16074 = pi171 & new_n1989 ;
  assign new_n16075 = pi174 & new_n1979 ;
  assign new_n16076 = ~new_n16074 & ~new_n16075 ;
  assign new_n16077 = new_n16073 & new_n16076 ;
  assign new_n16078 = new_n16070 & new_n16077 ;
  assign new_n16079 = new_n16060 & new_n16078 ;
  assign new_n16080 = new_n15621 & ~new_n16079 ;
  assign new_n16081 = ~new_n16055 & ~new_n16080 ;
  assign new_n16082 = lo0154 & ~new_n15621 ;
  assign new_n16083 = lo1010 & new_n15621 ;
  assign new_n16084 = ~new_n16082 & ~new_n16083 ;
  assign new_n16085 = lo0155 & ~new_n15621 ;
  assign new_n16086 = pi180 & new_n1989 ;
  assign new_n16087 = pi178 & new_n1979 ;
  assign new_n16088 = pi179 & new_n1987 ;
  assign new_n16089 = ~new_n16087 & ~new_n16088 ;
  assign new_n16090 = ~new_n16086 & new_n16089 ;
  assign new_n16091 = lo0917 & lo1011 ;
  assign new_n16092 = lo0864 & ~lo0917 ;
  assign new_n16093 = ~new_n16091 & ~new_n16092 ;
  assign new_n16094 = new_n15154 & ~new_n16093 ;
  assign new_n16095 = pi184 & new_n1991 ;
  assign new_n16096 = ~new_n16094 & ~new_n16095 ;
  assign new_n16097 = pi182 & new_n1976 ;
  assign new_n16098 = pi183 & new_n1982 ;
  assign new_n16099 = ~new_n16097 & ~new_n16098 ;
  assign new_n16100 = pi177 & new_n1973 ;
  assign new_n16101 = pi181 & new_n1985 ;
  assign new_n16102 = ~new_n16100 & ~new_n16101 ;
  assign new_n16103 = new_n16099 & new_n16102 ;
  assign new_n16104 = new_n16096 & new_n16103 ;
  assign new_n16105 = new_n16090 & new_n16104 ;
  assign new_n16106 = new_n15621 & ~new_n16105 ;
  assign new_n16107 = ~new_n16085 & ~new_n16106 ;
  assign new_n16108 = lo0156 & ~new_n15621 ;
  assign new_n16109 = pi189 & new_n1982 ;
  assign new_n16110 = pi185 & new_n1987 ;
  assign new_n16111 = pi186 & new_n1989 ;
  assign new_n16112 = ~new_n16110 & ~new_n16111 ;
  assign new_n16113 = ~new_n16109 & new_n16112 ;
  assign new_n16114 = pi192 & new_n1991 ;
  assign new_n16115 = lo1012 & new_n14668 ;
  assign new_n16116 = lo1013 & new_n15207 ;
  assign new_n16117 = ~new_n16115 & ~new_n16116 ;
  assign new_n16118 = ~new_n16114 & new_n16117 ;
  assign new_n16119 = pi190 & new_n1985 ;
  assign new_n16120 = pi191 & new_n1973 ;
  assign new_n16121 = ~new_n16119 & ~new_n16120 ;
  assign new_n16122 = pi187 & new_n1976 ;
  assign new_n16123 = pi188 & new_n1979 ;
  assign new_n16124 = ~new_n16122 & ~new_n16123 ;
  assign new_n16125 = new_n16121 & new_n16124 ;
  assign new_n16126 = new_n16118 & new_n16125 ;
  assign new_n16127 = new_n16113 & new_n16126 ;
  assign new_n16128 = new_n15621 & ~new_n16127 ;
  assign new_n16129 = ~new_n16108 & ~new_n16128 ;
  assign new_n16130 = lo0157 & ~new_n15621 ;
  assign new_n16131 = lo1014 & new_n15621 ;
  assign new_n16132 = ~new_n16130 & ~new_n16131 ;
  assign new_n16133 = lo0158 & ~new_n15621 ;
  assign new_n16134 = pi196 & new_n1989 ;
  assign new_n16135 = pi194 & new_n1979 ;
  assign new_n16136 = pi195 & new_n1987 ;
  assign new_n16137 = ~new_n16135 & ~new_n16136 ;
  assign new_n16138 = ~new_n16134 & new_n16137 ;
  assign new_n16139 = lo0917 & lo1015 ;
  assign new_n16140 = lo0862 & ~lo0917 ;
  assign new_n16141 = ~new_n16139 & ~new_n16140 ;
  assign new_n16142 = new_n15154 & ~new_n16141 ;
  assign new_n16143 = pi200 & new_n1991 ;
  assign new_n16144 = ~new_n16142 & ~new_n16143 ;
  assign new_n16145 = pi198 & new_n1976 ;
  assign new_n16146 = pi199 & new_n1982 ;
  assign new_n16147 = ~new_n16145 & ~new_n16146 ;
  assign new_n16148 = pi193 & new_n1973 ;
  assign new_n16149 = pi197 & new_n1985 ;
  assign new_n16150 = ~new_n16148 & ~new_n16149 ;
  assign new_n16151 = new_n16147 & new_n16150 ;
  assign new_n16152 = new_n16144 & new_n16151 ;
  assign new_n16153 = new_n16138 & new_n16152 ;
  assign new_n16154 = new_n15621 & ~new_n16153 ;
  assign new_n16155 = ~new_n16133 & ~new_n16154 ;
  assign new_n16156 = lo0159 & ~new_n15621 ;
  assign new_n16157 = pi205 & new_n1982 ;
  assign new_n16158 = pi201 & new_n1987 ;
  assign new_n16159 = pi202 & new_n1989 ;
  assign new_n16160 = ~new_n16158 & ~new_n16159 ;
  assign new_n16161 = ~new_n16157 & new_n16160 ;
  assign new_n16162 = pi208 & new_n1991 ;
  assign new_n16163 = lo1016 & new_n14668 ;
  assign new_n16164 = lo1017 & new_n15207 ;
  assign new_n16165 = ~new_n16163 & ~new_n16164 ;
  assign new_n16166 = ~new_n16162 & new_n16165 ;
  assign new_n16167 = pi206 & new_n1985 ;
  assign new_n16168 = pi207 & new_n1973 ;
  assign new_n16169 = ~new_n16167 & ~new_n16168 ;
  assign new_n16170 = pi203 & new_n1976 ;
  assign new_n16171 = pi204 & new_n1979 ;
  assign new_n16172 = ~new_n16170 & ~new_n16171 ;
  assign new_n16173 = new_n16169 & new_n16172 ;
  assign new_n16174 = new_n16166 & new_n16173 ;
  assign new_n16175 = new_n16161 & new_n16174 ;
  assign new_n16176 = new_n15621 & ~new_n16175 ;
  assign new_n16177 = ~new_n16156 & ~new_n16176 ;
  assign new_n16178 = lo0160 & ~new_n15621 ;
  assign new_n16179 = lo1018 & new_n15621 ;
  assign new_n16180 = ~new_n16178 & ~new_n16179 ;
  assign new_n16181 = lo0161 & ~new_n15621 ;
  assign new_n16182 = ~new_n15262 & new_n15621 ;
  assign new_n16183 = ~new_n16181 & ~new_n16182 ;
  assign new_n16184 = lo0162 & ~new_n15621 ;
  assign new_n16185 = ~new_n15170 & new_n15621 ;
  assign new_n16186 = ~new_n16184 & ~new_n16185 ;
  assign new_n16187 = lo0163 & ~new_n15621 ;
  assign new_n16188 = lo1019 & new_n15621 ;
  assign new_n16189 = ~new_n16187 & ~new_n16188 ;
  assign new_n16190 = lo0164 & ~new_n15621 ;
  assign new_n16191 = pi209 & new_n1987 ;
  assign new_n16192 = pi210 & new_n1991 ;
  assign new_n16193 = pi216 & new_n1985 ;
  assign new_n16194 = ~new_n16192 & ~new_n16193 ;
  assign new_n16195 = ~new_n16191 & new_n16194 ;
  assign new_n16196 = pi215 & new_n1982 ;
  assign new_n16197 = lo0917 & lo1020 ;
  assign new_n16198 = ~lo0917 & ~lo1440 ;
  assign new_n16199 = ~new_n16197 & ~new_n16198 ;
  assign new_n16200 = new_n15154 & ~new_n16199 ;
  assign new_n16201 = pi007 & new_n2187 ;
  assign new_n16202 = ~lo0051 & lo1023 ;
  assign new_n16203 = ~lo0054 & new_n16202 ;
  assign new_n16204 = ~lo0051 & lo1022 ;
  assign new_n16205 = lo0054 & new_n16204 ;
  assign new_n16206 = ~new_n15236 & ~new_n16205 ;
  assign new_n16207 = ~new_n16203 & new_n16206 ;
  assign new_n16208 = ~lo0051 & ~new_n16207 ;
  assign new_n16209 = lo0051 & new_n16207 ;
  assign new_n16210 = ~new_n16208 & ~new_n16209 ;
  assign new_n16211 = lo1021 & ~new_n16210 ;
  assign new_n16212 = ~lo1021 & new_n16208 ;
  assign new_n16213 = lo0051 & lo1024 ;
  assign new_n16214 = ~new_n16207 & new_n16213 ;
  assign new_n16215 = ~new_n16212 & ~new_n16214 ;
  assign new_n16216 = ~new_n16211 & new_n16215 ;
  assign new_n16217 = new_n14668 & ~new_n16216 ;
  assign new_n16218 = ~new_n16201 & ~new_n16217 ;
  assign new_n16219 = ~new_n16200 & new_n16218 ;
  assign new_n16220 = ~new_n16196 & new_n16219 ;
  assign new_n16221 = pi212 & new_n1973 ;
  assign new_n16222 = pi213 & new_n1976 ;
  assign new_n16223 = ~new_n16221 & ~new_n16222 ;
  assign new_n16224 = pi211 & new_n1989 ;
  assign new_n16225 = pi214 & new_n1979 ;
  assign new_n16226 = ~new_n16224 & ~new_n16225 ;
  assign new_n16227 = new_n16223 & new_n16226 ;
  assign new_n16228 = new_n16220 & new_n16227 ;
  assign new_n16229 = new_n16195 & new_n16228 ;
  assign new_n16230 = new_n15621 & ~new_n16229 ;
  assign new_n16231 = ~new_n16190 & ~new_n16230 ;
  assign new_n16232 = lo0165 & ~new_n15621 ;
  assign new_n16233 = pi220 & new_n1982 ;
  assign new_n16234 = pi217 & new_n1973 ;
  assign new_n16235 = pi218 & new_n1976 ;
  assign new_n16236 = ~new_n16234 & ~new_n16235 ;
  assign new_n16237 = ~new_n16233 & new_n16236 ;
  assign new_n16238 = pi224 & new_n1991 ;
  assign new_n16239 = lo0917 & lo1026 ;
  assign new_n16240 = lo0184 & ~lo0917 ;
  assign new_n16241 = ~new_n16239 & ~new_n16240 ;
  assign new_n16242 = new_n15154 & ~new_n16241 ;
  assign new_n16243 = lo1025 & new_n14668 ;
  assign new_n16244 = ~new_n16242 & ~new_n16243 ;
  assign new_n16245 = ~new_n16238 & new_n16244 ;
  assign new_n16246 = pi221 & new_n1985 ;
  assign new_n16247 = pi222 & new_n1987 ;
  assign new_n16248 = ~new_n16246 & ~new_n16247 ;
  assign new_n16249 = pi219 & new_n1979 ;
  assign new_n16250 = pi223 & new_n1989 ;
  assign new_n16251 = ~new_n16249 & ~new_n16250 ;
  assign new_n16252 = new_n16248 & new_n16251 ;
  assign new_n16253 = new_n16245 & new_n16252 ;
  assign new_n16254 = new_n16237 & new_n16253 ;
  assign new_n16255 = new_n15621 & ~new_n16254 ;
  assign new_n16256 = ~new_n16232 & ~new_n16255 ;
  assign new_n16257 = lo0166 & ~new_n15621 ;
  assign new_n16258 = lo1027 & new_n15621 ;
  assign new_n16259 = ~new_n16257 & ~new_n16258 ;
  assign new_n16260 = lo0167 & ~new_n15621 ;
  assign new_n16261 = pi225 & new_n1987 ;
  assign new_n16262 = pi226 & new_n1991 ;
  assign new_n16263 = pi232 & new_n1985 ;
  assign new_n16264 = ~new_n16262 & ~new_n16263 ;
  assign new_n16265 = ~new_n16261 & new_n16264 ;
  assign new_n16266 = pi231 & new_n1982 ;
  assign new_n16267 = lo0917 & lo1028 ;
  assign new_n16268 = ~lo0917 & ~lo1441 ;
  assign new_n16269 = ~new_n16267 & ~new_n16268 ;
  assign new_n16270 = new_n15154 & ~new_n16269 ;
  assign new_n16271 = pi008 & new_n2187 ;
  assign new_n16272 = ~lo0051 & lo1031 ;
  assign new_n16273 = ~lo0054 & new_n16272 ;
  assign new_n16274 = ~lo0051 & lo1030 ;
  assign new_n16275 = lo0054 & new_n16274 ;
  assign new_n16276 = ~new_n15236 & ~new_n16275 ;
  assign new_n16277 = ~new_n16273 & new_n16276 ;
  assign new_n16278 = ~lo0051 & ~new_n16277 ;
  assign new_n16279 = lo0051 & new_n16277 ;
  assign new_n16280 = ~new_n16278 & ~new_n16279 ;
  assign new_n16281 = lo1029 & ~new_n16280 ;
  assign new_n16282 = ~lo1029 & new_n16278 ;
  assign new_n16283 = lo0051 & lo1032 ;
  assign new_n16284 = ~new_n16277 & new_n16283 ;
  assign new_n16285 = ~new_n16282 & ~new_n16284 ;
  assign new_n16286 = ~new_n16281 & new_n16285 ;
  assign new_n16287 = new_n14668 & ~new_n16286 ;
  assign new_n16288 = ~new_n16271 & ~new_n16287 ;
  assign new_n16289 = ~new_n16270 & new_n16288 ;
  assign new_n16290 = ~new_n16266 & new_n16289 ;
  assign new_n16291 = pi228 & new_n1973 ;
  assign new_n16292 = pi229 & new_n1976 ;
  assign new_n16293 = ~new_n16291 & ~new_n16292 ;
  assign new_n16294 = pi227 & new_n1989 ;
  assign new_n16295 = pi230 & new_n1979 ;
  assign new_n16296 = ~new_n16294 & ~new_n16295 ;
  assign new_n16297 = new_n16293 & new_n16296 ;
  assign new_n16298 = new_n16290 & new_n16297 ;
  assign new_n16299 = new_n16265 & new_n16298 ;
  assign new_n16300 = new_n15621 & ~new_n16299 ;
  assign new_n16301 = ~new_n16260 & ~new_n16300 ;
  assign new_n16302 = lo0168 & ~new_n15621 ;
  assign new_n16303 = pi233 & new_n1987 ;
  assign new_n16304 = pi234 & new_n1991 ;
  assign new_n16305 = pi240 & new_n1985 ;
  assign new_n16306 = ~new_n16304 & ~new_n16305 ;
  assign new_n16307 = ~new_n16303 & new_n16306 ;
  assign new_n16308 = pi239 & new_n1982 ;
  assign new_n16309 = lo0917 & lo1033 ;
  assign new_n16310 = lo0871 & ~lo0917 ;
  assign new_n16311 = ~new_n16309 & ~new_n16310 ;
  assign new_n16312 = new_n15154 & ~new_n16311 ;
  assign new_n16313 = pi009 & new_n2187 ;
  assign new_n16314 = lo1034 & new_n14668 ;
  assign new_n16315 = ~new_n16313 & ~new_n16314 ;
  assign new_n16316 = ~new_n16312 & new_n16315 ;
  assign new_n16317 = ~new_n16308 & new_n16316 ;
  assign new_n16318 = pi236 & new_n1973 ;
  assign new_n16319 = pi237 & new_n1976 ;
  assign new_n16320 = ~new_n16318 & ~new_n16319 ;
  assign new_n16321 = pi235 & new_n1989 ;
  assign new_n16322 = pi238 & new_n1979 ;
  assign new_n16323 = ~new_n16321 & ~new_n16322 ;
  assign new_n16324 = new_n16320 & new_n16323 ;
  assign new_n16325 = new_n16317 & new_n16324 ;
  assign new_n16326 = new_n16307 & new_n16325 ;
  assign new_n16327 = new_n15621 & ~new_n16326 ;
  assign new_n16328 = ~new_n16302 & ~new_n16327 ;
  assign new_n16329 = lo0169 & ~new_n15621 ;
  assign new_n16330 = lo1035 & new_n15621 ;
  assign new_n16331 = ~new_n16329 & ~new_n16330 ;
  assign new_n16332 = lo0170 & ~new_n15621 ;
  assign new_n16333 = pi241 & new_n1987 ;
  assign new_n16334 = pi242 & new_n1991 ;
  assign new_n16335 = pi248 & new_n1985 ;
  assign new_n16336 = ~new_n16334 & ~new_n16335 ;
  assign new_n16337 = ~new_n16333 & new_n16336 ;
  assign new_n16338 = pi247 & new_n1982 ;
  assign new_n16339 = lo0917 & lo1036 ;
  assign new_n16340 = ~lo0917 & ~lo1442 ;
  assign new_n16341 = ~new_n16339 & ~new_n16340 ;
  assign new_n16342 = new_n15154 & ~new_n16341 ;
  assign new_n16343 = pi010 & new_n2187 ;
  assign new_n16344 = ~lo0051 & lo1039 ;
  assign new_n16345 = ~lo0054 & new_n16344 ;
  assign new_n16346 = ~lo0051 & lo1038 ;
  assign new_n16347 = lo0054 & new_n16346 ;
  assign new_n16348 = ~new_n15236 & ~new_n16347 ;
  assign new_n16349 = ~new_n16345 & new_n16348 ;
  assign new_n16350 = ~lo0051 & ~new_n16349 ;
  assign new_n16351 = lo0051 & new_n16349 ;
  assign new_n16352 = ~new_n16350 & ~new_n16351 ;
  assign new_n16353 = lo1037 & ~new_n16352 ;
  assign new_n16354 = ~lo1037 & new_n16350 ;
  assign new_n16355 = lo0051 & lo1040 ;
  assign new_n16356 = ~new_n16349 & new_n16355 ;
  assign new_n16357 = ~new_n16354 & ~new_n16356 ;
  assign new_n16358 = ~new_n16353 & new_n16357 ;
  assign new_n16359 = new_n14668 & ~new_n16358 ;
  assign new_n16360 = ~new_n16343 & ~new_n16359 ;
  assign new_n16361 = ~new_n16342 & new_n16360 ;
  assign new_n16362 = ~new_n16338 & new_n16361 ;
  assign new_n16363 = pi244 & new_n1973 ;
  assign new_n16364 = pi245 & new_n1976 ;
  assign new_n16365 = ~new_n16363 & ~new_n16364 ;
  assign new_n16366 = pi243 & new_n1989 ;
  assign new_n16367 = pi246 & new_n1979 ;
  assign new_n16368 = ~new_n16366 & ~new_n16367 ;
  assign new_n16369 = new_n16365 & new_n16368 ;
  assign new_n16370 = new_n16362 & new_n16369 ;
  assign new_n16371 = new_n16337 & new_n16370 ;
  assign new_n16372 = new_n15621 & ~new_n16371 ;
  assign new_n16373 = ~new_n16332 & ~new_n16372 ;
  assign new_n16374 = lo0171 & ~new_n15621 ;
  assign new_n16375 = pi249 & new_n1987 ;
  assign new_n16376 = pi250 & new_n1991 ;
  assign new_n16377 = pi256 & new_n1985 ;
  assign new_n16378 = ~new_n16376 & ~new_n16377 ;
  assign new_n16379 = ~new_n16375 & new_n16378 ;
  assign new_n16380 = pi255 & new_n1982 ;
  assign new_n16381 = lo0917 & lo1041 ;
  assign new_n16382 = lo0188 & ~lo0917 ;
  assign new_n16383 = ~new_n16381 & ~new_n16382 ;
  assign new_n16384 = new_n15154 & ~new_n16383 ;
  assign new_n16385 = pi011 & new_n2187 ;
  assign new_n16386 = lo1042 & new_n14668 ;
  assign new_n16387 = ~new_n16385 & ~new_n16386 ;
  assign new_n16388 = ~new_n16384 & new_n16387 ;
  assign new_n16389 = ~new_n16380 & new_n16388 ;
  assign new_n16390 = pi252 & new_n1973 ;
  assign new_n16391 = pi253 & new_n1976 ;
  assign new_n16392 = ~new_n16390 & ~new_n16391 ;
  assign new_n16393 = pi251 & new_n1989 ;
  assign new_n16394 = pi254 & new_n1979 ;
  assign new_n16395 = ~new_n16393 & ~new_n16394 ;
  assign new_n16396 = new_n16392 & new_n16395 ;
  assign new_n16397 = new_n16389 & new_n16396 ;
  assign new_n16398 = new_n16379 & new_n16397 ;
  assign new_n16399 = new_n15621 & ~new_n16398 ;
  assign new_n16400 = ~new_n16374 & ~new_n16399 ;
  assign new_n16401 = lo0172 & ~new_n15621 ;
  assign new_n16402 = lo1043 & new_n15621 ;
  assign new_n16403 = ~new_n16401 & ~new_n16402 ;
  assign new_n16404 = lo0173 & ~new_n15621 ;
  assign new_n16405 = pi257 & new_n1987 ;
  assign new_n16406 = pi258 & new_n1991 ;
  assign new_n16407 = pi264 & new_n1985 ;
  assign new_n16408 = ~new_n16406 & ~new_n16407 ;
  assign new_n16409 = ~new_n16405 & new_n16408 ;
  assign new_n16410 = pi263 & new_n1982 ;
  assign new_n16411 = lo0917 & lo1044 ;
  assign new_n16412 = ~lo0917 & ~lo1443 ;
  assign new_n16413 = ~new_n16411 & ~new_n16412 ;
  assign new_n16414 = new_n15154 & ~new_n16413 ;
  assign new_n16415 = pi012 & new_n2187 ;
  assign new_n16416 = ~lo0054 & lo1047 ;
  assign new_n16417 = ~lo0051 & new_n16416 ;
  assign new_n16418 = ~lo0054 & lo1046 ;
  assign new_n16419 = lo0051 & new_n16418 ;
  assign new_n16420 = ~new_n15236 & ~new_n16419 ;
  assign new_n16421 = ~new_n16417 & new_n16420 ;
  assign new_n16422 = ~lo0054 & ~new_n16421 ;
  assign new_n16423 = lo0054 & new_n16421 ;
  assign new_n16424 = ~new_n16422 & ~new_n16423 ;
  assign new_n16425 = lo1045 & ~new_n16424 ;
  assign new_n16426 = ~lo1045 & new_n16422 ;
  assign new_n16427 = lo0054 & lo1048 ;
  assign new_n16428 = ~new_n16421 & new_n16427 ;
  assign new_n16429 = ~new_n16426 & ~new_n16428 ;
  assign new_n16430 = ~new_n16425 & new_n16429 ;
  assign new_n16431 = new_n14668 & ~new_n16430 ;
  assign new_n16432 = ~new_n16415 & ~new_n16431 ;
  assign new_n16433 = ~new_n16414 & new_n16432 ;
  assign new_n16434 = ~new_n16410 & new_n16433 ;
  assign new_n16435 = pi260 & new_n1973 ;
  assign new_n16436 = pi261 & new_n1976 ;
  assign new_n16437 = ~new_n16435 & ~new_n16436 ;
  assign new_n16438 = pi259 & new_n1989 ;
  assign new_n16439 = pi262 & new_n1979 ;
  assign new_n16440 = ~new_n16438 & ~new_n16439 ;
  assign new_n16441 = new_n16437 & new_n16440 ;
  assign new_n16442 = new_n16434 & new_n16441 ;
  assign new_n16443 = new_n16409 & new_n16442 ;
  assign new_n16444 = new_n15621 & ~new_n16443 ;
  assign new_n16445 = ~new_n16404 & ~new_n16444 ;
  assign new_n16446 = lo0174 & ~new_n15621 ;
  assign new_n16447 = pi265 & new_n1987 ;
  assign new_n16448 = pi266 & new_n1991 ;
  assign new_n16449 = pi272 & new_n1985 ;
  assign new_n16450 = ~new_n16448 & ~new_n16449 ;
  assign new_n16451 = ~new_n16447 & new_n16450 ;
  assign new_n16452 = pi271 & new_n1982 ;
  assign new_n16453 = lo0917 & lo1049 ;
  assign new_n16454 = lo0869 & ~lo0917 ;
  assign new_n16455 = ~new_n16453 & ~new_n16454 ;
  assign new_n16456 = new_n15154 & ~new_n16455 ;
  assign new_n16457 = pi013 & new_n2187 ;
  assign new_n16458 = lo1050 & new_n14668 ;
  assign new_n16459 = ~new_n16457 & ~new_n16458 ;
  assign new_n16460 = ~new_n16456 & new_n16459 ;
  assign new_n16461 = ~new_n16452 & new_n16460 ;
  assign new_n16462 = pi268 & new_n1973 ;
  assign new_n16463 = pi269 & new_n1976 ;
  assign new_n16464 = ~new_n16462 & ~new_n16463 ;
  assign new_n16465 = pi267 & new_n1989 ;
  assign new_n16466 = pi270 & new_n1979 ;
  assign new_n16467 = ~new_n16465 & ~new_n16466 ;
  assign new_n16468 = new_n16464 & new_n16467 ;
  assign new_n16469 = new_n16461 & new_n16468 ;
  assign new_n16470 = new_n16451 & new_n16469 ;
  assign new_n16471 = new_n15621 & ~new_n16470 ;
  assign new_n16472 = ~new_n16446 & ~new_n16471 ;
  assign new_n16473 = new_n2264 & new_n12325 ;
  assign new_n16474 = ~new_n15374 & ~new_n16473 ;
  assign new_n16475 = ~new_n2252 & new_n15373 ;
  assign new_n16476 = ~new_n16474 & new_n16475 ;
  assign new_n16477 = new_n2436 & new_n16476 ;
  assign new_n16478 = lo0175 & ~new_n16477 ;
  assign new_n16479 = ~lo0917 & ~new_n2249 ;
  assign new_n16480 = new_n15154 & new_n16479 ;
  assign new_n16481 = new_n2002 & new_n16480 ;
  assign new_n16482 = lo1052 & new_n16481 ;
  assign new_n16483 = lo0018 & ~new_n2249 ;
  assign new_n16484 = lo0043 & lo0045 ;
  assign new_n16485 = lo0892 & ~lo1051 ;
  assign new_n16486 = ~lo0046 & new_n16485 ;
  assign new_n16487 = new_n16484 & new_n16486 ;
  assign new_n16488 = ~lo0043 & lo0892 ;
  assign new_n16489 = ~lo0045 & new_n16488 ;
  assign new_n16490 = ~lo0892 & ~lo0893 ;
  assign new_n16491 = new_n16484 & ~new_n16490 ;
  assign new_n16492 = ~new_n16489 & ~new_n16491 ;
  assign new_n16493 = lo0046 & lo1051 ;
  assign new_n16494 = ~new_n16492 & new_n16493 ;
  assign new_n16495 = ~new_n16487 & ~new_n16494 ;
  assign new_n16496 = new_n16483 & ~new_n16495 ;
  assign new_n16497 = ~new_n16482 & ~new_n16496 ;
  assign new_n16498 = ~new_n16478 & new_n16497 ;
  assign new_n16499 = lo1053 & new_n1993 ;
  assign new_n16500 = new_n16480 & new_n16499 ;
  assign new_n16501 = lo0176 & ~new_n16476 ;
  assign new_n16502 = ~new_n16500 & ~new_n16501 ;
  assign new_n16503 = lo1054 & new_n16481 ;
  assign new_n16504 = new_n2413 & new_n16476 ;
  assign new_n16505 = lo0177 & ~new_n16504 ;
  assign new_n16506 = ~new_n16503 & ~new_n16505 ;
  assign new_n16507 = lo0178 & new_n2252 ;
  assign new_n16508 = new_n12495 & new_n13863 ;
  assign new_n16509 = ~new_n12737 & ~new_n16508 ;
  assign new_n16510 = ~new_n2252 & ~new_n12452 ;
  assign new_n16511 = new_n13809 & new_n16510 ;
  assign new_n16512 = ~new_n16509 & new_n16511 ;
  assign new_n16513 = ~new_n16507 & ~new_n16512 ;
  assign new_n16514 = new_n2437 & new_n16476 ;
  assign new_n16515 = lo0179 & ~new_n16514 ;
  assign new_n16516 = lo1055 & new_n16481 ;
  assign new_n16517 = lo1433 & lo1435 ;
  assign new_n16518 = lo1432 & lo1438 ;
  assign new_n16519 = new_n16517 & new_n16518 ;
  assign new_n16520 = lo1431 & lo1439 ;
  assign new_n16521 = lo1436 & lo1437 ;
  assign new_n16522 = new_n16520 & new_n16521 ;
  assign new_n16523 = lo1442 & lo1443 ;
  assign new_n16524 = lo1440 & lo1441 ;
  assign new_n16525 = new_n16523 & new_n16524 ;
  assign new_n16526 = new_n16522 & new_n16525 ;
  assign new_n16527 = new_n16519 & new_n16526 ;
  assign new_n16528 = ~new_n16516 & ~new_n16527 ;
  assign new_n16529 = ~new_n16515 & new_n16528 ;
  assign new_n16530 = new_n2435 & new_n16504 ;
  assign new_n16531 = lo0180 & ~new_n16530 ;
  assign new_n16532 = lo1061 & new_n16481 ;
  assign new_n16533 = ~lo0031 & lo0918 ;
  assign new_n16534 = lo0930 & ~new_n16533 ;
  assign new_n16535 = ~lo0965 & lo1060 ;
  assign new_n16536 = lo0031 & ~lo0918 ;
  assign new_n16537 = ~new_n16535 & ~new_n16536 ;
  assign new_n16538 = ~lo0029 & lo0983 ;
  assign new_n16539 = lo0965 & ~lo1060 ;
  assign new_n16540 = ~new_n16538 & ~new_n16539 ;
  assign new_n16541 = new_n16537 & new_n16540 ;
  assign new_n16542 = new_n16534 & new_n16541 ;
  assign new_n16543 = ~lo0032 & lo1026 ;
  assign new_n16544 = lo0020 & ~lo0981 ;
  assign new_n16545 = ~new_n16543 & ~new_n16544 ;
  assign new_n16546 = ~lo0040 & lo0990 ;
  assign new_n16547 = lo0032 & ~lo1026 ;
  assign new_n16548 = ~new_n16546 & ~new_n16547 ;
  assign new_n16549 = new_n16545 & new_n16548 ;
  assign new_n16550 = ~lo0042 & lo0986 ;
  assign new_n16551 = lo0029 & ~lo0983 ;
  assign new_n16552 = ~new_n16550 & ~new_n16551 ;
  assign new_n16553 = ~lo0020 & lo0981 ;
  assign new_n16554 = lo0042 & ~lo0986 ;
  assign new_n16555 = ~new_n16553 & ~new_n16554 ;
  assign new_n16556 = new_n16552 & new_n16555 ;
  assign new_n16557 = new_n16549 & new_n16556 ;
  assign new_n16558 = ~lo0022 & lo1049 ;
  assign new_n16559 = lo1020 & ~lo1059 ;
  assign new_n16560 = ~new_n16558 & ~new_n16559 ;
  assign new_n16561 = ~lo0038 & lo0919 ;
  assign new_n16562 = lo0022 & ~lo1049 ;
  assign new_n16563 = ~new_n16561 & ~new_n16562 ;
  assign new_n16564 = new_n16560 & new_n16563 ;
  assign new_n16565 = ~lo0030 & lo0929 ;
  assign new_n16566 = lo0040 & ~lo0990 ;
  assign new_n16567 = ~new_n16565 & ~new_n16566 ;
  assign new_n16568 = ~lo1020 & lo1059 ;
  assign new_n16569 = lo0030 & ~lo0929 ;
  assign new_n16570 = ~new_n16568 & ~new_n16569 ;
  assign new_n16571 = new_n16567 & new_n16570 ;
  assign new_n16572 = new_n16564 & new_n16571 ;
  assign new_n16573 = new_n16557 & new_n16572 ;
  assign new_n16574 = new_n16542 & new_n16573 ;
  assign new_n16575 = lo0024 & ~lo0975 ;
  assign new_n16576 = lo0892 & ~lo1044 ;
  assign new_n16577 = ~new_n16575 & ~new_n16576 ;
  assign new_n16578 = lo1036 & ~lo1056 ;
  assign new_n16579 = ~lo1036 & lo1056 ;
  assign new_n16580 = ~new_n16578 & ~new_n16579 ;
  assign new_n16581 = new_n16577 & new_n16580 ;
  assign new_n16582 = ~lo0994 & lo1057 ;
  assign new_n16583 = lo0023 & ~lo0921 ;
  assign new_n16584 = ~new_n16582 & ~new_n16583 ;
  assign new_n16585 = ~lo0892 & lo1044 ;
  assign new_n16586 = lo0994 & ~lo1057 ;
  assign new_n16587 = ~new_n16585 & ~new_n16586 ;
  assign new_n16588 = new_n16584 & new_n16587 ;
  assign new_n16589 = new_n16581 & new_n16588 ;
  assign new_n16590 = ~lo0024 & lo0975 ;
  assign new_n16591 = lo0041 & ~lo1015 ;
  assign new_n16592 = ~lo0041 & lo1015 ;
  assign new_n16593 = ~new_n16591 & ~new_n16592 ;
  assign new_n16594 = ~new_n16590 & new_n16593 ;
  assign new_n16595 = new_n16483 & new_n16594 ;
  assign new_n16596 = new_n16589 & new_n16595 ;
  assign new_n16597 = ~lo0036 & lo1008 ;
  assign new_n16598 = lo0025 & ~lo1013 ;
  assign new_n16599 = ~new_n16597 & ~new_n16598 ;
  assign new_n16600 = ~lo0035 & lo0970 ;
  assign new_n16601 = lo0036 & ~lo1008 ;
  assign new_n16602 = ~new_n16600 & ~new_n16601 ;
  assign new_n16603 = new_n16599 & new_n16602 ;
  assign new_n16604 = ~lo0028 & lo0992 ;
  assign new_n16605 = lo0922 & ~lo1058 ;
  assign new_n16606 = ~new_n16604 & ~new_n16605 ;
  assign new_n16607 = ~lo0025 & lo1013 ;
  assign new_n16608 = lo0028 & ~lo0992 ;
  assign new_n16609 = ~new_n16607 & ~new_n16608 ;
  assign new_n16610 = new_n16606 & new_n16609 ;
  assign new_n16611 = new_n16603 & new_n16610 ;
  assign new_n16612 = ~lo0039 & lo0973 ;
  assign new_n16613 = lo0019 & ~lo0927 ;
  assign new_n16614 = ~new_n16612 & ~new_n16613 ;
  assign new_n16615 = ~lo0023 & lo0921 ;
  assign new_n16616 = lo0039 & ~lo0973 ;
  assign new_n16617 = ~new_n16615 & ~new_n16616 ;
  assign new_n16618 = new_n16614 & new_n16617 ;
  assign new_n16619 = ~lo0917 & lo1003 ;
  assign new_n16620 = lo0035 & ~lo0970 ;
  assign new_n16621 = ~new_n16619 & ~new_n16620 ;
  assign new_n16622 = ~lo0019 & lo0927 ;
  assign new_n16623 = lo0917 & ~lo1003 ;
  assign new_n16624 = ~new_n16622 & ~new_n16623 ;
  assign new_n16625 = new_n16621 & new_n16624 ;
  assign new_n16626 = new_n16618 & new_n16625 ;
  assign new_n16627 = new_n16611 & new_n16626 ;
  assign new_n16628 = ~lo0033 & lo1000 ;
  assign new_n16629 = lo0034 & ~lo1041 ;
  assign new_n16630 = ~new_n16628 & ~new_n16629 ;
  assign new_n16631 = ~lo0027 & lo0988 ;
  assign new_n16632 = lo0033 & ~lo1000 ;
  assign new_n16633 = ~new_n16631 & ~new_n16632 ;
  assign new_n16634 = new_n16630 & new_n16633 ;
  assign new_n16635 = ~lo0893 & lo1028 ;
  assign new_n16636 = lo0038 & ~lo0919 ;
  assign new_n16637 = ~new_n16635 & ~new_n16636 ;
  assign new_n16638 = ~lo0034 & lo1041 ;
  assign new_n16639 = lo0893 & ~lo1028 ;
  assign new_n16640 = ~new_n16638 & ~new_n16639 ;
  assign new_n16641 = new_n16637 & new_n16640 ;
  assign new_n16642 = new_n16634 & new_n16641 ;
  assign new_n16643 = ~lo0037 & lo1033 ;
  assign new_n16644 = lo0026 & ~lo1017 ;
  assign new_n16645 = ~new_n16643 & ~new_n16644 ;
  assign new_n16646 = ~lo0922 & lo1058 ;
  assign new_n16647 = lo0037 & ~lo1033 ;
  assign new_n16648 = ~new_n16646 & ~new_n16647 ;
  assign new_n16649 = new_n16645 & new_n16648 ;
  assign new_n16650 = ~lo0021 & lo1011 ;
  assign new_n16651 = lo0027 & ~lo0988 ;
  assign new_n16652 = ~new_n16650 & ~new_n16651 ;
  assign new_n16653 = ~lo0026 & lo1017 ;
  assign new_n16654 = lo0021 & ~lo1011 ;
  assign new_n16655 = ~new_n16653 & ~new_n16654 ;
  assign new_n16656 = new_n16652 & new_n16655 ;
  assign new_n16657 = new_n16649 & new_n16656 ;
  assign new_n16658 = new_n16642 & new_n16657 ;
  assign new_n16659 = new_n16627 & new_n16658 ;
  assign new_n16660 = new_n16596 & new_n16659 ;
  assign new_n16661 = new_n16574 & new_n16660 ;
  assign new_n16662 = ~new_n16532 & ~new_n16661 ;
  assign new_n16663 = ~new_n16531 & new_n16662 ;
  assign new_n16664 = new_n12358 & new_n15372 ;
  assign new_n16665 = new_n2465 & new_n12910 ;
  assign new_n16666 = new_n16664 & new_n16665 ;
  assign new_n16667 = ~lo0858 & ~lo0859 ;
  assign new_n16668 = ~new_n16666 & new_n16667 ;
  assign new_n16669 = ~new_n2252 & ~new_n16668 ;
  assign new_n16670 = ~new_n15375 & ~new_n16669 ;
  assign new_n16671 = lo0181 & new_n16670 ;
  assign new_n16672 = lo0954 & new_n11591 ;
  assign new_n16673 = new_n11591 & ~new_n16672 ;
  assign new_n16674 = ~new_n8446 & ~new_n16673 ;
  assign new_n16675 = ~lo0954 & new_n8446 ;
  assign new_n16676 = ~new_n11591 & new_n16675 ;
  assign new_n16677 = ~new_n16674 & ~new_n16676 ;
  assign new_n16678 = lo0859 & ~new_n16677 ;
  assign new_n16679 = ~lo0859 & ~new_n5743 ;
  assign new_n16680 = ~new_n16678 & ~new_n16679 ;
  assign new_n16681 = ~new_n16666 & ~new_n16680 ;
  assign new_n16682 = lo1062 & new_n16666 ;
  assign new_n16683 = ~new_n15375 & ~new_n16682 ;
  assign new_n16684 = ~new_n16681 & new_n16683 ;
  assign new_n16685 = ~new_n16670 & ~new_n16684 ;
  assign new_n16686 = ~new_n16671 & ~new_n16685 ;
  assign new_n16687 = lo0044 & new_n16480 ;
  assign new_n16688 = lo0182 & ~new_n16687 ;
  assign new_n16689 = lo1444 & new_n16687 ;
  assign new_n16690 = ~new_n16688 & ~new_n16689 ;
  assign new_n16691 = lo0183 & new_n16670 ;
  assign new_n16692 = lo0954 & new_n11639 ;
  assign new_n16693 = new_n11639 & ~new_n16692 ;
  assign new_n16694 = ~new_n8572 & ~new_n16693 ;
  assign new_n16695 = ~lo0954 & new_n8572 ;
  assign new_n16696 = ~new_n11639 & new_n16695 ;
  assign new_n16697 = ~new_n16694 & ~new_n16696 ;
  assign new_n16698 = lo0859 & ~new_n16697 ;
  assign new_n16699 = ~lo0859 & new_n5977 ;
  assign new_n16700 = ~new_n16698 & ~new_n16699 ;
  assign new_n16701 = ~new_n16666 & ~new_n16700 ;
  assign new_n16702 = lo1063 & new_n16666 ;
  assign new_n16703 = ~new_n15375 & ~new_n16702 ;
  assign new_n16704 = ~new_n16701 & new_n16703 ;
  assign new_n16705 = ~new_n16670 & ~new_n16704 ;
  assign new_n16706 = ~new_n16691 & ~new_n16705 ;
  assign new_n16707 = lo0184 & ~new_n16687 ;
  assign new_n16708 = lo1445 & new_n16687 ;
  assign new_n16709 = ~new_n16707 & ~new_n16708 ;
  assign new_n16710 = lo0185 & new_n16670 ;
  assign new_n16711 = lo0954 & new_n11690 ;
  assign new_n16712 = new_n11690 & ~new_n16711 ;
  assign new_n16713 = ~new_n8693 & ~new_n16712 ;
  assign new_n16714 = ~lo0954 & new_n8693 ;
  assign new_n16715 = ~new_n11690 & new_n16714 ;
  assign new_n16716 = ~new_n16713 & ~new_n16715 ;
  assign new_n16717 = lo0859 & ~new_n16716 ;
  assign new_n16718 = ~lo0859 & new_n6202 ;
  assign new_n16719 = ~new_n16717 & ~new_n16718 ;
  assign new_n16720 = ~new_n16666 & ~new_n16719 ;
  assign new_n16721 = lo1064 & new_n16666 ;
  assign new_n16722 = ~new_n15375 & ~new_n16721 ;
  assign new_n16723 = ~new_n16720 & new_n16722 ;
  assign new_n16724 = ~new_n16670 & ~new_n16723 ;
  assign new_n16725 = ~new_n16710 & ~new_n16724 ;
  assign new_n16726 = lo0186 & ~new_n16687 ;
  assign new_n16727 = lo1446 & new_n16687 ;
  assign new_n16728 = ~new_n16726 & ~new_n16727 ;
  assign new_n16729 = lo0187 & new_n16670 ;
  assign new_n16730 = lo0954 & new_n11840 ;
  assign new_n16731 = new_n11840 & ~new_n16730 ;
  assign new_n16732 = ~new_n8815 & ~new_n16731 ;
  assign new_n16733 = ~lo0954 & new_n8815 ;
  assign new_n16734 = ~new_n11840 & new_n16733 ;
  assign new_n16735 = ~new_n16732 & ~new_n16734 ;
  assign new_n16736 = lo0859 & ~new_n16735 ;
  assign new_n16737 = ~lo0859 & new_n6433 ;
  assign new_n16738 = ~new_n16736 & ~new_n16737 ;
  assign new_n16739 = ~new_n16666 & ~new_n16738 ;
  assign new_n16740 = lo1065 & new_n16666 ;
  assign new_n16741 = ~new_n15375 & ~new_n16740 ;
  assign new_n16742 = ~new_n16739 & new_n16741 ;
  assign new_n16743 = ~new_n16670 & ~new_n16742 ;
  assign new_n16744 = ~new_n16729 & ~new_n16743 ;
  assign new_n16745 = lo0188 & ~new_n16687 ;
  assign new_n16746 = lo1284 & new_n16687 ;
  assign new_n16747 = ~new_n16745 & ~new_n16746 ;
  assign new_n16748 = lo0189 & ~new_n15612 ;
  assign new_n16749 = ~new_n2448 & new_n15612 ;
  assign new_n16750 = ~new_n16748 & ~new_n16749 ;
  assign new_n16751 = lo0190 & ~new_n15612 ;
  assign new_n16752 = ~new_n2452 & new_n15612 ;
  assign new_n16753 = ~new_n16751 & ~new_n16752 ;
  assign new_n16754 = lo0191 & ~new_n15612 ;
  assign new_n16755 = ~new_n12327 & new_n15612 ;
  assign new_n16756 = ~new_n16754 & ~new_n16755 ;
  assign new_n16757 = lo0192 & ~new_n15612 ;
  assign new_n16758 = new_n12355 & new_n15612 ;
  assign new_n16759 = ~new_n16757 & ~new_n16758 ;
  assign new_n16760 = lo0193 & ~new_n15612 ;
  assign new_n16761 = ~new_n12322 & new_n15612 ;
  assign new_n16762 = ~new_n16760 & ~new_n16761 ;
  assign new_n16763 = lo0194 & ~new_n15612 ;
  assign new_n16764 = ~new_n2463 & new_n15612 ;
  assign new_n16765 = ~new_n16763 & ~new_n16764 ;
  assign new_n16766 = lo0195 & ~new_n15612 ;
  assign new_n16767 = ~new_n12364 & new_n15612 ;
  assign new_n16768 = ~new_n16766 & ~new_n16767 ;
  assign new_n16769 = lo0196 & new_n2252 ;
  assign new_n16770 = ~new_n2252 & ~new_n12675 ;
  assign new_n16771 = ~new_n16769 & ~new_n16770 ;
  assign new_n16772 = lo0197 & new_n2252 ;
  assign new_n16773 = ~new_n2252 & ~new_n12589 ;
  assign new_n16774 = ~new_n16772 & ~new_n16773 ;
  assign new_n16775 = lo0198 & new_n2252 ;
  assign new_n16776 = ~new_n2252 & ~new_n12834 ;
  assign new_n16777 = ~new_n16775 & ~new_n16776 ;
  assign new_n16778 = lo0199 & new_n2252 ;
  assign new_n16779 = ~new_n2252 & ~new_n12928 ;
  assign new_n16780 = ~new_n16778 & ~new_n16779 ;
  assign new_n16781 = lo0200 & new_n2252 ;
  assign new_n16782 = ~new_n2252 & ~new_n12729 ;
  assign new_n16783 = ~new_n16781 & ~new_n16782 ;
  assign new_n16784 = lo0201 & ~new_n15033 ;
  assign new_n16785 = new_n6433 & ~new_n15036 ;
  assign new_n16786 = new_n15036 & ~new_n16735 ;
  assign new_n16787 = ~new_n16785 & ~new_n16786 ;
  assign new_n16788 = new_n15033 & ~new_n16787 ;
  assign new_n16789 = ~new_n16784 & ~new_n16788 ;
  assign new_n16790 = lo0202 & ~new_n14848 ;
  assign new_n16791 = new_n6433 & ~new_n14853 ;
  assign new_n16792 = new_n14853 & ~new_n16735 ;
  assign new_n16793 = ~new_n16791 & ~new_n16792 ;
  assign new_n16794 = new_n14848 & ~new_n16793 ;
  assign new_n16795 = ~new_n16790 & ~new_n16794 ;
  assign new_n16796 = lo0203 & ~new_n14869 ;
  assign new_n16797 = new_n6433 & ~new_n14872 ;
  assign new_n16798 = new_n14872 & ~new_n16735 ;
  assign new_n16799 = ~new_n16797 & ~new_n16798 ;
  assign new_n16800 = new_n14869 & ~new_n16799 ;
  assign new_n16801 = ~new_n16796 & ~new_n16800 ;
  assign new_n16802 = lo0204 & ~new_n14886 ;
  assign new_n16803 = new_n6433 & ~new_n14889 ;
  assign new_n16804 = new_n14889 & ~new_n16735 ;
  assign new_n16805 = ~new_n16803 & ~new_n16804 ;
  assign new_n16806 = new_n14886 & ~new_n16805 ;
  assign new_n16807 = ~new_n16802 & ~new_n16806 ;
  assign new_n16808 = lo0205 & ~new_n14903 ;
  assign new_n16809 = new_n6433 & ~new_n14906 ;
  assign new_n16810 = new_n14906 & ~new_n16735 ;
  assign new_n16811 = ~new_n16809 & ~new_n16810 ;
  assign new_n16812 = new_n14903 & ~new_n16811 ;
  assign new_n16813 = ~new_n16808 & ~new_n16812 ;
  assign new_n16814 = lo0206 & ~new_n14924 ;
  assign new_n16815 = new_n6433 & ~new_n14927 ;
  assign new_n16816 = new_n14927 & ~new_n16735 ;
  assign new_n16817 = ~new_n16815 & ~new_n16816 ;
  assign new_n16818 = new_n14924 & ~new_n16817 ;
  assign new_n16819 = ~new_n16814 & ~new_n16818 ;
  assign new_n16820 = lo0207 & ~new_n14943 ;
  assign new_n16821 = new_n6433 & ~new_n14946 ;
  assign new_n16822 = new_n14946 & ~new_n16735 ;
  assign new_n16823 = ~new_n16821 & ~new_n16822 ;
  assign new_n16824 = new_n14943 & ~new_n16823 ;
  assign new_n16825 = ~new_n16820 & ~new_n16824 ;
  assign new_n16826 = lo0208 & ~new_n14960 ;
  assign new_n16827 = new_n6433 & ~new_n14963 ;
  assign new_n16828 = new_n14963 & ~new_n16735 ;
  assign new_n16829 = ~new_n16827 & ~new_n16828 ;
  assign new_n16830 = new_n14960 & ~new_n16829 ;
  assign new_n16831 = ~new_n16826 & ~new_n16830 ;
  assign new_n16832 = lo0209 & ~new_n14977 ;
  assign new_n16833 = new_n6433 & ~new_n14980 ;
  assign new_n16834 = new_n14980 & ~new_n16735 ;
  assign new_n16835 = ~new_n16833 & ~new_n16834 ;
  assign new_n16836 = new_n14977 & ~new_n16835 ;
  assign new_n16837 = ~new_n16832 & ~new_n16836 ;
  assign new_n16838 = lo0210 & ~new_n14997 ;
  assign new_n16839 = new_n6433 & ~new_n15000 ;
  assign new_n16840 = new_n15000 & ~new_n16735 ;
  assign new_n16841 = ~new_n16839 & ~new_n16840 ;
  assign new_n16842 = new_n14997 & ~new_n16841 ;
  assign new_n16843 = ~new_n16838 & ~new_n16842 ;
  assign new_n16844 = lo0211 & ~new_n15016 ;
  assign new_n16845 = new_n6433 & ~new_n15019 ;
  assign new_n16846 = new_n15019 & ~new_n16735 ;
  assign new_n16847 = ~new_n16845 & ~new_n16846 ;
  assign new_n16848 = new_n15016 & ~new_n16847 ;
  assign new_n16849 = ~new_n16844 & ~new_n16848 ;
  assign new_n16850 = lo0212 & ~new_n15050 ;
  assign new_n16851 = new_n6433 & ~new_n15053 ;
  assign new_n16852 = new_n15053 & ~new_n16735 ;
  assign new_n16853 = ~new_n16851 & ~new_n16852 ;
  assign new_n16854 = new_n15050 & ~new_n16853 ;
  assign new_n16855 = ~new_n16850 & ~new_n16854 ;
  assign new_n16856 = lo0213 & ~new_n15071 ;
  assign new_n16857 = new_n6433 & ~new_n15074 ;
  assign new_n16858 = new_n15074 & ~new_n16735 ;
  assign new_n16859 = ~new_n16857 & ~new_n16858 ;
  assign new_n16860 = new_n15071 & ~new_n16859 ;
  assign new_n16861 = ~new_n16856 & ~new_n16860 ;
  assign new_n16862 = lo0214 & ~new_n15090 ;
  assign new_n16863 = new_n6433 & ~new_n15093 ;
  assign new_n16864 = new_n15093 & ~new_n16735 ;
  assign new_n16865 = ~new_n16863 & ~new_n16864 ;
  assign new_n16866 = new_n15090 & ~new_n16865 ;
  assign new_n16867 = ~new_n16862 & ~new_n16866 ;
  assign new_n16868 = lo0215 & ~new_n15107 ;
  assign new_n16869 = new_n6433 & ~new_n15110 ;
  assign new_n16870 = new_n15110 & ~new_n16735 ;
  assign new_n16871 = ~new_n16869 & ~new_n16870 ;
  assign new_n16872 = new_n15107 & ~new_n16871 ;
  assign new_n16873 = ~new_n16868 & ~new_n16872 ;
  assign new_n16874 = lo0216 & ~new_n15124 ;
  assign new_n16875 = new_n6433 & ~new_n15127 ;
  assign new_n16876 = new_n15127 & ~new_n16735 ;
  assign new_n16877 = ~new_n16875 & ~new_n16876 ;
  assign new_n16878 = new_n15124 & ~new_n16877 ;
  assign new_n16879 = ~new_n16874 & ~new_n16878 ;
  assign new_n16880 = lo0217 & ~new_n15137 ;
  assign new_n16881 = new_n15137 & ~new_n16175 ;
  assign new_n16882 = ~new_n16880 & ~new_n16881 ;
  assign new_n16883 = lo0218 & ~new_n15137 ;
  assign new_n16884 = new_n15137 & ~new_n16398 ;
  assign new_n16885 = ~new_n16883 & ~new_n16884 ;
  assign new_n16886 = lo0219 & ~new_n15137 ;
  assign new_n16887 = new_n15137 & ~new_n16153 ;
  assign new_n16888 = ~new_n16886 & ~new_n16887 ;
  assign new_n16889 = lo0220 & ~new_n15137 ;
  assign new_n16890 = new_n15137 & ~new_n16371 ;
  assign new_n16891 = ~new_n16889 & ~new_n16890 ;
  assign new_n16892 = lo0221 & new_n2252 ;
  assign new_n16893 = ~new_n2252 & ~new_n12420 ;
  assign new_n16894 = ~new_n16892 & ~new_n16893 ;
  assign new_n16895 = lo0222 & new_n2252 ;
  assign new_n16896 = ~new_n12329 & ~new_n15469 ;
  assign new_n16897 = new_n12325 & new_n15644 ;
  assign new_n16898 = new_n13286 & new_n16897 ;
  assign new_n16899 = new_n2454 & new_n16898 ;
  assign new_n16900 = ~new_n16896 & ~new_n16899 ;
  assign new_n16901 = ~new_n12698 & ~new_n12768 ;
  assign new_n16902 = ~new_n2252 & new_n16901 ;
  assign new_n16903 = ~new_n16900 & new_n16902 ;
  assign new_n16904 = ~new_n16895 & ~new_n16903 ;
  assign new_n16905 = lo0223 & new_n2252 ;
  assign new_n16906 = ~new_n16510 & ~new_n16905 ;
  assign new_n16907 = lo0224 & new_n2252 ;
  assign new_n16908 = ~new_n2252 & ~new_n12460 ;
  assign new_n16909 = ~new_n16907 & ~new_n16908 ;
  assign new_n16910 = lo0225 & ~new_n15365 ;
  assign new_n16911 = lo0952 & ~new_n16735 ;
  assign new_n16912 = ~lo0952 & new_n6433 ;
  assign new_n16913 = ~new_n16911 & ~new_n16912 ;
  assign new_n16914 = new_n15365 & ~new_n16913 ;
  assign new_n16915 = ~new_n16910 & ~new_n16914 ;
  assign new_n16916 = lo0226 & new_n15454 ;
  assign new_n16917 = lo0958 & ~new_n16735 ;
  assign new_n16918 = lo0226 & ~new_n13945 ;
  assign new_n16919 = ~lo0226 & new_n13945 ;
  assign new_n16920 = ~new_n16918 & ~new_n16919 ;
  assign new_n16921 = ~lo0958 & ~new_n16920 ;
  assign new_n16922 = ~new_n16917 & ~new_n16921 ;
  assign new_n16923 = ~new_n15454 & ~new_n16922 ;
  assign new_n16924 = ~new_n16916 & ~new_n16923 ;
  assign new_n16925 = lo0227 & ~new_n15033 ;
  assign new_n16926 = new_n4257 & ~new_n15036 ;
  assign new_n16927 = ~new_n14366 & new_n15036 ;
  assign new_n16928 = ~new_n16926 & ~new_n16927 ;
  assign new_n16929 = new_n15033 & ~new_n16928 ;
  assign new_n16930 = ~new_n16925 & ~new_n16929 ;
  assign new_n16931 = lo0228 & new_n2252 ;
  assign new_n16932 = ~new_n2252 & new_n12506 ;
  assign new_n16933 = new_n2455 & new_n16932 ;
  assign new_n16934 = new_n15644 & new_n16933 ;
  assign new_n16935 = ~new_n16931 & ~new_n16934 ;
  assign new_n16936 = lo0229 & new_n2252 ;
  assign new_n16937 = ~new_n2252 & ~new_n12357 ;
  assign new_n16938 = ~new_n16936 & ~new_n16937 ;
  assign new_n16939 = lo0230 & ~new_n14924 ;
  assign new_n16940 = new_n4257 & ~new_n14927 ;
  assign new_n16941 = ~new_n14366 & new_n14927 ;
  assign new_n16942 = ~new_n16940 & ~new_n16941 ;
  assign new_n16943 = new_n14924 & ~new_n16942 ;
  assign new_n16944 = ~new_n16939 & ~new_n16943 ;
  assign new_n16945 = lo0231 & ~new_n14869 ;
  assign new_n16946 = new_n4257 & ~new_n14872 ;
  assign new_n16947 = ~new_n14366 & new_n14872 ;
  assign new_n16948 = ~new_n16946 & ~new_n16947 ;
  assign new_n16949 = new_n14869 & ~new_n16948 ;
  assign new_n16950 = ~new_n16945 & ~new_n16949 ;
  assign new_n16951 = lo0232 & ~new_n15016 ;
  assign new_n16952 = new_n4257 & ~new_n15019 ;
  assign new_n16953 = ~new_n14366 & new_n15019 ;
  assign new_n16954 = ~new_n16952 & ~new_n16953 ;
  assign new_n16955 = new_n15016 & ~new_n16954 ;
  assign new_n16956 = ~new_n16951 & ~new_n16955 ;
  assign new_n16957 = lo0233 & ~new_n15071 ;
  assign new_n16958 = new_n4257 & ~new_n15074 ;
  assign new_n16959 = ~new_n14366 & new_n15074 ;
  assign new_n16960 = ~new_n16958 & ~new_n16959 ;
  assign new_n16961 = new_n15071 & ~new_n16960 ;
  assign new_n16962 = ~new_n16957 & ~new_n16961 ;
  assign new_n16963 = lo0234 & ~new_n14848 ;
  assign new_n16964 = new_n4257 & ~new_n14853 ;
  assign new_n16965 = ~new_n14366 & new_n14853 ;
  assign new_n16966 = ~new_n16964 & ~new_n16965 ;
  assign new_n16967 = new_n14848 & ~new_n16966 ;
  assign new_n16968 = ~new_n16963 & ~new_n16967 ;
  assign new_n16969 = lo0235 & ~new_n14943 ;
  assign new_n16970 = new_n4257 & ~new_n14946 ;
  assign new_n16971 = ~new_n14366 & new_n14946 ;
  assign new_n16972 = ~new_n16970 & ~new_n16971 ;
  assign new_n16973 = new_n14943 & ~new_n16972 ;
  assign new_n16974 = ~new_n16969 & ~new_n16973 ;
  assign new_n16975 = lo0236 & ~new_n14997 ;
  assign new_n16976 = new_n4257 & ~new_n15000 ;
  assign new_n16977 = ~new_n14366 & new_n15000 ;
  assign new_n16978 = ~new_n16976 & ~new_n16977 ;
  assign new_n16979 = new_n14997 & ~new_n16978 ;
  assign new_n16980 = ~new_n16975 & ~new_n16979 ;
  assign new_n16981 = lo0237 & ~new_n15090 ;
  assign new_n16982 = new_n4257 & ~new_n15093 ;
  assign new_n16983 = ~new_n14366 & new_n15093 ;
  assign new_n16984 = ~new_n16982 & ~new_n16983 ;
  assign new_n16985 = new_n15090 & ~new_n16984 ;
  assign new_n16986 = ~new_n16981 & ~new_n16985 ;
  assign new_n16987 = lo0238 & ~new_n14886 ;
  assign new_n16988 = new_n4257 & ~new_n14889 ;
  assign new_n16989 = ~new_n14366 & new_n14889 ;
  assign new_n16990 = ~new_n16988 & ~new_n16989 ;
  assign new_n16991 = new_n14886 & ~new_n16990 ;
  assign new_n16992 = ~new_n16987 & ~new_n16991 ;
  assign new_n16993 = lo0239 & ~new_n14960 ;
  assign new_n16994 = new_n4257 & ~new_n14963 ;
  assign new_n16995 = ~new_n14366 & new_n14963 ;
  assign new_n16996 = ~new_n16994 & ~new_n16995 ;
  assign new_n16997 = new_n14960 & ~new_n16996 ;
  assign new_n16998 = ~new_n16993 & ~new_n16997 ;
  assign new_n16999 = lo0240 & ~new_n15107 ;
  assign new_n17000 = new_n4257 & ~new_n15110 ;
  assign new_n17001 = ~new_n14366 & new_n15110 ;
  assign new_n17002 = ~new_n17000 & ~new_n17001 ;
  assign new_n17003 = new_n15107 & ~new_n17002 ;
  assign new_n17004 = ~new_n16999 & ~new_n17003 ;
  assign new_n17005 = lo0241 & ~new_n14977 ;
  assign new_n17006 = new_n4257 & ~new_n14980 ;
  assign new_n17007 = ~new_n14366 & new_n14980 ;
  assign new_n17008 = ~new_n17006 & ~new_n17007 ;
  assign new_n17009 = new_n14977 & ~new_n17008 ;
  assign new_n17010 = ~new_n17005 & ~new_n17009 ;
  assign new_n17011 = lo0242 & ~new_n14903 ;
  assign new_n17012 = new_n4257 & ~new_n14906 ;
  assign new_n17013 = ~new_n14366 & new_n14906 ;
  assign new_n17014 = ~new_n17012 & ~new_n17013 ;
  assign new_n17015 = new_n14903 & ~new_n17014 ;
  assign new_n17016 = ~new_n17011 & ~new_n17015 ;
  assign new_n17017 = lo0243 & ~new_n15050 ;
  assign new_n17018 = new_n4257 & ~new_n15053 ;
  assign new_n17019 = ~new_n14366 & new_n15053 ;
  assign new_n17020 = ~new_n17018 & ~new_n17019 ;
  assign new_n17021 = new_n15050 & ~new_n17020 ;
  assign new_n17022 = ~new_n17017 & ~new_n17021 ;
  assign new_n17023 = lo0244 & ~new_n15124 ;
  assign new_n17024 = new_n4257 & ~new_n15127 ;
  assign new_n17025 = ~new_n14366 & new_n15127 ;
  assign new_n17026 = ~new_n17024 & ~new_n17025 ;
  assign new_n17027 = new_n15124 & ~new_n17026 ;
  assign new_n17028 = ~new_n17023 & ~new_n17027 ;
  assign new_n17029 = lo0245 & new_n15454 ;
  assign new_n17030 = lo0958 & ~new_n14366 ;
  assign new_n17031 = ~lo0958 & ~new_n14369 ;
  assign new_n17032 = ~new_n17030 & ~new_n17031 ;
  assign new_n17033 = ~new_n15454 & ~new_n17032 ;
  assign new_n17034 = ~new_n17029 & ~new_n17033 ;
  assign new_n17035 = lo0246 & ~new_n15365 ;
  assign new_n17036 = lo0952 & ~new_n14366 ;
  assign new_n17037 = ~lo0952 & new_n4257 ;
  assign new_n17038 = ~new_n17036 & ~new_n17037 ;
  assign new_n17039 = new_n15365 & ~new_n17038 ;
  assign new_n17040 = ~new_n17035 & ~new_n17039 ;
  assign new_n17041 = lo0247 & new_n2252 ;
  assign new_n17042 = ~new_n2252 & ~new_n13574 ;
  assign new_n17043 = ~new_n17041 & ~new_n17042 ;
  assign new_n17044 = lo0248 & new_n2252 ;
  assign new_n17045 = ~new_n12329 & new_n15451 ;
  assign new_n17046 = new_n2446 & new_n12523 ;
  assign new_n17047 = new_n12745 & new_n17046 ;
  assign new_n17048 = ~new_n2446 & new_n12370 ;
  assign new_n17049 = ~new_n17047 & ~new_n17048 ;
  assign new_n17050 = ~new_n2252 & new_n12376 ;
  assign new_n17051 = new_n2455 & new_n17050 ;
  assign new_n17052 = ~new_n17049 & new_n17051 ;
  assign new_n17053 = new_n17045 & new_n17052 ;
  assign new_n17054 = ~new_n17044 & ~new_n17053 ;
  assign new_n17055 = lo0249 & ~new_n14699 ;
  assign new_n17056 = ~new_n13508 & new_n14699 ;
  assign new_n17057 = ~new_n17055 & ~new_n17056 ;
  assign new_n17058 = lo0250 & ~new_n14699 ;
  assign new_n17059 = ~new_n13702 & new_n14699 ;
  assign new_n17060 = ~new_n17058 & ~new_n17059 ;
  assign new_n17061 = lo0251 & ~new_n14699 ;
  assign new_n17062 = ~new_n13617 & new_n14699 ;
  assign new_n17063 = ~new_n17061 & ~new_n17062 ;
  assign new_n17064 = lo0252 & ~new_n14699 ;
  assign new_n17065 = ~new_n13662 & new_n14699 ;
  assign new_n17066 = ~new_n17064 & ~new_n17065 ;
  assign new_n17067 = lo0253 & new_n2252 ;
  assign new_n17068 = new_n12395 & new_n12472 ;
  assign new_n17069 = new_n12325 & new_n12471 ;
  assign new_n17070 = ~new_n17068 & ~new_n17069 ;
  assign new_n17071 = new_n16475 & ~new_n17070 ;
  assign new_n17072 = new_n15451 & new_n17071 ;
  assign new_n17073 = ~new_n17067 & ~new_n17072 ;
  assign new_n17074 = lo0254 & new_n2252 ;
  assign new_n17075 = new_n2264 & new_n12370 ;
  assign new_n17076 = ~new_n12863 & ~new_n17075 ;
  assign new_n17077 = new_n15348 & ~new_n17076 ;
  assign new_n17078 = ~new_n17074 & ~new_n17077 ;
  assign new_n17079 = lo0255 & new_n2252 ;
  assign new_n17080 = ~new_n2252 & new_n12860 ;
  assign new_n17081 = new_n16664 & new_n17080 ;
  assign new_n17082 = ~new_n17079 & ~new_n17081 ;
  assign new_n17083 = lo0256 & new_n2252 ;
  assign new_n17084 = new_n12522 & new_n14742 ;
  assign new_n17085 = new_n2446 & new_n13768 ;
  assign new_n17086 = ~new_n2446 & new_n12507 ;
  assign new_n17087 = ~new_n17085 & ~new_n17086 ;
  assign new_n17088 = new_n12329 & ~new_n17087 ;
  assign new_n17089 = ~new_n17084 & ~new_n17088 ;
  assign new_n17090 = new_n2455 & ~new_n17089 ;
  assign new_n17091 = new_n12405 & new_n15442 ;
  assign new_n17092 = ~new_n12402 & ~new_n17091 ;
  assign new_n17093 = ~new_n17090 & new_n17092 ;
  assign new_n17094 = new_n2454 & ~new_n17093 ;
  assign new_n17095 = ~new_n2454 & new_n17093 ;
  assign new_n17096 = ~new_n17094 & ~new_n17095 ;
  assign new_n17097 = ~new_n2446 & ~new_n17096 ;
  assign new_n17098 = new_n2446 & new_n17094 ;
  assign new_n17099 = new_n12357 & new_n12395 ;
  assign new_n17100 = ~new_n12329 & new_n17099 ;
  assign new_n17101 = new_n2264 & ~new_n2454 ;
  assign new_n17102 = ~new_n2446 & new_n17101 ;
  assign new_n17103 = ~new_n17100 & new_n17102 ;
  assign new_n17104 = ~new_n17093 & new_n17103 ;
  assign new_n17105 = ~new_n17098 & ~new_n17104 ;
  assign new_n17106 = ~new_n17097 & new_n17105 ;
  assign new_n17107 = ~new_n2252 & ~new_n17106 ;
  assign new_n17108 = ~new_n17083 & ~new_n17107 ;
  assign new_n17109 = lo0257 & new_n2252 ;
  assign new_n17110 = ~new_n2252 & new_n14813 ;
  assign new_n17111 = ~new_n17109 & ~new_n17110 ;
  assign new_n17112 = lo0258 & ~new_n14943 ;
  assign new_n17113 = new_n3538 & ~new_n14946 ;
  assign new_n17114 = ~new_n14313 & new_n14946 ;
  assign new_n17115 = ~new_n17113 & ~new_n17114 ;
  assign new_n17116 = new_n14943 & ~new_n17115 ;
  assign new_n17117 = ~new_n17112 & ~new_n17116 ;
  assign new_n17118 = lo0259 & ~new_n14848 ;
  assign new_n17119 = new_n3538 & ~new_n14853 ;
  assign new_n17120 = ~new_n14313 & new_n14853 ;
  assign new_n17121 = ~new_n17119 & ~new_n17120 ;
  assign new_n17122 = new_n14848 & ~new_n17121 ;
  assign new_n17123 = ~new_n17118 & ~new_n17122 ;
  assign new_n17124 = lo0260 & ~new_n14997 ;
  assign new_n17125 = new_n3538 & ~new_n15000 ;
  assign new_n17126 = ~new_n14313 & new_n15000 ;
  assign new_n17127 = ~new_n17125 & ~new_n17126 ;
  assign new_n17128 = new_n14997 & ~new_n17127 ;
  assign new_n17129 = ~new_n17124 & ~new_n17128 ;
  assign new_n17130 = lo0261 & ~new_n15090 ;
  assign new_n17131 = new_n3538 & ~new_n15093 ;
  assign new_n17132 = ~new_n14313 & new_n15093 ;
  assign new_n17133 = ~new_n17131 & ~new_n17132 ;
  assign new_n17134 = new_n15090 & ~new_n17133 ;
  assign new_n17135 = ~new_n17130 & ~new_n17134 ;
  assign new_n17136 = lo0262 & ~new_n14869 ;
  assign new_n17137 = new_n3538 & ~new_n14872 ;
  assign new_n17138 = ~new_n14313 & new_n14872 ;
  assign new_n17139 = ~new_n17137 & ~new_n17138 ;
  assign new_n17140 = new_n14869 & ~new_n17139 ;
  assign new_n17141 = ~new_n17136 & ~new_n17140 ;
  assign new_n17142 = lo0263 & ~new_n14924 ;
  assign new_n17143 = new_n3538 & ~new_n14927 ;
  assign new_n17144 = ~new_n14313 & new_n14927 ;
  assign new_n17145 = ~new_n17143 & ~new_n17144 ;
  assign new_n17146 = new_n14924 & ~new_n17145 ;
  assign new_n17147 = ~new_n17142 & ~new_n17146 ;
  assign new_n17148 = lo0264 & ~new_n15016 ;
  assign new_n17149 = new_n3538 & ~new_n15019 ;
  assign new_n17150 = ~new_n14313 & new_n15019 ;
  assign new_n17151 = ~new_n17149 & ~new_n17150 ;
  assign new_n17152 = new_n15016 & ~new_n17151 ;
  assign new_n17153 = ~new_n17148 & ~new_n17152 ;
  assign new_n17154 = lo0265 & ~new_n15071 ;
  assign new_n17155 = new_n3538 & ~new_n15074 ;
  assign new_n17156 = ~new_n14313 & new_n15074 ;
  assign new_n17157 = ~new_n17155 & ~new_n17156 ;
  assign new_n17158 = new_n15071 & ~new_n17157 ;
  assign new_n17159 = ~new_n17154 & ~new_n17158 ;
  assign new_n17160 = lo0266 & ~new_n14960 ;
  assign new_n17161 = new_n3538 & ~new_n14963 ;
  assign new_n17162 = ~new_n14313 & new_n14963 ;
  assign new_n17163 = ~new_n17161 & ~new_n17162 ;
  assign new_n17164 = new_n14960 & ~new_n17163 ;
  assign new_n17165 = ~new_n17160 & ~new_n17164 ;
  assign new_n17166 = lo0267 & ~new_n14886 ;
  assign new_n17167 = new_n3538 & ~new_n14889 ;
  assign new_n17168 = ~new_n14313 & new_n14889 ;
  assign new_n17169 = ~new_n17167 & ~new_n17168 ;
  assign new_n17170 = new_n14886 & ~new_n17169 ;
  assign new_n17171 = ~new_n17166 & ~new_n17170 ;
  assign new_n17172 = lo0268 & ~new_n15033 ;
  assign new_n17173 = new_n3538 & ~new_n15036 ;
  assign new_n17174 = ~new_n14313 & new_n15036 ;
  assign new_n17175 = ~new_n17173 & ~new_n17174 ;
  assign new_n17176 = new_n15033 & ~new_n17175 ;
  assign new_n17177 = ~new_n17172 & ~new_n17176 ;
  assign new_n17178 = lo0269 & ~new_n15107 ;
  assign new_n17179 = new_n3538 & ~new_n15110 ;
  assign new_n17180 = ~new_n14313 & new_n15110 ;
  assign new_n17181 = ~new_n17179 & ~new_n17180 ;
  assign new_n17182 = new_n15107 & ~new_n17181 ;
  assign new_n17183 = ~new_n17178 & ~new_n17182 ;
  assign new_n17184 = lo0270 & ~new_n14903 ;
  assign new_n17185 = new_n3538 & ~new_n14906 ;
  assign new_n17186 = ~new_n14313 & new_n14906 ;
  assign new_n17187 = ~new_n17185 & ~new_n17186 ;
  assign new_n17188 = new_n14903 & ~new_n17187 ;
  assign new_n17189 = ~new_n17184 & ~new_n17188 ;
  assign new_n17190 = lo0271 & ~new_n14977 ;
  assign new_n17191 = new_n3538 & ~new_n14980 ;
  assign new_n17192 = ~new_n14313 & new_n14980 ;
  assign new_n17193 = ~new_n17191 & ~new_n17192 ;
  assign new_n17194 = new_n14977 & ~new_n17193 ;
  assign new_n17195 = ~new_n17190 & ~new_n17194 ;
  assign new_n17196 = lo0272 & ~new_n15050 ;
  assign new_n17197 = new_n3538 & ~new_n15053 ;
  assign new_n17198 = ~new_n14313 & new_n15053 ;
  assign new_n17199 = ~new_n17197 & ~new_n17198 ;
  assign new_n17200 = new_n15050 & ~new_n17199 ;
  assign new_n17201 = ~new_n17196 & ~new_n17200 ;
  assign new_n17202 = lo0273 & ~new_n15124 ;
  assign new_n17203 = new_n3538 & ~new_n15127 ;
  assign new_n17204 = ~new_n14313 & new_n15127 ;
  assign new_n17205 = ~new_n17203 & ~new_n17204 ;
  assign new_n17206 = new_n15124 & ~new_n17205 ;
  assign new_n17207 = ~new_n17202 & ~new_n17206 ;
  assign new_n17208 = lo0274 & ~new_n15137 ;
  assign new_n17209 = new_n15137 & ~new_n16254 ;
  assign new_n17210 = ~new_n17208 & ~new_n17209 ;
  assign new_n17211 = lo0275 & new_n15454 ;
  assign new_n17212 = lo0958 & ~new_n14313 ;
  assign new_n17213 = ~lo0958 & ~new_n14316 ;
  assign new_n17214 = ~new_n17212 & ~new_n17213 ;
  assign new_n17215 = ~new_n15454 & ~new_n17214 ;
  assign new_n17216 = ~new_n17211 & ~new_n17215 ;
  assign new_n17217 = lo0276 & ~new_n15365 ;
  assign new_n17218 = lo0952 & ~new_n14313 ;
  assign new_n17219 = ~lo0952 & new_n3538 ;
  assign new_n17220 = ~new_n17218 & ~new_n17219 ;
  assign new_n17221 = new_n15365 & ~new_n17220 ;
  assign new_n17222 = ~new_n17217 & ~new_n17221 ;
  assign new_n17223 = lo1066 & ~new_n2252 ;
  assign new_n17224 = lo0277 & ~new_n17223 ;
  assign new_n17225 = ~new_n14313 & new_n17223 ;
  assign new_n17226 = ~new_n17224 & ~new_n17225 ;
  assign new_n17227 = lo0278 & ~new_n14924 ;
  assign new_n17228 = new_n3453 & ~new_n14927 ;
  assign new_n17229 = ~new_n14154 & new_n14927 ;
  assign new_n17230 = ~new_n17228 & ~new_n17229 ;
  assign new_n17231 = new_n14924 & ~new_n17230 ;
  assign new_n17232 = ~new_n17227 & ~new_n17231 ;
  assign new_n17233 = lo0279 & ~new_n14869 ;
  assign new_n17234 = new_n3453 & ~new_n14872 ;
  assign new_n17235 = ~new_n14154 & new_n14872 ;
  assign new_n17236 = ~new_n17234 & ~new_n17235 ;
  assign new_n17237 = new_n14869 & ~new_n17236 ;
  assign new_n17238 = ~new_n17233 & ~new_n17237 ;
  assign new_n17239 = lo0280 & ~new_n15016 ;
  assign new_n17240 = new_n3453 & ~new_n15019 ;
  assign new_n17241 = ~new_n14154 & new_n15019 ;
  assign new_n17242 = ~new_n17240 & ~new_n17241 ;
  assign new_n17243 = new_n15016 & ~new_n17242 ;
  assign new_n17244 = ~new_n17239 & ~new_n17243 ;
  assign new_n17245 = lo0281 & ~new_n15071 ;
  assign new_n17246 = new_n3453 & ~new_n15074 ;
  assign new_n17247 = ~new_n14154 & new_n15074 ;
  assign new_n17248 = ~new_n17246 & ~new_n17247 ;
  assign new_n17249 = new_n15071 & ~new_n17248 ;
  assign new_n17250 = ~new_n17245 & ~new_n17249 ;
  assign new_n17251 = lo0282 & ~new_n14848 ;
  assign new_n17252 = new_n3453 & ~new_n14853 ;
  assign new_n17253 = ~new_n14154 & new_n14853 ;
  assign new_n17254 = ~new_n17252 & ~new_n17253 ;
  assign new_n17255 = new_n14848 & ~new_n17254 ;
  assign new_n17256 = ~new_n17251 & ~new_n17255 ;
  assign new_n17257 = lo0283 & ~new_n14943 ;
  assign new_n17258 = new_n3453 & ~new_n14946 ;
  assign new_n17259 = ~new_n14154 & new_n14946 ;
  assign new_n17260 = ~new_n17258 & ~new_n17259 ;
  assign new_n17261 = new_n14943 & ~new_n17260 ;
  assign new_n17262 = ~new_n17257 & ~new_n17261 ;
  assign new_n17263 = lo0284 & ~new_n14997 ;
  assign new_n17264 = new_n3453 & ~new_n15000 ;
  assign new_n17265 = ~new_n14154 & new_n15000 ;
  assign new_n17266 = ~new_n17264 & ~new_n17265 ;
  assign new_n17267 = new_n14997 & ~new_n17266 ;
  assign new_n17268 = ~new_n17263 & ~new_n17267 ;
  assign new_n17269 = lo0285 & ~new_n15090 ;
  assign new_n17270 = new_n3453 & ~new_n15093 ;
  assign new_n17271 = ~new_n14154 & new_n15093 ;
  assign new_n17272 = ~new_n17270 & ~new_n17271 ;
  assign new_n17273 = new_n15090 & ~new_n17272 ;
  assign new_n17274 = ~new_n17269 & ~new_n17273 ;
  assign new_n17275 = lo0286 & ~new_n14886 ;
  assign new_n17276 = new_n3453 & ~new_n14889 ;
  assign new_n17277 = ~new_n14154 & new_n14889 ;
  assign new_n17278 = ~new_n17276 & ~new_n17277 ;
  assign new_n17279 = new_n14886 & ~new_n17278 ;
  assign new_n17280 = ~new_n17275 & ~new_n17279 ;
  assign new_n17281 = lo0287 & ~new_n14960 ;
  assign new_n17282 = new_n3453 & ~new_n14963 ;
  assign new_n17283 = ~new_n14154 & new_n14963 ;
  assign new_n17284 = ~new_n17282 & ~new_n17283 ;
  assign new_n17285 = new_n14960 & ~new_n17284 ;
  assign new_n17286 = ~new_n17281 & ~new_n17285 ;
  assign new_n17287 = lo0288 & ~new_n15033 ;
  assign new_n17288 = new_n3453 & ~new_n15036 ;
  assign new_n17289 = ~new_n14154 & new_n15036 ;
  assign new_n17290 = ~new_n17288 & ~new_n17289 ;
  assign new_n17291 = new_n15033 & ~new_n17290 ;
  assign new_n17292 = ~new_n17287 & ~new_n17291 ;
  assign new_n17293 = lo0289 & ~new_n15107 ;
  assign new_n17294 = new_n3453 & ~new_n15110 ;
  assign new_n17295 = ~new_n14154 & new_n15110 ;
  assign new_n17296 = ~new_n17294 & ~new_n17295 ;
  assign new_n17297 = new_n15107 & ~new_n17296 ;
  assign new_n17298 = ~new_n17293 & ~new_n17297 ;
  assign new_n17299 = lo0290 & ~new_n14977 ;
  assign new_n17300 = new_n3453 & ~new_n14980 ;
  assign new_n17301 = ~new_n14154 & new_n14980 ;
  assign new_n17302 = ~new_n17300 & ~new_n17301 ;
  assign new_n17303 = new_n14977 & ~new_n17302 ;
  assign new_n17304 = ~new_n17299 & ~new_n17303 ;
  assign new_n17305 = lo0291 & ~new_n14903 ;
  assign new_n17306 = new_n3453 & ~new_n14906 ;
  assign new_n17307 = ~new_n14154 & new_n14906 ;
  assign new_n17308 = ~new_n17306 & ~new_n17307 ;
  assign new_n17309 = new_n14903 & ~new_n17308 ;
  assign new_n17310 = ~new_n17305 & ~new_n17309 ;
  assign new_n17311 = lo0292 & ~new_n15050 ;
  assign new_n17312 = new_n3453 & ~new_n15053 ;
  assign new_n17313 = ~new_n14154 & new_n15053 ;
  assign new_n17314 = ~new_n17312 & ~new_n17313 ;
  assign new_n17315 = new_n15050 & ~new_n17314 ;
  assign new_n17316 = ~new_n17311 & ~new_n17315 ;
  assign new_n17317 = lo0293 & ~new_n15124 ;
  assign new_n17318 = new_n3453 & ~new_n15127 ;
  assign new_n17319 = ~new_n14154 & new_n15127 ;
  assign new_n17320 = ~new_n17318 & ~new_n17319 ;
  assign new_n17321 = new_n15124 & ~new_n17320 ;
  assign new_n17322 = ~new_n17317 & ~new_n17321 ;
  assign new_n17323 = lo0294 & new_n15454 ;
  assign new_n17324 = lo0958 & ~new_n14154 ;
  assign new_n17325 = ~lo0958 & ~new_n14157 ;
  assign new_n17326 = ~new_n17324 & ~new_n17325 ;
  assign new_n17327 = ~new_n15454 & ~new_n17326 ;
  assign new_n17328 = ~new_n17323 & ~new_n17327 ;
  assign new_n17329 = lo0295 & ~new_n15365 ;
  assign new_n17330 = lo0952 & ~new_n14154 ;
  assign new_n17331 = ~lo0952 & new_n3453 ;
  assign new_n17332 = ~new_n17330 & ~new_n17331 ;
  assign new_n17333 = new_n15365 & ~new_n17332 ;
  assign new_n17334 = ~new_n17329 & ~new_n17333 ;
  assign new_n17335 = lo0296 & ~new_n17223 ;
  assign new_n17336 = ~new_n14154 & new_n17223 ;
  assign new_n17337 = ~new_n17335 & ~new_n17336 ;
  assign new_n17338 = lo0297 & ~new_n14699 ;
  assign new_n17339 = new_n13809 & new_n15451 ;
  assign new_n17340 = new_n12441 & new_n17339 ;
  assign new_n17341 = new_n12509 & new_n17340 ;
  assign new_n17342 = new_n14699 & new_n17341 ;
  assign new_n17343 = ~new_n17338 & ~new_n17342 ;
  assign new_n17344 = lo0298 & ~new_n14699 ;
  assign new_n17345 = ~new_n12460 & ~new_n12509 ;
  assign new_n17346 = new_n12460 & new_n12720 ;
  assign new_n17347 = ~new_n17345 & ~new_n17346 ;
  assign new_n17348 = new_n12549 & new_n14699 ;
  assign new_n17349 = new_n17347 & new_n17348 ;
  assign new_n17350 = new_n17339 & new_n17349 ;
  assign new_n17351 = ~new_n17344 & ~new_n17350 ;
  assign new_n17352 = lo0299 & ~new_n14699 ;
  assign new_n17353 = new_n12402 & new_n12508 ;
  assign new_n17354 = ~new_n13809 & ~new_n17353 ;
  assign new_n17355 = new_n12441 & ~new_n17354 ;
  assign new_n17356 = new_n15451 & new_n17355 ;
  assign new_n17357 = new_n2450 & ~new_n12467 ;
  assign new_n17358 = new_n17347 & new_n17357 ;
  assign new_n17359 = ~new_n2450 & new_n12429 ;
  assign new_n17360 = new_n12553 & new_n17359 ;
  assign new_n17361 = ~new_n17358 & ~new_n17360 ;
  assign new_n17362 = new_n14699 & ~new_n17361 ;
  assign new_n17363 = new_n17356 & new_n17362 ;
  assign new_n17364 = ~new_n17352 & ~new_n17363 ;
  assign new_n17365 = lo0300 & ~new_n14699 ;
  assign new_n17366 = ~new_n12460 & new_n14699 ;
  assign new_n17367 = new_n17341 & new_n17366 ;
  assign new_n17368 = ~new_n17365 & ~new_n17367 ;
  assign new_n17369 = lo0301 & ~new_n14848 ;
  assign new_n17370 = new_n4619 & ~new_n14853 ;
  assign new_n17371 = ~new_n14393 & new_n14853 ;
  assign new_n17372 = ~new_n17370 & ~new_n17371 ;
  assign new_n17373 = new_n14848 & ~new_n17372 ;
  assign new_n17374 = ~new_n17369 & ~new_n17373 ;
  assign new_n17375 = lo0302 & ~new_n14869 ;
  assign new_n17376 = new_n4619 & ~new_n14872 ;
  assign new_n17377 = ~new_n14393 & new_n14872 ;
  assign new_n17378 = ~new_n17376 & ~new_n17377 ;
  assign new_n17379 = new_n14869 & ~new_n17378 ;
  assign new_n17380 = ~new_n17375 & ~new_n17379 ;
  assign new_n17381 = lo0303 & ~new_n14886 ;
  assign new_n17382 = new_n4619 & ~new_n14889 ;
  assign new_n17383 = ~new_n14393 & new_n14889 ;
  assign new_n17384 = ~new_n17382 & ~new_n17383 ;
  assign new_n17385 = new_n14886 & ~new_n17384 ;
  assign new_n17386 = ~new_n17381 & ~new_n17385 ;
  assign new_n17387 = lo0304 & ~new_n14903 ;
  assign new_n17388 = new_n4619 & ~new_n14906 ;
  assign new_n17389 = ~new_n14393 & new_n14906 ;
  assign new_n17390 = ~new_n17388 & ~new_n17389 ;
  assign new_n17391 = new_n14903 & ~new_n17390 ;
  assign new_n17392 = ~new_n17387 & ~new_n17391 ;
  assign new_n17393 = lo0305 & ~new_n14924 ;
  assign new_n17394 = new_n4619 & ~new_n14927 ;
  assign new_n17395 = ~new_n14393 & new_n14927 ;
  assign new_n17396 = ~new_n17394 & ~new_n17395 ;
  assign new_n17397 = new_n14924 & ~new_n17396 ;
  assign new_n17398 = ~new_n17393 & ~new_n17397 ;
  assign new_n17399 = lo0306 & ~new_n14943 ;
  assign new_n17400 = new_n4619 & ~new_n14946 ;
  assign new_n17401 = ~new_n14393 & new_n14946 ;
  assign new_n17402 = ~new_n17400 & ~new_n17401 ;
  assign new_n17403 = new_n14943 & ~new_n17402 ;
  assign new_n17404 = ~new_n17399 & ~new_n17403 ;
  assign new_n17405 = lo0307 & ~new_n14960 ;
  assign new_n17406 = new_n4619 & ~new_n14963 ;
  assign new_n17407 = ~new_n14393 & new_n14963 ;
  assign new_n17408 = ~new_n17406 & ~new_n17407 ;
  assign new_n17409 = new_n14960 & ~new_n17408 ;
  assign new_n17410 = ~new_n17405 & ~new_n17409 ;
  assign new_n17411 = lo0308 & ~new_n14977 ;
  assign new_n17412 = new_n4619 & ~new_n14980 ;
  assign new_n17413 = ~new_n14393 & new_n14980 ;
  assign new_n17414 = ~new_n17412 & ~new_n17413 ;
  assign new_n17415 = new_n14977 & ~new_n17414 ;
  assign new_n17416 = ~new_n17411 & ~new_n17415 ;
  assign new_n17417 = lo0309 & ~new_n14997 ;
  assign new_n17418 = new_n4619 & ~new_n15000 ;
  assign new_n17419 = ~new_n14393 & new_n15000 ;
  assign new_n17420 = ~new_n17418 & ~new_n17419 ;
  assign new_n17421 = new_n14997 & ~new_n17420 ;
  assign new_n17422 = ~new_n17417 & ~new_n17421 ;
  assign new_n17423 = lo0310 & ~new_n15016 ;
  assign new_n17424 = new_n4619 & ~new_n15019 ;
  assign new_n17425 = ~new_n14393 & new_n15019 ;
  assign new_n17426 = ~new_n17424 & ~new_n17425 ;
  assign new_n17427 = new_n15016 & ~new_n17426 ;
  assign new_n17428 = ~new_n17423 & ~new_n17427 ;
  assign new_n17429 = lo0311 & ~new_n15033 ;
  assign new_n17430 = new_n4619 & ~new_n15036 ;
  assign new_n17431 = ~new_n14393 & new_n15036 ;
  assign new_n17432 = ~new_n17430 & ~new_n17431 ;
  assign new_n17433 = new_n15033 & ~new_n17432 ;
  assign new_n17434 = ~new_n17429 & ~new_n17433 ;
  assign new_n17435 = lo0312 & ~new_n15050 ;
  assign new_n17436 = new_n4619 & ~new_n15053 ;
  assign new_n17437 = ~new_n14393 & new_n15053 ;
  assign new_n17438 = ~new_n17436 & ~new_n17437 ;
  assign new_n17439 = new_n15050 & ~new_n17438 ;
  assign new_n17440 = ~new_n17435 & ~new_n17439 ;
  assign new_n17441 = lo0313 & ~new_n15071 ;
  assign new_n17442 = new_n4619 & ~new_n15074 ;
  assign new_n17443 = ~new_n14393 & new_n15074 ;
  assign new_n17444 = ~new_n17442 & ~new_n17443 ;
  assign new_n17445 = new_n15071 & ~new_n17444 ;
  assign new_n17446 = ~new_n17441 & ~new_n17445 ;
  assign new_n17447 = lo0314 & ~new_n15090 ;
  assign new_n17448 = new_n4619 & ~new_n15093 ;
  assign new_n17449 = ~new_n14393 & new_n15093 ;
  assign new_n17450 = ~new_n17448 & ~new_n17449 ;
  assign new_n17451 = new_n15090 & ~new_n17450 ;
  assign new_n17452 = ~new_n17447 & ~new_n17451 ;
  assign new_n17453 = lo0315 & ~new_n15107 ;
  assign new_n17454 = new_n4619 & ~new_n15110 ;
  assign new_n17455 = ~new_n14393 & new_n15110 ;
  assign new_n17456 = ~new_n17454 & ~new_n17455 ;
  assign new_n17457 = new_n15107 & ~new_n17456 ;
  assign new_n17458 = ~new_n17453 & ~new_n17457 ;
  assign new_n17459 = lo0316 & ~new_n15124 ;
  assign new_n17460 = new_n4619 & ~new_n15127 ;
  assign new_n17461 = ~new_n14393 & new_n15127 ;
  assign new_n17462 = ~new_n17460 & ~new_n17461 ;
  assign new_n17463 = new_n15124 & ~new_n17462 ;
  assign new_n17464 = ~new_n17459 & ~new_n17463 ;
  assign new_n17465 = lo0317 & ~new_n15137 ;
  assign new_n17466 = new_n15137 & ~new_n15723 ;
  assign new_n17467 = ~new_n17465 & ~new_n17466 ;
  assign new_n17468 = lo0318 & new_n15454 ;
  assign new_n17469 = lo0958 & ~new_n14393 ;
  assign new_n17470 = ~lo0958 & ~new_n14397 ;
  assign new_n17471 = ~new_n17469 & ~new_n17470 ;
  assign new_n17472 = ~new_n15454 & ~new_n17471 ;
  assign new_n17473 = ~new_n17468 & ~new_n17472 ;
  assign new_n17474 = lo0319 & ~new_n15365 ;
  assign new_n17475 = lo0952 & ~new_n14393 ;
  assign new_n17476 = ~lo0952 & new_n4619 ;
  assign new_n17477 = ~new_n17475 & ~new_n17476 ;
  assign new_n17478 = new_n15365 & ~new_n17477 ;
  assign new_n17479 = ~new_n17474 & ~new_n17478 ;
  assign new_n17480 = lo0320 & ~new_n17223 ;
  assign new_n17481 = ~new_n14393 & new_n17223 ;
  assign new_n17482 = ~new_n17480 & ~new_n17481 ;
  assign new_n17483 = lo0321 & ~new_n17223 ;
  assign new_n17484 = ~new_n16735 & new_n17223 ;
  assign new_n17485 = ~new_n17483 & ~new_n17484 ;
  assign new_n17486 = lo0322 & ~new_n14943 ;
  assign new_n17487 = new_n4981 & ~new_n14946 ;
  assign new_n17488 = ~new_n14419 & new_n14946 ;
  assign new_n17489 = ~new_n17487 & ~new_n17488 ;
  assign new_n17490 = new_n14943 & ~new_n17489 ;
  assign new_n17491 = ~new_n17486 & ~new_n17490 ;
  assign new_n17492 = lo0323 & ~new_n14848 ;
  assign new_n17493 = new_n4981 & ~new_n14853 ;
  assign new_n17494 = ~new_n14419 & new_n14853 ;
  assign new_n17495 = ~new_n17493 & ~new_n17494 ;
  assign new_n17496 = new_n14848 & ~new_n17495 ;
  assign new_n17497 = ~new_n17492 & ~new_n17496 ;
  assign new_n17498 = lo0324 & ~new_n14997 ;
  assign new_n17499 = new_n4981 & ~new_n15000 ;
  assign new_n17500 = ~new_n14419 & new_n15000 ;
  assign new_n17501 = ~new_n17499 & ~new_n17500 ;
  assign new_n17502 = new_n14997 & ~new_n17501 ;
  assign new_n17503 = ~new_n17498 & ~new_n17502 ;
  assign new_n17504 = lo0325 & ~new_n15090 ;
  assign new_n17505 = new_n4981 & ~new_n15093 ;
  assign new_n17506 = ~new_n14419 & new_n15093 ;
  assign new_n17507 = ~new_n17505 & ~new_n17506 ;
  assign new_n17508 = new_n15090 & ~new_n17507 ;
  assign new_n17509 = ~new_n17504 & ~new_n17508 ;
  assign new_n17510 = lo0326 & ~new_n14869 ;
  assign new_n17511 = new_n4981 & ~new_n14872 ;
  assign new_n17512 = ~new_n14419 & new_n14872 ;
  assign new_n17513 = ~new_n17511 & ~new_n17512 ;
  assign new_n17514 = new_n14869 & ~new_n17513 ;
  assign new_n17515 = ~new_n17510 & ~new_n17514 ;
  assign new_n17516 = lo0327 & ~new_n14924 ;
  assign new_n17517 = new_n4981 & ~new_n14927 ;
  assign new_n17518 = ~new_n14419 & new_n14927 ;
  assign new_n17519 = ~new_n17517 & ~new_n17518 ;
  assign new_n17520 = new_n14924 & ~new_n17519 ;
  assign new_n17521 = ~new_n17516 & ~new_n17520 ;
  assign new_n17522 = lo0328 & ~new_n15016 ;
  assign new_n17523 = new_n4981 & ~new_n15019 ;
  assign new_n17524 = ~new_n14419 & new_n15019 ;
  assign new_n17525 = ~new_n17523 & ~new_n17524 ;
  assign new_n17526 = new_n15016 & ~new_n17525 ;
  assign new_n17527 = ~new_n17522 & ~new_n17526 ;
  assign new_n17528 = lo0329 & ~new_n15071 ;
  assign new_n17529 = new_n4981 & ~new_n15074 ;
  assign new_n17530 = ~new_n14419 & new_n15074 ;
  assign new_n17531 = ~new_n17529 & ~new_n17530 ;
  assign new_n17532 = new_n15071 & ~new_n17531 ;
  assign new_n17533 = ~new_n17528 & ~new_n17532 ;
  assign new_n17534 = lo0330 & ~new_n14960 ;
  assign new_n17535 = new_n4981 & ~new_n14963 ;
  assign new_n17536 = ~new_n14419 & new_n14963 ;
  assign new_n17537 = ~new_n17535 & ~new_n17536 ;
  assign new_n17538 = new_n14960 & ~new_n17537 ;
  assign new_n17539 = ~new_n17534 & ~new_n17538 ;
  assign new_n17540 = lo0331 & ~new_n14886 ;
  assign new_n17541 = new_n4981 & ~new_n14889 ;
  assign new_n17542 = ~new_n14419 & new_n14889 ;
  assign new_n17543 = ~new_n17541 & ~new_n17542 ;
  assign new_n17544 = new_n14886 & ~new_n17543 ;
  assign new_n17545 = ~new_n17540 & ~new_n17544 ;
  assign new_n17546 = lo0332 & ~new_n15033 ;
  assign new_n17547 = new_n4981 & ~new_n15036 ;
  assign new_n17548 = ~new_n14419 & new_n15036 ;
  assign new_n17549 = ~new_n17547 & ~new_n17548 ;
  assign new_n17550 = new_n15033 & ~new_n17549 ;
  assign new_n17551 = ~new_n17546 & ~new_n17550 ;
  assign new_n17552 = lo0333 & ~new_n15107 ;
  assign new_n17553 = new_n4981 & ~new_n15110 ;
  assign new_n17554 = ~new_n14419 & new_n15110 ;
  assign new_n17555 = ~new_n17553 & ~new_n17554 ;
  assign new_n17556 = new_n15107 & ~new_n17555 ;
  assign new_n17557 = ~new_n17552 & ~new_n17556 ;
  assign new_n17558 = lo0334 & ~new_n14903 ;
  assign new_n17559 = new_n4981 & ~new_n14906 ;
  assign new_n17560 = ~new_n14419 & new_n14906 ;
  assign new_n17561 = ~new_n17559 & ~new_n17560 ;
  assign new_n17562 = new_n14903 & ~new_n17561 ;
  assign new_n17563 = ~new_n17558 & ~new_n17562 ;
  assign new_n17564 = lo0335 & ~new_n14977 ;
  assign new_n17565 = new_n4981 & ~new_n14980 ;
  assign new_n17566 = ~new_n14419 & new_n14980 ;
  assign new_n17567 = ~new_n17565 & ~new_n17566 ;
  assign new_n17568 = new_n14977 & ~new_n17567 ;
  assign new_n17569 = ~new_n17564 & ~new_n17568 ;
  assign new_n17570 = lo0336 & ~new_n15050 ;
  assign new_n17571 = new_n4981 & ~new_n15053 ;
  assign new_n17572 = ~new_n14419 & new_n15053 ;
  assign new_n17573 = ~new_n17571 & ~new_n17572 ;
  assign new_n17574 = new_n15050 & ~new_n17573 ;
  assign new_n17575 = ~new_n17570 & ~new_n17574 ;
  assign new_n17576 = lo0337 & ~new_n15124 ;
  assign new_n17577 = new_n4981 & ~new_n15127 ;
  assign new_n17578 = ~new_n14419 & new_n15127 ;
  assign new_n17579 = ~new_n17577 & ~new_n17578 ;
  assign new_n17580 = new_n15124 & ~new_n17579 ;
  assign new_n17581 = ~new_n17576 & ~new_n17580 ;
  assign new_n17582 = lo0338 & ~new_n15137 ;
  assign new_n17583 = new_n15137 & ~new_n16079 ;
  assign new_n17584 = ~new_n17582 & ~new_n17583 ;
  assign new_n17585 = lo0339 & new_n15454 ;
  assign new_n17586 = lo0958 & ~new_n14419 ;
  assign new_n17587 = ~lo0958 & ~new_n14422 ;
  assign new_n17588 = ~new_n17586 & ~new_n17587 ;
  assign new_n17589 = ~new_n15454 & ~new_n17588 ;
  assign new_n17590 = ~new_n17585 & ~new_n17589 ;
  assign new_n17591 = lo0340 & ~new_n15365 ;
  assign new_n17592 = lo0952 & ~new_n14419 ;
  assign new_n17593 = ~lo0952 & new_n4981 ;
  assign new_n17594 = ~new_n17592 & ~new_n17593 ;
  assign new_n17595 = new_n15365 & ~new_n17594 ;
  assign new_n17596 = ~new_n17591 & ~new_n17595 ;
  assign new_n17597 = lo0341 & ~new_n17223 ;
  assign new_n17598 = ~new_n14419 & new_n17223 ;
  assign new_n17599 = ~new_n17597 & ~new_n17598 ;
  assign new_n17600 = lo0342 & ~new_n14848 ;
  assign new_n17601 = ~new_n4168 & ~new_n14853 ;
  assign new_n17602 = ~new_n14552 & new_n14853 ;
  assign new_n17603 = ~new_n17601 & ~new_n17602 ;
  assign new_n17604 = new_n14848 & ~new_n17603 ;
  assign new_n17605 = ~new_n17600 & ~new_n17604 ;
  assign new_n17606 = lo0343 & ~new_n14869 ;
  assign new_n17607 = ~new_n4168 & ~new_n14872 ;
  assign new_n17608 = ~new_n14552 & new_n14872 ;
  assign new_n17609 = ~new_n17607 & ~new_n17608 ;
  assign new_n17610 = new_n14869 & ~new_n17609 ;
  assign new_n17611 = ~new_n17606 & ~new_n17610 ;
  assign new_n17612 = lo0344 & ~new_n14886 ;
  assign new_n17613 = ~new_n4168 & ~new_n14889 ;
  assign new_n17614 = ~new_n14552 & new_n14889 ;
  assign new_n17615 = ~new_n17613 & ~new_n17614 ;
  assign new_n17616 = new_n14886 & ~new_n17615 ;
  assign new_n17617 = ~new_n17612 & ~new_n17616 ;
  assign new_n17618 = lo0345 & ~new_n14903 ;
  assign new_n17619 = ~new_n4168 & ~new_n14906 ;
  assign new_n17620 = ~new_n14552 & new_n14906 ;
  assign new_n17621 = ~new_n17619 & ~new_n17620 ;
  assign new_n17622 = new_n14903 & ~new_n17621 ;
  assign new_n17623 = ~new_n17618 & ~new_n17622 ;
  assign new_n17624 = lo0346 & ~new_n14924 ;
  assign new_n17625 = ~new_n4168 & ~new_n14927 ;
  assign new_n17626 = ~new_n14552 & new_n14927 ;
  assign new_n17627 = ~new_n17625 & ~new_n17626 ;
  assign new_n17628 = new_n14924 & ~new_n17627 ;
  assign new_n17629 = ~new_n17624 & ~new_n17628 ;
  assign new_n17630 = lo0347 & ~new_n14943 ;
  assign new_n17631 = ~new_n4168 & ~new_n14946 ;
  assign new_n17632 = ~new_n14552 & new_n14946 ;
  assign new_n17633 = ~new_n17631 & ~new_n17632 ;
  assign new_n17634 = new_n14943 & ~new_n17633 ;
  assign new_n17635 = ~new_n17630 & ~new_n17634 ;
  assign new_n17636 = lo0348 & ~new_n14960 ;
  assign new_n17637 = ~new_n4168 & ~new_n14963 ;
  assign new_n17638 = ~new_n14552 & new_n14963 ;
  assign new_n17639 = ~new_n17637 & ~new_n17638 ;
  assign new_n17640 = new_n14960 & ~new_n17639 ;
  assign new_n17641 = ~new_n17636 & ~new_n17640 ;
  assign new_n17642 = lo0349 & ~new_n14977 ;
  assign new_n17643 = ~new_n4168 & ~new_n14980 ;
  assign new_n17644 = ~new_n14552 & new_n14980 ;
  assign new_n17645 = ~new_n17643 & ~new_n17644 ;
  assign new_n17646 = new_n14977 & ~new_n17645 ;
  assign new_n17647 = ~new_n17642 & ~new_n17646 ;
  assign new_n17648 = lo0350 & ~new_n14997 ;
  assign new_n17649 = ~new_n4168 & ~new_n15000 ;
  assign new_n17650 = ~new_n14552 & new_n15000 ;
  assign new_n17651 = ~new_n17649 & ~new_n17650 ;
  assign new_n17652 = new_n14997 & ~new_n17651 ;
  assign new_n17653 = ~new_n17648 & ~new_n17652 ;
  assign new_n17654 = lo0351 & ~new_n15016 ;
  assign new_n17655 = ~new_n4168 & ~new_n15019 ;
  assign new_n17656 = ~new_n14552 & new_n15019 ;
  assign new_n17657 = ~new_n17655 & ~new_n17656 ;
  assign new_n17658 = new_n15016 & ~new_n17657 ;
  assign new_n17659 = ~new_n17654 & ~new_n17658 ;
  assign new_n17660 = lo0352 & ~new_n15050 ;
  assign new_n17661 = ~new_n4168 & ~new_n15053 ;
  assign new_n17662 = ~new_n14552 & new_n15053 ;
  assign new_n17663 = ~new_n17661 & ~new_n17662 ;
  assign new_n17664 = new_n15050 & ~new_n17663 ;
  assign new_n17665 = ~new_n17660 & ~new_n17664 ;
  assign new_n17666 = lo0353 & ~new_n15071 ;
  assign new_n17667 = ~new_n4168 & ~new_n15074 ;
  assign new_n17668 = ~new_n14552 & new_n15074 ;
  assign new_n17669 = ~new_n17667 & ~new_n17668 ;
  assign new_n17670 = new_n15071 & ~new_n17669 ;
  assign new_n17671 = ~new_n17666 & ~new_n17670 ;
  assign new_n17672 = lo0354 & ~new_n15090 ;
  assign new_n17673 = ~new_n4168 & ~new_n15093 ;
  assign new_n17674 = ~new_n14552 & new_n15093 ;
  assign new_n17675 = ~new_n17673 & ~new_n17674 ;
  assign new_n17676 = new_n15090 & ~new_n17675 ;
  assign new_n17677 = ~new_n17672 & ~new_n17676 ;
  assign new_n17678 = lo0355 & ~new_n15107 ;
  assign new_n17679 = ~new_n4168 & ~new_n15110 ;
  assign new_n17680 = ~new_n14552 & new_n15110 ;
  assign new_n17681 = ~new_n17679 & ~new_n17680 ;
  assign new_n17682 = new_n15107 & ~new_n17681 ;
  assign new_n17683 = ~new_n17678 & ~new_n17682 ;
  assign new_n17684 = lo0356 & ~new_n15124 ;
  assign new_n17685 = ~new_n4168 & ~new_n15127 ;
  assign new_n17686 = ~new_n14552 & new_n15127 ;
  assign new_n17687 = ~new_n17685 & ~new_n17686 ;
  assign new_n17688 = new_n15124 & ~new_n17687 ;
  assign new_n17689 = ~new_n17684 & ~new_n17688 ;
  assign new_n17690 = lo0357 & new_n15454 ;
  assign new_n17691 = lo0958 & ~new_n14552 ;
  assign new_n17692 = ~lo0958 & ~new_n14556 ;
  assign new_n17693 = ~new_n17691 & ~new_n17692 ;
  assign new_n17694 = ~new_n15454 & ~new_n17693 ;
  assign new_n17695 = ~new_n17690 & ~new_n17694 ;
  assign new_n17696 = lo0358 & ~new_n15365 ;
  assign new_n17697 = lo0952 & ~new_n14552 ;
  assign new_n17698 = ~lo0952 & ~new_n4168 ;
  assign new_n17699 = ~new_n17697 & ~new_n17698 ;
  assign new_n17700 = new_n15365 & ~new_n17699 ;
  assign new_n17701 = ~new_n17696 & ~new_n17700 ;
  assign new_n17702 = lo0359 & ~new_n17223 ;
  assign new_n17703 = ~new_n14552 & new_n17223 ;
  assign new_n17704 = ~new_n17702 & ~new_n17703 ;
  assign new_n17705 = ~lo0955 & ~lo0956 ;
  assign new_n17706 = ~new_n2252 & ~new_n17705 ;
  assign new_n17707 = lo0360 & ~new_n17706 ;
  assign new_n17708 = lo0955 & ~new_n14552 ;
  assign new_n17709 = ~lo0955 & ~new_n4168 ;
  assign new_n17710 = ~new_n17708 & ~new_n17709 ;
  assign new_n17711 = new_n17706 & ~new_n17710 ;
  assign new_n17712 = ~new_n17707 & ~new_n17711 ;
  assign new_n17713 = lo0361 & ~new_n14943 ;
  assign new_n17714 = new_n3897 & ~new_n14946 ;
  assign new_n17715 = ~new_n14340 & new_n14946 ;
  assign new_n17716 = ~new_n17714 & ~new_n17715 ;
  assign new_n17717 = new_n14943 & ~new_n17716 ;
  assign new_n17718 = ~new_n17713 & ~new_n17717 ;
  assign new_n17719 = lo0362 & ~new_n14924 ;
  assign new_n17720 = new_n3897 & ~new_n14927 ;
  assign new_n17721 = ~new_n14340 & new_n14927 ;
  assign new_n17722 = ~new_n17720 & ~new_n17721 ;
  assign new_n17723 = new_n14924 & ~new_n17722 ;
  assign new_n17724 = ~new_n17719 & ~new_n17723 ;
  assign new_n17725 = lo0363 & ~new_n14960 ;
  assign new_n17726 = new_n3897 & ~new_n14963 ;
  assign new_n17727 = ~new_n14340 & new_n14963 ;
  assign new_n17728 = ~new_n17726 & ~new_n17727 ;
  assign new_n17729 = new_n14960 & ~new_n17728 ;
  assign new_n17730 = ~new_n17725 & ~new_n17729 ;
  assign new_n17731 = lo0364 & ~new_n14977 ;
  assign new_n17732 = new_n3897 & ~new_n14980 ;
  assign new_n17733 = ~new_n14340 & new_n14980 ;
  assign new_n17734 = ~new_n17732 & ~new_n17733 ;
  assign new_n17735 = new_n14977 & ~new_n17734 ;
  assign new_n17736 = ~new_n17731 & ~new_n17735 ;
  assign new_n17737 = lo0365 & ~new_n14869 ;
  assign new_n17738 = new_n3897 & ~new_n14872 ;
  assign new_n17739 = ~new_n14340 & new_n14872 ;
  assign new_n17740 = ~new_n17738 & ~new_n17739 ;
  assign new_n17741 = new_n14869 & ~new_n17740 ;
  assign new_n17742 = ~new_n17737 & ~new_n17741 ;
  assign new_n17743 = lo0366 & ~new_n14848 ;
  assign new_n17744 = new_n3897 & ~new_n14853 ;
  assign new_n17745 = ~new_n14340 & new_n14853 ;
  assign new_n17746 = ~new_n17744 & ~new_n17745 ;
  assign new_n17747 = new_n14848 & ~new_n17746 ;
  assign new_n17748 = ~new_n17743 & ~new_n17747 ;
  assign new_n17749 = lo0367 & ~new_n14886 ;
  assign new_n17750 = new_n3897 & ~new_n14889 ;
  assign new_n17751 = ~new_n14340 & new_n14889 ;
  assign new_n17752 = ~new_n17750 & ~new_n17751 ;
  assign new_n17753 = new_n14886 & ~new_n17752 ;
  assign new_n17754 = ~new_n17749 & ~new_n17753 ;
  assign new_n17755 = lo0368 & ~new_n14903 ;
  assign new_n17756 = new_n3897 & ~new_n14906 ;
  assign new_n17757 = ~new_n14340 & new_n14906 ;
  assign new_n17758 = ~new_n17756 & ~new_n17757 ;
  assign new_n17759 = new_n14903 & ~new_n17758 ;
  assign new_n17760 = ~new_n17755 & ~new_n17759 ;
  assign new_n17761 = lo0369 & ~new_n15016 ;
  assign new_n17762 = new_n3897 & ~new_n15019 ;
  assign new_n17763 = ~new_n14340 & new_n15019 ;
  assign new_n17764 = ~new_n17762 & ~new_n17763 ;
  assign new_n17765 = new_n15016 & ~new_n17764 ;
  assign new_n17766 = ~new_n17761 & ~new_n17765 ;
  assign new_n17767 = lo0370 & ~new_n14997 ;
  assign new_n17768 = new_n3897 & ~new_n15000 ;
  assign new_n17769 = ~new_n14340 & new_n15000 ;
  assign new_n17770 = ~new_n17768 & ~new_n17769 ;
  assign new_n17771 = new_n14997 & ~new_n17770 ;
  assign new_n17772 = ~new_n17767 & ~new_n17771 ;
  assign new_n17773 = lo0371 & ~new_n15033 ;
  assign new_n17774 = new_n3897 & ~new_n15036 ;
  assign new_n17775 = ~new_n14340 & new_n15036 ;
  assign new_n17776 = ~new_n17774 & ~new_n17775 ;
  assign new_n17777 = new_n15033 & ~new_n17776 ;
  assign new_n17778 = ~new_n17773 & ~new_n17777 ;
  assign new_n17779 = lo0372 & ~new_n15050 ;
  assign new_n17780 = new_n3897 & ~new_n15053 ;
  assign new_n17781 = ~new_n14340 & new_n15053 ;
  assign new_n17782 = ~new_n17780 & ~new_n17781 ;
  assign new_n17783 = new_n15050 & ~new_n17782 ;
  assign new_n17784 = ~new_n17779 & ~new_n17783 ;
  assign new_n17785 = lo0373 & ~new_n15090 ;
  assign new_n17786 = new_n3897 & ~new_n15093 ;
  assign new_n17787 = ~new_n14340 & new_n15093 ;
  assign new_n17788 = ~new_n17786 & ~new_n17787 ;
  assign new_n17789 = new_n15090 & ~new_n17788 ;
  assign new_n17790 = ~new_n17785 & ~new_n17789 ;
  assign new_n17791 = lo0374 & ~new_n15071 ;
  assign new_n17792 = new_n3897 & ~new_n15074 ;
  assign new_n17793 = ~new_n14340 & new_n15074 ;
  assign new_n17794 = ~new_n17792 & ~new_n17793 ;
  assign new_n17795 = new_n15071 & ~new_n17794 ;
  assign new_n17796 = ~new_n17791 & ~new_n17795 ;
  assign new_n17797 = lo0375 & ~new_n15107 ;
  assign new_n17798 = new_n3897 & ~new_n15110 ;
  assign new_n17799 = ~new_n14340 & new_n15110 ;
  assign new_n17800 = ~new_n17798 & ~new_n17799 ;
  assign new_n17801 = new_n15107 & ~new_n17800 ;
  assign new_n17802 = ~new_n17797 & ~new_n17801 ;
  assign new_n17803 = lo0376 & ~new_n15124 ;
  assign new_n17804 = new_n3897 & ~new_n15127 ;
  assign new_n17805 = ~new_n14340 & new_n15127 ;
  assign new_n17806 = ~new_n17804 & ~new_n17805 ;
  assign new_n17807 = new_n15124 & ~new_n17806 ;
  assign new_n17808 = ~new_n17803 & ~new_n17807 ;
  assign new_n17809 = lo0377 & ~new_n15137 ;
  assign new_n17810 = new_n15137 & ~new_n15998 ;
  assign new_n17811 = ~new_n17809 & ~new_n17810 ;
  assign new_n17812 = lo0378 & new_n15454 ;
  assign new_n17813 = lo0958 & ~new_n14340 ;
  assign new_n17814 = ~lo0958 & ~new_n14344 ;
  assign new_n17815 = ~new_n17813 & ~new_n17814 ;
  assign new_n17816 = ~new_n15454 & ~new_n17815 ;
  assign new_n17817 = ~new_n17812 & ~new_n17816 ;
  assign new_n17818 = lo0379 & ~new_n15365 ;
  assign new_n17819 = lo0952 & ~new_n14340 ;
  assign new_n17820 = ~lo0952 & new_n3897 ;
  assign new_n17821 = ~new_n17819 & ~new_n17820 ;
  assign new_n17822 = new_n15365 & ~new_n17821 ;
  assign new_n17823 = ~new_n17818 & ~new_n17822 ;
  assign new_n17824 = lo0380 & ~new_n17223 ;
  assign new_n17825 = ~new_n14340 & new_n17223 ;
  assign new_n17826 = ~new_n17824 & ~new_n17825 ;
  assign new_n17827 = lo0381 & ~new_n17223 ;
  assign new_n17828 = ~new_n14366 & new_n17223 ;
  assign new_n17829 = ~new_n17827 & ~new_n17828 ;
  assign new_n17830 = lo0382 & ~new_n14943 ;
  assign new_n17831 = ~new_n5743 & ~new_n14946 ;
  assign new_n17832 = new_n14946 & ~new_n16677 ;
  assign new_n17833 = ~new_n17831 & ~new_n17832 ;
  assign new_n17834 = new_n14943 & ~new_n17833 ;
  assign new_n17835 = ~new_n17830 & ~new_n17834 ;
  assign new_n17836 = lo0383 & ~new_n14848 ;
  assign new_n17837 = ~new_n5743 & ~new_n14853 ;
  assign new_n17838 = new_n14853 & ~new_n16677 ;
  assign new_n17839 = ~new_n17837 & ~new_n17838 ;
  assign new_n17840 = new_n14848 & ~new_n17839 ;
  assign new_n17841 = ~new_n17836 & ~new_n17840 ;
  assign new_n17842 = lo0384 & ~new_n14997 ;
  assign new_n17843 = ~new_n5743 & ~new_n15000 ;
  assign new_n17844 = new_n15000 & ~new_n16677 ;
  assign new_n17845 = ~new_n17843 & ~new_n17844 ;
  assign new_n17846 = new_n14997 & ~new_n17845 ;
  assign new_n17847 = ~new_n17842 & ~new_n17846 ;
  assign new_n17848 = lo0385 & ~new_n15090 ;
  assign new_n17849 = ~new_n5743 & ~new_n15093 ;
  assign new_n17850 = new_n15093 & ~new_n16677 ;
  assign new_n17851 = ~new_n17849 & ~new_n17850 ;
  assign new_n17852 = new_n15090 & ~new_n17851 ;
  assign new_n17853 = ~new_n17848 & ~new_n17852 ;
  assign new_n17854 = lo0386 & ~new_n14869 ;
  assign new_n17855 = ~new_n5743 & ~new_n14872 ;
  assign new_n17856 = new_n14872 & ~new_n16677 ;
  assign new_n17857 = ~new_n17855 & ~new_n17856 ;
  assign new_n17858 = new_n14869 & ~new_n17857 ;
  assign new_n17859 = ~new_n17854 & ~new_n17858 ;
  assign new_n17860 = lo0387 & ~new_n14924 ;
  assign new_n17861 = ~new_n5743 & ~new_n14927 ;
  assign new_n17862 = new_n14927 & ~new_n16677 ;
  assign new_n17863 = ~new_n17861 & ~new_n17862 ;
  assign new_n17864 = new_n14924 & ~new_n17863 ;
  assign new_n17865 = ~new_n17860 & ~new_n17864 ;
  assign new_n17866 = lo0388 & ~new_n15016 ;
  assign new_n17867 = ~new_n5743 & ~new_n15019 ;
  assign new_n17868 = new_n15019 & ~new_n16677 ;
  assign new_n17869 = ~new_n17867 & ~new_n17868 ;
  assign new_n17870 = new_n15016 & ~new_n17869 ;
  assign new_n17871 = ~new_n17866 & ~new_n17870 ;
  assign new_n17872 = lo0389 & ~new_n15071 ;
  assign new_n17873 = ~new_n5743 & ~new_n15074 ;
  assign new_n17874 = new_n15074 & ~new_n16677 ;
  assign new_n17875 = ~new_n17873 & ~new_n17874 ;
  assign new_n17876 = new_n15071 & ~new_n17875 ;
  assign new_n17877 = ~new_n17872 & ~new_n17876 ;
  assign new_n17878 = lo0390 & ~new_n14960 ;
  assign new_n17879 = ~new_n5743 & ~new_n14963 ;
  assign new_n17880 = new_n14963 & ~new_n16677 ;
  assign new_n17881 = ~new_n17879 & ~new_n17880 ;
  assign new_n17882 = new_n14960 & ~new_n17881 ;
  assign new_n17883 = ~new_n17878 & ~new_n17882 ;
  assign new_n17884 = lo0391 & ~new_n14886 ;
  assign new_n17885 = ~new_n5743 & ~new_n14889 ;
  assign new_n17886 = new_n14889 & ~new_n16677 ;
  assign new_n17887 = ~new_n17885 & ~new_n17886 ;
  assign new_n17888 = new_n14886 & ~new_n17887 ;
  assign new_n17889 = ~new_n17884 & ~new_n17888 ;
  assign new_n17890 = lo0392 & ~new_n15033 ;
  assign new_n17891 = ~new_n5743 & ~new_n15036 ;
  assign new_n17892 = new_n15036 & ~new_n16677 ;
  assign new_n17893 = ~new_n17891 & ~new_n17892 ;
  assign new_n17894 = new_n15033 & ~new_n17893 ;
  assign new_n17895 = ~new_n17890 & ~new_n17894 ;
  assign new_n17896 = lo0393 & ~new_n15107 ;
  assign new_n17897 = ~new_n5743 & ~new_n15110 ;
  assign new_n17898 = new_n15110 & ~new_n16677 ;
  assign new_n17899 = ~new_n17897 & ~new_n17898 ;
  assign new_n17900 = new_n15107 & ~new_n17899 ;
  assign new_n17901 = ~new_n17896 & ~new_n17900 ;
  assign new_n17902 = lo0394 & ~new_n14903 ;
  assign new_n17903 = ~new_n5743 & ~new_n14906 ;
  assign new_n17904 = new_n14906 & ~new_n16677 ;
  assign new_n17905 = ~new_n17903 & ~new_n17904 ;
  assign new_n17906 = new_n14903 & ~new_n17905 ;
  assign new_n17907 = ~new_n17902 & ~new_n17906 ;
  assign new_n17908 = lo0395 & ~new_n14977 ;
  assign new_n17909 = ~new_n5743 & ~new_n14980 ;
  assign new_n17910 = new_n14980 & ~new_n16677 ;
  assign new_n17911 = ~new_n17909 & ~new_n17910 ;
  assign new_n17912 = new_n14977 & ~new_n17911 ;
  assign new_n17913 = ~new_n17908 & ~new_n17912 ;
  assign new_n17914 = lo0396 & ~new_n15050 ;
  assign new_n17915 = ~new_n5743 & ~new_n15053 ;
  assign new_n17916 = new_n15053 & ~new_n16677 ;
  assign new_n17917 = ~new_n17915 & ~new_n17916 ;
  assign new_n17918 = new_n15050 & ~new_n17917 ;
  assign new_n17919 = ~new_n17914 & ~new_n17918 ;
  assign new_n17920 = lo0397 & ~new_n15124 ;
  assign new_n17921 = ~new_n5743 & ~new_n15127 ;
  assign new_n17922 = new_n15127 & ~new_n16677 ;
  assign new_n17923 = ~new_n17921 & ~new_n17922 ;
  assign new_n17924 = new_n15124 & ~new_n17923 ;
  assign new_n17925 = ~new_n17920 & ~new_n17924 ;
  assign new_n17926 = lo0398 & new_n2252 ;
  assign new_n17927 = ~new_n2252 & ~new_n12467 ;
  assign new_n17928 = ~new_n17926 & ~new_n17927 ;
  assign new_n17929 = lo0399 & new_n15454 ;
  assign new_n17930 = lo0958 & ~new_n16677 ;
  assign new_n17931 = lo0399 & ~new_n13948 ;
  assign new_n17932 = ~lo0399 & new_n13948 ;
  assign new_n17933 = ~new_n17931 & ~new_n17932 ;
  assign new_n17934 = ~lo0958 & ~new_n17933 ;
  assign new_n17935 = ~new_n17930 & ~new_n17934 ;
  assign new_n17936 = ~new_n15454 & ~new_n17935 ;
  assign new_n17937 = ~new_n17929 & ~new_n17936 ;
  assign new_n17938 = lo0400 & ~new_n15365 ;
  assign new_n17939 = lo0952 & ~new_n16677 ;
  assign new_n17940 = ~lo0952 & ~new_n5743 ;
  assign new_n17941 = ~new_n17939 & ~new_n17940 ;
  assign new_n17942 = new_n15365 & ~new_n17941 ;
  assign new_n17943 = ~new_n17938 & ~new_n17942 ;
  assign new_n17944 = lo0401 & ~new_n15033 ;
  assign new_n17945 = new_n2899 & ~new_n15036 ;
  assign new_n17946 = ~new_n14472 & new_n15036 ;
  assign new_n17947 = ~new_n17945 & ~new_n17946 ;
  assign new_n17948 = new_n15033 & ~new_n17947 ;
  assign new_n17949 = ~new_n17944 & ~new_n17948 ;
  assign new_n17950 = lo0402 & ~new_n14943 ;
  assign new_n17951 = new_n2899 & ~new_n14946 ;
  assign new_n17952 = ~new_n14472 & new_n14946 ;
  assign new_n17953 = ~new_n17951 & ~new_n17952 ;
  assign new_n17954 = new_n14943 & ~new_n17953 ;
  assign new_n17955 = ~new_n17950 & ~new_n17954 ;
  assign new_n17956 = lo0403 & ~new_n14848 ;
  assign new_n17957 = new_n2899 & ~new_n14853 ;
  assign new_n17958 = ~new_n14472 & new_n14853 ;
  assign new_n17959 = ~new_n17957 & ~new_n17958 ;
  assign new_n17960 = new_n14848 & ~new_n17959 ;
  assign new_n17961 = ~new_n17956 & ~new_n17960 ;
  assign new_n17962 = lo0404 & ~new_n14997 ;
  assign new_n17963 = new_n2899 & ~new_n15000 ;
  assign new_n17964 = ~new_n14472 & new_n15000 ;
  assign new_n17965 = ~new_n17963 & ~new_n17964 ;
  assign new_n17966 = new_n14997 & ~new_n17965 ;
  assign new_n17967 = ~new_n17962 & ~new_n17966 ;
  assign new_n17968 = lo0405 & ~new_n15090 ;
  assign new_n17969 = new_n2899 & ~new_n15093 ;
  assign new_n17970 = ~new_n14472 & new_n15093 ;
  assign new_n17971 = ~new_n17969 & ~new_n17970 ;
  assign new_n17972 = new_n15090 & ~new_n17971 ;
  assign new_n17973 = ~new_n17968 & ~new_n17972 ;
  assign new_n17974 = lo0406 & ~new_n14869 ;
  assign new_n17975 = new_n2899 & ~new_n14872 ;
  assign new_n17976 = ~new_n14472 & new_n14872 ;
  assign new_n17977 = ~new_n17975 & ~new_n17976 ;
  assign new_n17978 = new_n14869 & ~new_n17977 ;
  assign new_n17979 = ~new_n17974 & ~new_n17978 ;
  assign new_n17980 = lo0407 & ~new_n14924 ;
  assign new_n17981 = new_n2899 & ~new_n14927 ;
  assign new_n17982 = ~new_n14472 & new_n14927 ;
  assign new_n17983 = ~new_n17981 & ~new_n17982 ;
  assign new_n17984 = new_n14924 & ~new_n17983 ;
  assign new_n17985 = ~new_n17980 & ~new_n17984 ;
  assign new_n17986 = lo0408 & ~new_n15016 ;
  assign new_n17987 = new_n2899 & ~new_n15019 ;
  assign new_n17988 = ~new_n14472 & new_n15019 ;
  assign new_n17989 = ~new_n17987 & ~new_n17988 ;
  assign new_n17990 = new_n15016 & ~new_n17989 ;
  assign new_n17991 = ~new_n17986 & ~new_n17990 ;
  assign new_n17992 = lo0409 & ~new_n15071 ;
  assign new_n17993 = new_n2899 & ~new_n15074 ;
  assign new_n17994 = ~new_n14472 & new_n15074 ;
  assign new_n17995 = ~new_n17993 & ~new_n17994 ;
  assign new_n17996 = new_n15071 & ~new_n17995 ;
  assign new_n17997 = ~new_n17992 & ~new_n17996 ;
  assign new_n17998 = lo0410 & ~new_n14960 ;
  assign new_n17999 = new_n2899 & ~new_n14963 ;
  assign new_n18000 = ~new_n14472 & new_n14963 ;
  assign new_n18001 = ~new_n17999 & ~new_n18000 ;
  assign new_n18002 = new_n14960 & ~new_n18001 ;
  assign new_n18003 = ~new_n17998 & ~new_n18002 ;
  assign new_n18004 = lo0411 & ~new_n14886 ;
  assign new_n18005 = new_n2899 & ~new_n14889 ;
  assign new_n18006 = ~new_n14472 & new_n14889 ;
  assign new_n18007 = ~new_n18005 & ~new_n18006 ;
  assign new_n18008 = new_n14886 & ~new_n18007 ;
  assign new_n18009 = ~new_n18004 & ~new_n18008 ;
  assign new_n18010 = lo0412 & ~new_n15107 ;
  assign new_n18011 = new_n2899 & ~new_n15110 ;
  assign new_n18012 = ~new_n14472 & new_n15110 ;
  assign new_n18013 = ~new_n18011 & ~new_n18012 ;
  assign new_n18014 = new_n15107 & ~new_n18013 ;
  assign new_n18015 = ~new_n18010 & ~new_n18014 ;
  assign new_n18016 = lo0413 & ~new_n14903 ;
  assign new_n18017 = new_n2899 & ~new_n14906 ;
  assign new_n18018 = ~new_n14472 & new_n14906 ;
  assign new_n18019 = ~new_n18017 & ~new_n18018 ;
  assign new_n18020 = new_n14903 & ~new_n18019 ;
  assign new_n18021 = ~new_n18016 & ~new_n18020 ;
  assign new_n18022 = lo0414 & ~new_n14977 ;
  assign new_n18023 = new_n2899 & ~new_n14980 ;
  assign new_n18024 = ~new_n14472 & new_n14980 ;
  assign new_n18025 = ~new_n18023 & ~new_n18024 ;
  assign new_n18026 = new_n14977 & ~new_n18025 ;
  assign new_n18027 = ~new_n18022 & ~new_n18026 ;
  assign new_n18028 = lo0415 & ~new_n15050 ;
  assign new_n18029 = new_n2899 & ~new_n15053 ;
  assign new_n18030 = ~new_n14472 & new_n15053 ;
  assign new_n18031 = ~new_n18029 & ~new_n18030 ;
  assign new_n18032 = new_n15050 & ~new_n18031 ;
  assign new_n18033 = ~new_n18028 & ~new_n18032 ;
  assign new_n18034 = lo0416 & ~new_n15124 ;
  assign new_n18035 = new_n2899 & ~new_n15127 ;
  assign new_n18036 = ~new_n14472 & new_n15127 ;
  assign new_n18037 = ~new_n18035 & ~new_n18036 ;
  assign new_n18038 = new_n15124 & ~new_n18037 ;
  assign new_n18039 = ~new_n18034 & ~new_n18038 ;
  assign new_n18040 = lo0417 & new_n15454 ;
  assign new_n18041 = lo0958 & ~new_n14472 ;
  assign new_n18042 = ~lo0958 & ~new_n14475 ;
  assign new_n18043 = ~new_n18041 & ~new_n18042 ;
  assign new_n18044 = ~new_n15454 & ~new_n18043 ;
  assign new_n18045 = ~new_n18040 & ~new_n18044 ;
  assign new_n18046 = lo0418 & ~new_n15365 ;
  assign new_n18047 = lo0952 & ~new_n14472 ;
  assign new_n18048 = ~lo0952 & new_n2899 ;
  assign new_n18049 = ~new_n18047 & ~new_n18048 ;
  assign new_n18050 = new_n15365 & ~new_n18049 ;
  assign new_n18051 = ~new_n18046 & ~new_n18050 ;
  assign new_n18052 = lo0419 & ~new_n14943 ;
  assign new_n18053 = ~new_n3372 & ~new_n14946 ;
  assign new_n18054 = ~new_n14499 & new_n14946 ;
  assign new_n18055 = ~new_n18053 & ~new_n18054 ;
  assign new_n18056 = new_n14943 & ~new_n18055 ;
  assign new_n18057 = ~new_n18052 & ~new_n18056 ;
  assign new_n18058 = lo0420 & ~new_n14924 ;
  assign new_n18059 = ~new_n3372 & ~new_n14927 ;
  assign new_n18060 = ~new_n14499 & new_n14927 ;
  assign new_n18061 = ~new_n18059 & ~new_n18060 ;
  assign new_n18062 = new_n14924 & ~new_n18061 ;
  assign new_n18063 = ~new_n18058 & ~new_n18062 ;
  assign new_n18064 = lo0421 & ~new_n14960 ;
  assign new_n18065 = ~new_n3372 & ~new_n14963 ;
  assign new_n18066 = ~new_n14499 & new_n14963 ;
  assign new_n18067 = ~new_n18065 & ~new_n18066 ;
  assign new_n18068 = new_n14960 & ~new_n18067 ;
  assign new_n18069 = ~new_n18064 & ~new_n18068 ;
  assign new_n18070 = lo0422 & ~new_n14977 ;
  assign new_n18071 = ~new_n3372 & ~new_n14980 ;
  assign new_n18072 = ~new_n14499 & new_n14980 ;
  assign new_n18073 = ~new_n18071 & ~new_n18072 ;
  assign new_n18074 = new_n14977 & ~new_n18073 ;
  assign new_n18075 = ~new_n18070 & ~new_n18074 ;
  assign new_n18076 = lo0423 & ~new_n14869 ;
  assign new_n18077 = ~new_n3372 & ~new_n14872 ;
  assign new_n18078 = ~new_n14499 & new_n14872 ;
  assign new_n18079 = ~new_n18077 & ~new_n18078 ;
  assign new_n18080 = new_n14869 & ~new_n18079 ;
  assign new_n18081 = ~new_n18076 & ~new_n18080 ;
  assign new_n18082 = lo0424 & ~new_n14848 ;
  assign new_n18083 = ~new_n3372 & ~new_n14853 ;
  assign new_n18084 = ~new_n14499 & new_n14853 ;
  assign new_n18085 = ~new_n18083 & ~new_n18084 ;
  assign new_n18086 = new_n14848 & ~new_n18085 ;
  assign new_n18087 = ~new_n18082 & ~new_n18086 ;
  assign new_n18088 = lo0425 & ~new_n14886 ;
  assign new_n18089 = ~new_n3372 & ~new_n14889 ;
  assign new_n18090 = ~new_n14499 & new_n14889 ;
  assign new_n18091 = ~new_n18089 & ~new_n18090 ;
  assign new_n18092 = new_n14886 & ~new_n18091 ;
  assign new_n18093 = ~new_n18088 & ~new_n18092 ;
  assign new_n18094 = lo0426 & ~new_n14903 ;
  assign new_n18095 = ~new_n3372 & ~new_n14906 ;
  assign new_n18096 = ~new_n14499 & new_n14906 ;
  assign new_n18097 = ~new_n18095 & ~new_n18096 ;
  assign new_n18098 = new_n14903 & ~new_n18097 ;
  assign new_n18099 = ~new_n18094 & ~new_n18098 ;
  assign new_n18100 = lo0427 & ~new_n15016 ;
  assign new_n18101 = ~new_n3372 & ~new_n15019 ;
  assign new_n18102 = ~new_n14499 & new_n15019 ;
  assign new_n18103 = ~new_n18101 & ~new_n18102 ;
  assign new_n18104 = new_n15016 & ~new_n18103 ;
  assign new_n18105 = ~new_n18100 & ~new_n18104 ;
  assign new_n18106 = lo0428 & ~new_n14997 ;
  assign new_n18107 = ~new_n3372 & ~new_n15000 ;
  assign new_n18108 = ~new_n14499 & new_n15000 ;
  assign new_n18109 = ~new_n18107 & ~new_n18108 ;
  assign new_n18110 = new_n14997 & ~new_n18109 ;
  assign new_n18111 = ~new_n18106 & ~new_n18110 ;
  assign new_n18112 = lo0429 & ~new_n15033 ;
  assign new_n18113 = ~new_n3372 & ~new_n15036 ;
  assign new_n18114 = ~new_n14499 & new_n15036 ;
  assign new_n18115 = ~new_n18113 & ~new_n18114 ;
  assign new_n18116 = new_n15033 & ~new_n18115 ;
  assign new_n18117 = ~new_n18112 & ~new_n18116 ;
  assign new_n18118 = lo0430 & ~new_n15050 ;
  assign new_n18119 = ~new_n3372 & ~new_n15053 ;
  assign new_n18120 = ~new_n14499 & new_n15053 ;
  assign new_n18121 = ~new_n18119 & ~new_n18120 ;
  assign new_n18122 = new_n15050 & ~new_n18121 ;
  assign new_n18123 = ~new_n18118 & ~new_n18122 ;
  assign new_n18124 = lo0431 & ~new_n15090 ;
  assign new_n18125 = ~new_n3372 & ~new_n15093 ;
  assign new_n18126 = ~new_n14499 & new_n15093 ;
  assign new_n18127 = ~new_n18125 & ~new_n18126 ;
  assign new_n18128 = new_n15090 & ~new_n18127 ;
  assign new_n18129 = ~new_n18124 & ~new_n18128 ;
  assign new_n18130 = lo0432 & ~new_n15071 ;
  assign new_n18131 = ~new_n3372 & ~new_n15074 ;
  assign new_n18132 = ~new_n14499 & new_n15074 ;
  assign new_n18133 = ~new_n18131 & ~new_n18132 ;
  assign new_n18134 = new_n15071 & ~new_n18133 ;
  assign new_n18135 = ~new_n18130 & ~new_n18134 ;
  assign new_n18136 = lo0433 & ~new_n15107 ;
  assign new_n18137 = ~new_n3372 & ~new_n15110 ;
  assign new_n18138 = ~new_n14499 & new_n15110 ;
  assign new_n18139 = ~new_n18137 & ~new_n18138 ;
  assign new_n18140 = new_n15107 & ~new_n18139 ;
  assign new_n18141 = ~new_n18136 & ~new_n18140 ;
  assign new_n18142 = lo0434 & ~new_n15124 ;
  assign new_n18143 = ~new_n3372 & ~new_n15127 ;
  assign new_n18144 = ~new_n14499 & new_n15127 ;
  assign new_n18145 = ~new_n18143 & ~new_n18144 ;
  assign new_n18146 = new_n15124 & ~new_n18145 ;
  assign new_n18147 = ~new_n18142 & ~new_n18146 ;
  assign new_n18148 = lo0435 & ~new_n15137 ;
  assign new_n18149 = new_n15137 & ~new_n15749 ;
  assign new_n18150 = ~new_n18148 & ~new_n18149 ;
  assign new_n18151 = lo0436 & ~new_n15137 ;
  assign new_n18152 = new_n15137 & ~new_n15771 ;
  assign new_n18153 = ~new_n18151 & ~new_n18152 ;
  assign new_n18154 = lo0437 & new_n15454 ;
  assign new_n18155 = lo0958 & ~new_n14499 ;
  assign new_n18156 = ~lo0958 & ~new_n14503 ;
  assign new_n18157 = ~new_n18155 & ~new_n18156 ;
  assign new_n18158 = ~new_n15454 & ~new_n18157 ;
  assign new_n18159 = ~new_n18154 & ~new_n18158 ;
  assign new_n18160 = lo0438 & ~new_n15365 ;
  assign new_n18161 = lo0952 & ~new_n14499 ;
  assign new_n18162 = ~lo0952 & ~new_n3372 ;
  assign new_n18163 = ~new_n18161 & ~new_n18162 ;
  assign new_n18164 = new_n15365 & ~new_n18163 ;
  assign new_n18165 = ~new_n18160 & ~new_n18164 ;
  assign new_n18166 = lo0439 & ~new_n17223 ;
  assign new_n18167 = ~new_n14499 & new_n17223 ;
  assign new_n18168 = ~new_n18166 & ~new_n18167 ;
  assign new_n18169 = lo0440 & ~new_n14943 ;
  assign new_n18170 = new_n2990 & ~new_n14946 ;
  assign new_n18171 = ~new_n14128 & new_n14946 ;
  assign new_n18172 = ~new_n18170 & ~new_n18171 ;
  assign new_n18173 = new_n14943 & ~new_n18172 ;
  assign new_n18174 = ~new_n18169 & ~new_n18173 ;
  assign new_n18175 = lo0441 & ~new_n14924 ;
  assign new_n18176 = new_n2990 & ~new_n14927 ;
  assign new_n18177 = ~new_n14128 & new_n14927 ;
  assign new_n18178 = ~new_n18176 & ~new_n18177 ;
  assign new_n18179 = new_n14924 & ~new_n18178 ;
  assign new_n18180 = ~new_n18175 & ~new_n18179 ;
  assign new_n18181 = lo0442 & ~new_n14960 ;
  assign new_n18182 = new_n2990 & ~new_n14963 ;
  assign new_n18183 = ~new_n14128 & new_n14963 ;
  assign new_n18184 = ~new_n18182 & ~new_n18183 ;
  assign new_n18185 = new_n14960 & ~new_n18184 ;
  assign new_n18186 = ~new_n18181 & ~new_n18185 ;
  assign new_n18187 = lo0443 & ~new_n14977 ;
  assign new_n18188 = new_n2990 & ~new_n14980 ;
  assign new_n18189 = ~new_n14128 & new_n14980 ;
  assign new_n18190 = ~new_n18188 & ~new_n18189 ;
  assign new_n18191 = new_n14977 & ~new_n18190 ;
  assign new_n18192 = ~new_n18187 & ~new_n18191 ;
  assign new_n18193 = lo0444 & ~new_n14869 ;
  assign new_n18194 = new_n2990 & ~new_n14872 ;
  assign new_n18195 = ~new_n14128 & new_n14872 ;
  assign new_n18196 = ~new_n18194 & ~new_n18195 ;
  assign new_n18197 = new_n14869 & ~new_n18196 ;
  assign new_n18198 = ~new_n18193 & ~new_n18197 ;
  assign new_n18199 = lo0445 & ~new_n14848 ;
  assign new_n18200 = new_n2990 & ~new_n14853 ;
  assign new_n18201 = ~new_n14128 & new_n14853 ;
  assign new_n18202 = ~new_n18200 & ~new_n18201 ;
  assign new_n18203 = new_n14848 & ~new_n18202 ;
  assign new_n18204 = ~new_n18199 & ~new_n18203 ;
  assign new_n18205 = lo0446 & ~new_n14886 ;
  assign new_n18206 = new_n2990 & ~new_n14889 ;
  assign new_n18207 = ~new_n14128 & new_n14889 ;
  assign new_n18208 = ~new_n18206 & ~new_n18207 ;
  assign new_n18209 = new_n14886 & ~new_n18208 ;
  assign new_n18210 = ~new_n18205 & ~new_n18209 ;
  assign new_n18211 = lo0447 & ~new_n14903 ;
  assign new_n18212 = new_n2990 & ~new_n14906 ;
  assign new_n18213 = ~new_n14128 & new_n14906 ;
  assign new_n18214 = ~new_n18212 & ~new_n18213 ;
  assign new_n18215 = new_n14903 & ~new_n18214 ;
  assign new_n18216 = ~new_n18211 & ~new_n18215 ;
  assign new_n18217 = lo0448 & ~new_n15016 ;
  assign new_n18218 = new_n2990 & ~new_n15019 ;
  assign new_n18219 = ~new_n14128 & new_n15019 ;
  assign new_n18220 = ~new_n18218 & ~new_n18219 ;
  assign new_n18221 = new_n15016 & ~new_n18220 ;
  assign new_n18222 = ~new_n18217 & ~new_n18221 ;
  assign new_n18223 = lo0449 & ~new_n14997 ;
  assign new_n18224 = new_n2990 & ~new_n15000 ;
  assign new_n18225 = ~new_n14128 & new_n15000 ;
  assign new_n18226 = ~new_n18224 & ~new_n18225 ;
  assign new_n18227 = new_n14997 & ~new_n18226 ;
  assign new_n18228 = ~new_n18223 & ~new_n18227 ;
  assign new_n18229 = lo0450 & ~new_n15033 ;
  assign new_n18230 = new_n2990 & ~new_n15036 ;
  assign new_n18231 = ~new_n14128 & new_n15036 ;
  assign new_n18232 = ~new_n18230 & ~new_n18231 ;
  assign new_n18233 = new_n15033 & ~new_n18232 ;
  assign new_n18234 = ~new_n18229 & ~new_n18233 ;
  assign new_n18235 = lo0451 & ~new_n15050 ;
  assign new_n18236 = new_n2990 & ~new_n15053 ;
  assign new_n18237 = ~new_n14128 & new_n15053 ;
  assign new_n18238 = ~new_n18236 & ~new_n18237 ;
  assign new_n18239 = new_n15050 & ~new_n18238 ;
  assign new_n18240 = ~new_n18235 & ~new_n18239 ;
  assign new_n18241 = lo0452 & ~new_n15090 ;
  assign new_n18242 = new_n2990 & ~new_n15093 ;
  assign new_n18243 = ~new_n14128 & new_n15093 ;
  assign new_n18244 = ~new_n18242 & ~new_n18243 ;
  assign new_n18245 = new_n15090 & ~new_n18244 ;
  assign new_n18246 = ~new_n18241 & ~new_n18245 ;
  assign new_n18247 = lo0453 & ~new_n15071 ;
  assign new_n18248 = new_n2990 & ~new_n15074 ;
  assign new_n18249 = ~new_n14128 & new_n15074 ;
  assign new_n18250 = ~new_n18248 & ~new_n18249 ;
  assign new_n18251 = new_n15071 & ~new_n18250 ;
  assign new_n18252 = ~new_n18247 & ~new_n18251 ;
  assign new_n18253 = lo0454 & ~new_n15107 ;
  assign new_n18254 = new_n2990 & ~new_n15110 ;
  assign new_n18255 = ~new_n14128 & new_n15110 ;
  assign new_n18256 = ~new_n18254 & ~new_n18255 ;
  assign new_n18257 = new_n15107 & ~new_n18256 ;
  assign new_n18258 = ~new_n18253 & ~new_n18257 ;
  assign new_n18259 = lo0455 & ~new_n15124 ;
  assign new_n18260 = new_n2990 & ~new_n15127 ;
  assign new_n18261 = ~new_n14128 & new_n15127 ;
  assign new_n18262 = ~new_n18260 & ~new_n18261 ;
  assign new_n18263 = new_n15124 & ~new_n18262 ;
  assign new_n18264 = ~new_n18259 & ~new_n18263 ;
  assign new_n18265 = lo0456 & ~new_n15137 ;
  assign new_n18266 = new_n15137 & ~new_n16127 ;
  assign new_n18267 = ~new_n18265 & ~new_n18266 ;
  assign new_n18268 = lo0457 & new_n15454 ;
  assign new_n18269 = lo0958 & ~new_n14128 ;
  assign new_n18270 = ~lo0958 & ~new_n14132 ;
  assign new_n18271 = ~new_n18269 & ~new_n18270 ;
  assign new_n18272 = ~new_n15454 & ~new_n18271 ;
  assign new_n18273 = ~new_n18268 & ~new_n18272 ;
  assign new_n18274 = lo0458 & ~new_n15365 ;
  assign new_n18275 = lo0952 & ~new_n14128 ;
  assign new_n18276 = ~lo0952 & new_n2990 ;
  assign new_n18277 = ~new_n18275 & ~new_n18276 ;
  assign new_n18278 = new_n15365 & ~new_n18277 ;
  assign new_n18279 = ~new_n18274 & ~new_n18278 ;
  assign new_n18280 = lo0459 & ~new_n17223 ;
  assign new_n18281 = ~new_n14128 & new_n17223 ;
  assign new_n18282 = ~new_n18280 & ~new_n18281 ;
  assign new_n18283 = lo0460 & ~new_n14848 ;
  assign new_n18284 = new_n2718 & ~new_n14853 ;
  assign new_n18285 = ~new_n14060 & new_n14853 ;
  assign new_n18286 = ~new_n18284 & ~new_n18285 ;
  assign new_n18287 = new_n14848 & ~new_n18286 ;
  assign new_n18288 = ~new_n18283 & ~new_n18287 ;
  assign new_n18289 = lo0461 & ~new_n14869 ;
  assign new_n18290 = new_n2718 & ~new_n14872 ;
  assign new_n18291 = ~new_n14060 & new_n14872 ;
  assign new_n18292 = ~new_n18290 & ~new_n18291 ;
  assign new_n18293 = new_n14869 & ~new_n18292 ;
  assign new_n18294 = ~new_n18289 & ~new_n18293 ;
  assign new_n18295 = lo0462 & ~new_n14886 ;
  assign new_n18296 = new_n2718 & ~new_n14889 ;
  assign new_n18297 = ~new_n14060 & new_n14889 ;
  assign new_n18298 = ~new_n18296 & ~new_n18297 ;
  assign new_n18299 = new_n14886 & ~new_n18298 ;
  assign new_n18300 = ~new_n18295 & ~new_n18299 ;
  assign new_n18301 = lo0463 & ~new_n14903 ;
  assign new_n18302 = new_n2718 & ~new_n14906 ;
  assign new_n18303 = ~new_n14060 & new_n14906 ;
  assign new_n18304 = ~new_n18302 & ~new_n18303 ;
  assign new_n18305 = new_n14903 & ~new_n18304 ;
  assign new_n18306 = ~new_n18301 & ~new_n18305 ;
  assign new_n18307 = lo0464 & ~new_n14924 ;
  assign new_n18308 = new_n2718 & ~new_n14927 ;
  assign new_n18309 = ~new_n14060 & new_n14927 ;
  assign new_n18310 = ~new_n18308 & ~new_n18309 ;
  assign new_n18311 = new_n14924 & ~new_n18310 ;
  assign new_n18312 = ~new_n18307 & ~new_n18311 ;
  assign new_n18313 = lo0465 & ~new_n14943 ;
  assign new_n18314 = new_n2718 & ~new_n14946 ;
  assign new_n18315 = ~new_n14060 & new_n14946 ;
  assign new_n18316 = ~new_n18314 & ~new_n18315 ;
  assign new_n18317 = new_n14943 & ~new_n18316 ;
  assign new_n18318 = ~new_n18313 & ~new_n18317 ;
  assign new_n18319 = lo0466 & ~new_n14960 ;
  assign new_n18320 = new_n2718 & ~new_n14963 ;
  assign new_n18321 = ~new_n14060 & new_n14963 ;
  assign new_n18322 = ~new_n18320 & ~new_n18321 ;
  assign new_n18323 = new_n14960 & ~new_n18322 ;
  assign new_n18324 = ~new_n18319 & ~new_n18323 ;
  assign new_n18325 = lo0467 & ~new_n14977 ;
  assign new_n18326 = new_n2718 & ~new_n14980 ;
  assign new_n18327 = ~new_n14060 & new_n14980 ;
  assign new_n18328 = ~new_n18326 & ~new_n18327 ;
  assign new_n18329 = new_n14977 & ~new_n18328 ;
  assign new_n18330 = ~new_n18325 & ~new_n18329 ;
  assign new_n18331 = lo0468 & ~new_n14997 ;
  assign new_n18332 = new_n2718 & ~new_n15000 ;
  assign new_n18333 = ~new_n14060 & new_n15000 ;
  assign new_n18334 = ~new_n18332 & ~new_n18333 ;
  assign new_n18335 = new_n14997 & ~new_n18334 ;
  assign new_n18336 = ~new_n18331 & ~new_n18335 ;
  assign new_n18337 = lo0469 & ~new_n15016 ;
  assign new_n18338 = new_n2718 & ~new_n15019 ;
  assign new_n18339 = ~new_n14060 & new_n15019 ;
  assign new_n18340 = ~new_n18338 & ~new_n18339 ;
  assign new_n18341 = new_n15016 & ~new_n18340 ;
  assign new_n18342 = ~new_n18337 & ~new_n18341 ;
  assign new_n18343 = lo0470 & ~new_n15033 ;
  assign new_n18344 = new_n2718 & ~new_n15036 ;
  assign new_n18345 = ~new_n14060 & new_n15036 ;
  assign new_n18346 = ~new_n18344 & ~new_n18345 ;
  assign new_n18347 = new_n15033 & ~new_n18346 ;
  assign new_n18348 = ~new_n18343 & ~new_n18347 ;
  assign new_n18349 = lo0471 & ~new_n15050 ;
  assign new_n18350 = new_n2718 & ~new_n15053 ;
  assign new_n18351 = ~new_n14060 & new_n15053 ;
  assign new_n18352 = ~new_n18350 & ~new_n18351 ;
  assign new_n18353 = new_n15050 & ~new_n18352 ;
  assign new_n18354 = ~new_n18349 & ~new_n18353 ;
  assign new_n18355 = lo0472 & ~new_n15071 ;
  assign new_n18356 = new_n2718 & ~new_n15074 ;
  assign new_n18357 = ~new_n14060 & new_n15074 ;
  assign new_n18358 = ~new_n18356 & ~new_n18357 ;
  assign new_n18359 = new_n15071 & ~new_n18358 ;
  assign new_n18360 = ~new_n18355 & ~new_n18359 ;
  assign new_n18361 = lo0473 & ~new_n15090 ;
  assign new_n18362 = new_n2718 & ~new_n15093 ;
  assign new_n18363 = ~new_n14060 & new_n15093 ;
  assign new_n18364 = ~new_n18362 & ~new_n18363 ;
  assign new_n18365 = new_n15090 & ~new_n18364 ;
  assign new_n18366 = ~new_n18361 & ~new_n18365 ;
  assign new_n18367 = lo0474 & ~new_n15107 ;
  assign new_n18368 = new_n2718 & ~new_n15110 ;
  assign new_n18369 = ~new_n14060 & new_n15110 ;
  assign new_n18370 = ~new_n18368 & ~new_n18369 ;
  assign new_n18371 = new_n15107 & ~new_n18370 ;
  assign new_n18372 = ~new_n18367 & ~new_n18371 ;
  assign new_n18373 = lo0475 & ~new_n15124 ;
  assign new_n18374 = new_n2718 & ~new_n15127 ;
  assign new_n18375 = ~new_n14060 & new_n15127 ;
  assign new_n18376 = ~new_n18374 & ~new_n18375 ;
  assign new_n18377 = new_n15124 & ~new_n18376 ;
  assign new_n18378 = ~new_n18373 & ~new_n18377 ;
  assign new_n18379 = lo0476 & new_n15454 ;
  assign new_n18380 = lo0958 & ~new_n14060 ;
  assign new_n18381 = ~lo0958 & ~new_n14079 ;
  assign new_n18382 = ~new_n18380 & ~new_n18381 ;
  assign new_n18383 = ~new_n15454 & ~new_n18382 ;
  assign new_n18384 = ~new_n18379 & ~new_n18383 ;
  assign new_n18385 = lo0477 & ~new_n15365 ;
  assign new_n18386 = lo0952 & ~new_n14060 ;
  assign new_n18387 = ~lo0952 & new_n2718 ;
  assign new_n18388 = ~new_n18386 & ~new_n18387 ;
  assign new_n18389 = new_n15365 & ~new_n18388 ;
  assign new_n18390 = ~new_n18385 & ~new_n18389 ;
  assign new_n18391 = lo0478 & ~new_n17223 ;
  assign new_n18392 = ~new_n14060 & new_n17223 ;
  assign new_n18393 = ~new_n18391 & ~new_n18392 ;
  assign new_n18394 = lo0479 & ~new_n14943 ;
  assign new_n18395 = new_n3081 & ~new_n14946 ;
  assign new_n18396 = ~new_n14101 & new_n14946 ;
  assign new_n18397 = ~new_n18395 & ~new_n18396 ;
  assign new_n18398 = new_n14943 & ~new_n18397 ;
  assign new_n18399 = ~new_n18394 & ~new_n18398 ;
  assign new_n18400 = lo0480 & ~new_n14848 ;
  assign new_n18401 = new_n3081 & ~new_n14853 ;
  assign new_n18402 = ~new_n14101 & new_n14853 ;
  assign new_n18403 = ~new_n18401 & ~new_n18402 ;
  assign new_n18404 = new_n14848 & ~new_n18403 ;
  assign new_n18405 = ~new_n18400 & ~new_n18404 ;
  assign new_n18406 = lo0481 & ~new_n14997 ;
  assign new_n18407 = new_n3081 & ~new_n15000 ;
  assign new_n18408 = ~new_n14101 & new_n15000 ;
  assign new_n18409 = ~new_n18407 & ~new_n18408 ;
  assign new_n18410 = new_n14997 & ~new_n18409 ;
  assign new_n18411 = ~new_n18406 & ~new_n18410 ;
  assign new_n18412 = lo0482 & ~new_n15090 ;
  assign new_n18413 = new_n3081 & ~new_n15093 ;
  assign new_n18414 = ~new_n14101 & new_n15093 ;
  assign new_n18415 = ~new_n18413 & ~new_n18414 ;
  assign new_n18416 = new_n15090 & ~new_n18415 ;
  assign new_n18417 = ~new_n18412 & ~new_n18416 ;
  assign new_n18418 = lo0483 & ~new_n14869 ;
  assign new_n18419 = new_n3081 & ~new_n14872 ;
  assign new_n18420 = ~new_n14101 & new_n14872 ;
  assign new_n18421 = ~new_n18419 & ~new_n18420 ;
  assign new_n18422 = new_n14869 & ~new_n18421 ;
  assign new_n18423 = ~new_n18418 & ~new_n18422 ;
  assign new_n18424 = lo0484 & ~new_n14924 ;
  assign new_n18425 = new_n3081 & ~new_n14927 ;
  assign new_n18426 = ~new_n14101 & new_n14927 ;
  assign new_n18427 = ~new_n18425 & ~new_n18426 ;
  assign new_n18428 = new_n14924 & ~new_n18427 ;
  assign new_n18429 = ~new_n18424 & ~new_n18428 ;
  assign new_n18430 = lo0485 & ~new_n15016 ;
  assign new_n18431 = new_n3081 & ~new_n15019 ;
  assign new_n18432 = ~new_n14101 & new_n15019 ;
  assign new_n18433 = ~new_n18431 & ~new_n18432 ;
  assign new_n18434 = new_n15016 & ~new_n18433 ;
  assign new_n18435 = ~new_n18430 & ~new_n18434 ;
  assign new_n18436 = lo0486 & ~new_n15071 ;
  assign new_n18437 = new_n3081 & ~new_n15074 ;
  assign new_n18438 = ~new_n14101 & new_n15074 ;
  assign new_n18439 = ~new_n18437 & ~new_n18438 ;
  assign new_n18440 = new_n15071 & ~new_n18439 ;
  assign new_n18441 = ~new_n18436 & ~new_n18440 ;
  assign new_n18442 = lo0487 & ~new_n14960 ;
  assign new_n18443 = new_n3081 & ~new_n14963 ;
  assign new_n18444 = ~new_n14101 & new_n14963 ;
  assign new_n18445 = ~new_n18443 & ~new_n18444 ;
  assign new_n18446 = new_n14960 & ~new_n18445 ;
  assign new_n18447 = ~new_n18442 & ~new_n18446 ;
  assign new_n18448 = lo0488 & ~new_n14886 ;
  assign new_n18449 = new_n3081 & ~new_n14889 ;
  assign new_n18450 = ~new_n14101 & new_n14889 ;
  assign new_n18451 = ~new_n18449 & ~new_n18450 ;
  assign new_n18452 = new_n14886 & ~new_n18451 ;
  assign new_n18453 = ~new_n18448 & ~new_n18452 ;
  assign new_n18454 = lo0489 & ~new_n15033 ;
  assign new_n18455 = new_n3081 & ~new_n15036 ;
  assign new_n18456 = ~new_n14101 & new_n15036 ;
  assign new_n18457 = ~new_n18455 & ~new_n18456 ;
  assign new_n18458 = new_n15033 & ~new_n18457 ;
  assign new_n18459 = ~new_n18454 & ~new_n18458 ;
  assign new_n18460 = lo0490 & ~new_n15107 ;
  assign new_n18461 = new_n3081 & ~new_n15110 ;
  assign new_n18462 = ~new_n14101 & new_n15110 ;
  assign new_n18463 = ~new_n18461 & ~new_n18462 ;
  assign new_n18464 = new_n15107 & ~new_n18463 ;
  assign new_n18465 = ~new_n18460 & ~new_n18464 ;
  assign new_n18466 = lo0491 & ~new_n14903 ;
  assign new_n18467 = new_n3081 & ~new_n14906 ;
  assign new_n18468 = ~new_n14101 & new_n14906 ;
  assign new_n18469 = ~new_n18467 & ~new_n18468 ;
  assign new_n18470 = new_n14903 & ~new_n18469 ;
  assign new_n18471 = ~new_n18466 & ~new_n18470 ;
  assign new_n18472 = lo0492 & ~new_n14977 ;
  assign new_n18473 = new_n3081 & ~new_n14980 ;
  assign new_n18474 = ~new_n14101 & new_n14980 ;
  assign new_n18475 = ~new_n18473 & ~new_n18474 ;
  assign new_n18476 = new_n14977 & ~new_n18475 ;
  assign new_n18477 = ~new_n18472 & ~new_n18476 ;
  assign new_n18478 = lo0493 & ~new_n15050 ;
  assign new_n18479 = new_n3081 & ~new_n15053 ;
  assign new_n18480 = ~new_n14101 & new_n15053 ;
  assign new_n18481 = ~new_n18479 & ~new_n18480 ;
  assign new_n18482 = new_n15050 & ~new_n18481 ;
  assign new_n18483 = ~new_n18478 & ~new_n18482 ;
  assign new_n18484 = lo0494 & ~new_n15124 ;
  assign new_n18485 = new_n3081 & ~new_n15127 ;
  assign new_n18486 = ~new_n14101 & new_n15127 ;
  assign new_n18487 = ~new_n18485 & ~new_n18486 ;
  assign new_n18488 = new_n15124 & ~new_n18487 ;
  assign new_n18489 = ~new_n18484 & ~new_n18488 ;
  assign new_n18490 = lo0495 & new_n15454 ;
  assign new_n18491 = lo0958 & ~new_n14101 ;
  assign new_n18492 = ~lo0958 & ~new_n14104 ;
  assign new_n18493 = ~new_n18491 & ~new_n18492 ;
  assign new_n18494 = ~new_n15454 & ~new_n18493 ;
  assign new_n18495 = ~new_n18490 & ~new_n18494 ;
  assign new_n18496 = lo0496 & ~new_n15365 ;
  assign new_n18497 = lo0952 & ~new_n14101 ;
  assign new_n18498 = ~lo0952 & new_n3081 ;
  assign new_n18499 = ~new_n18497 & ~new_n18498 ;
  assign new_n18500 = new_n15365 & ~new_n18499 ;
  assign new_n18501 = ~new_n18496 & ~new_n18500 ;
  assign new_n18502 = lo0497 & ~new_n17223 ;
  assign new_n18503 = ~new_n14101 & new_n17223 ;
  assign new_n18504 = ~new_n18502 & ~new_n18503 ;
  assign new_n18505 = lo0498 & ~new_n15033 ;
  assign new_n18506 = new_n5977 & ~new_n15036 ;
  assign new_n18507 = new_n15036 & ~new_n16697 ;
  assign new_n18508 = ~new_n18506 & ~new_n18507 ;
  assign new_n18509 = new_n15033 & ~new_n18508 ;
  assign new_n18510 = ~new_n18505 & ~new_n18509 ;
  assign new_n18511 = lo0499 & ~new_n14943 ;
  assign new_n18512 = new_n5977 & ~new_n14946 ;
  assign new_n18513 = new_n14946 & ~new_n16697 ;
  assign new_n18514 = ~new_n18512 & ~new_n18513 ;
  assign new_n18515 = new_n14943 & ~new_n18514 ;
  assign new_n18516 = ~new_n18511 & ~new_n18515 ;
  assign new_n18517 = lo0500 & ~new_n14924 ;
  assign new_n18518 = new_n5977 & ~new_n14927 ;
  assign new_n18519 = new_n14927 & ~new_n16697 ;
  assign new_n18520 = ~new_n18518 & ~new_n18519 ;
  assign new_n18521 = new_n14924 & ~new_n18520 ;
  assign new_n18522 = ~new_n18517 & ~new_n18521 ;
  assign new_n18523 = lo0501 & ~new_n14960 ;
  assign new_n18524 = new_n5977 & ~new_n14963 ;
  assign new_n18525 = new_n14963 & ~new_n16697 ;
  assign new_n18526 = ~new_n18524 & ~new_n18525 ;
  assign new_n18527 = new_n14960 & ~new_n18526 ;
  assign new_n18528 = ~new_n18523 & ~new_n18527 ;
  assign new_n18529 = lo0502 & ~new_n14977 ;
  assign new_n18530 = new_n5977 & ~new_n14980 ;
  assign new_n18531 = new_n14980 & ~new_n16697 ;
  assign new_n18532 = ~new_n18530 & ~new_n18531 ;
  assign new_n18533 = new_n14977 & ~new_n18532 ;
  assign new_n18534 = ~new_n18529 & ~new_n18533 ;
  assign new_n18535 = lo0503 & ~new_n14869 ;
  assign new_n18536 = new_n5977 & ~new_n14872 ;
  assign new_n18537 = new_n14872 & ~new_n16697 ;
  assign new_n18538 = ~new_n18536 & ~new_n18537 ;
  assign new_n18539 = new_n14869 & ~new_n18538 ;
  assign new_n18540 = ~new_n18535 & ~new_n18539 ;
  assign new_n18541 = lo0504 & ~new_n14848 ;
  assign new_n18542 = new_n5977 & ~new_n14853 ;
  assign new_n18543 = new_n14853 & ~new_n16697 ;
  assign new_n18544 = ~new_n18542 & ~new_n18543 ;
  assign new_n18545 = new_n14848 & ~new_n18544 ;
  assign new_n18546 = ~new_n18541 & ~new_n18545 ;
  assign new_n18547 = lo0505 & ~new_n14886 ;
  assign new_n18548 = new_n5977 & ~new_n14889 ;
  assign new_n18549 = new_n14889 & ~new_n16697 ;
  assign new_n18550 = ~new_n18548 & ~new_n18549 ;
  assign new_n18551 = new_n14886 & ~new_n18550 ;
  assign new_n18552 = ~new_n18547 & ~new_n18551 ;
  assign new_n18553 = lo0506 & ~new_n14903 ;
  assign new_n18554 = new_n5977 & ~new_n14906 ;
  assign new_n18555 = new_n14906 & ~new_n16697 ;
  assign new_n18556 = ~new_n18554 & ~new_n18555 ;
  assign new_n18557 = new_n14903 & ~new_n18556 ;
  assign new_n18558 = ~new_n18553 & ~new_n18557 ;
  assign new_n18559 = lo0507 & ~new_n15016 ;
  assign new_n18560 = new_n5977 & ~new_n15019 ;
  assign new_n18561 = new_n15019 & ~new_n16697 ;
  assign new_n18562 = ~new_n18560 & ~new_n18561 ;
  assign new_n18563 = new_n15016 & ~new_n18562 ;
  assign new_n18564 = ~new_n18559 & ~new_n18563 ;
  assign new_n18565 = lo0508 & ~new_n14997 ;
  assign new_n18566 = new_n5977 & ~new_n15000 ;
  assign new_n18567 = new_n15000 & ~new_n16697 ;
  assign new_n18568 = ~new_n18566 & ~new_n18567 ;
  assign new_n18569 = new_n14997 & ~new_n18568 ;
  assign new_n18570 = ~new_n18565 & ~new_n18569 ;
  assign new_n18571 = lo0509 & ~new_n15050 ;
  assign new_n18572 = new_n5977 & ~new_n15053 ;
  assign new_n18573 = new_n15053 & ~new_n16697 ;
  assign new_n18574 = ~new_n18572 & ~new_n18573 ;
  assign new_n18575 = new_n15050 & ~new_n18574 ;
  assign new_n18576 = ~new_n18571 & ~new_n18575 ;
  assign new_n18577 = lo0510 & ~new_n15090 ;
  assign new_n18578 = new_n5977 & ~new_n15093 ;
  assign new_n18579 = new_n15093 & ~new_n16697 ;
  assign new_n18580 = ~new_n18578 & ~new_n18579 ;
  assign new_n18581 = new_n15090 & ~new_n18580 ;
  assign new_n18582 = ~new_n18577 & ~new_n18581 ;
  assign new_n18583 = lo0511 & ~new_n15071 ;
  assign new_n18584 = new_n5977 & ~new_n15074 ;
  assign new_n18585 = new_n15074 & ~new_n16697 ;
  assign new_n18586 = ~new_n18584 & ~new_n18585 ;
  assign new_n18587 = new_n15071 & ~new_n18586 ;
  assign new_n18588 = ~new_n18583 & ~new_n18587 ;
  assign new_n18589 = lo0512 & ~new_n15107 ;
  assign new_n18590 = new_n5977 & ~new_n15110 ;
  assign new_n18591 = new_n15110 & ~new_n16697 ;
  assign new_n18592 = ~new_n18590 & ~new_n18591 ;
  assign new_n18593 = new_n15107 & ~new_n18592 ;
  assign new_n18594 = ~new_n18589 & ~new_n18593 ;
  assign new_n18595 = lo0513 & ~new_n15124 ;
  assign new_n18596 = new_n5977 & ~new_n15127 ;
  assign new_n18597 = new_n15127 & ~new_n16697 ;
  assign new_n18598 = ~new_n18596 & ~new_n18597 ;
  assign new_n18599 = new_n15124 & ~new_n18598 ;
  assign new_n18600 = ~new_n18595 & ~new_n18599 ;
  assign new_n18601 = lo0514 & ~new_n15137 ;
  assign new_n18602 = new_n15137 & ~new_n16229 ;
  assign new_n18603 = ~new_n18601 & ~new_n18602 ;
  assign new_n18604 = lo0515 & ~new_n15365 ;
  assign new_n18605 = lo0952 & ~new_n16697 ;
  assign new_n18606 = ~lo0952 & new_n5977 ;
  assign new_n18607 = ~new_n18605 & ~new_n18606 ;
  assign new_n18608 = new_n15365 & ~new_n18607 ;
  assign new_n18609 = ~new_n18604 & ~new_n18608 ;
  assign new_n18610 = lo0516 & new_n15454 ;
  assign new_n18611 = lo0958 & ~new_n16697 ;
  assign new_n18612 = lo0516 & ~new_n13947 ;
  assign new_n18613 = ~lo0516 & new_n13947 ;
  assign new_n18614 = ~new_n18612 & ~new_n18613 ;
  assign new_n18615 = ~lo0958 & ~new_n18614 ;
  assign new_n18616 = ~new_n18611 & ~new_n18615 ;
  assign new_n18617 = ~new_n15454 & ~new_n18616 ;
  assign new_n18618 = ~new_n18610 & ~new_n18617 ;
  assign new_n18619 = lo0517 & ~new_n17223 ;
  assign new_n18620 = ~new_n16697 & new_n17223 ;
  assign new_n18621 = ~new_n18619 & ~new_n18620 ;
  assign new_n18622 = lo0518 & ~new_n14924 ;
  assign new_n18623 = ~new_n3723 & ~new_n14927 ;
  assign new_n18624 = ~new_n14005 & new_n14927 ;
  assign new_n18625 = ~new_n18623 & ~new_n18624 ;
  assign new_n18626 = new_n14924 & ~new_n18625 ;
  assign new_n18627 = ~new_n18622 & ~new_n18626 ;
  assign new_n18628 = lo0519 & ~new_n14869 ;
  assign new_n18629 = ~new_n3723 & ~new_n14872 ;
  assign new_n18630 = ~new_n14005 & new_n14872 ;
  assign new_n18631 = ~new_n18629 & ~new_n18630 ;
  assign new_n18632 = new_n14869 & ~new_n18631 ;
  assign new_n18633 = ~new_n18628 & ~new_n18632 ;
  assign new_n18634 = lo0520 & ~new_n15016 ;
  assign new_n18635 = ~new_n3723 & ~new_n15019 ;
  assign new_n18636 = ~new_n14005 & new_n15019 ;
  assign new_n18637 = ~new_n18635 & ~new_n18636 ;
  assign new_n18638 = new_n15016 & ~new_n18637 ;
  assign new_n18639 = ~new_n18634 & ~new_n18638 ;
  assign new_n18640 = lo0521 & ~new_n15071 ;
  assign new_n18641 = ~new_n3723 & ~new_n15074 ;
  assign new_n18642 = ~new_n14005 & new_n15074 ;
  assign new_n18643 = ~new_n18641 & ~new_n18642 ;
  assign new_n18644 = new_n15071 & ~new_n18643 ;
  assign new_n18645 = ~new_n18640 & ~new_n18644 ;
  assign new_n18646 = lo0522 & ~new_n14848 ;
  assign new_n18647 = ~new_n3723 & ~new_n14853 ;
  assign new_n18648 = ~new_n14005 & new_n14853 ;
  assign new_n18649 = ~new_n18647 & ~new_n18648 ;
  assign new_n18650 = new_n14848 & ~new_n18649 ;
  assign new_n18651 = ~new_n18646 & ~new_n18650 ;
  assign new_n18652 = lo0523 & ~new_n14943 ;
  assign new_n18653 = ~new_n3723 & ~new_n14946 ;
  assign new_n18654 = ~new_n14005 & new_n14946 ;
  assign new_n18655 = ~new_n18653 & ~new_n18654 ;
  assign new_n18656 = new_n14943 & ~new_n18655 ;
  assign new_n18657 = ~new_n18652 & ~new_n18656 ;
  assign new_n18658 = lo0524 & ~new_n14997 ;
  assign new_n18659 = ~new_n3723 & ~new_n15000 ;
  assign new_n18660 = ~new_n14005 & new_n15000 ;
  assign new_n18661 = ~new_n18659 & ~new_n18660 ;
  assign new_n18662 = new_n14997 & ~new_n18661 ;
  assign new_n18663 = ~new_n18658 & ~new_n18662 ;
  assign new_n18664 = lo0525 & ~new_n15090 ;
  assign new_n18665 = ~new_n3723 & ~new_n15093 ;
  assign new_n18666 = ~new_n14005 & new_n15093 ;
  assign new_n18667 = ~new_n18665 & ~new_n18666 ;
  assign new_n18668 = new_n15090 & ~new_n18667 ;
  assign new_n18669 = ~new_n18664 & ~new_n18668 ;
  assign new_n18670 = lo0526 & ~new_n14886 ;
  assign new_n18671 = ~new_n3723 & ~new_n14889 ;
  assign new_n18672 = ~new_n14005 & new_n14889 ;
  assign new_n18673 = ~new_n18671 & ~new_n18672 ;
  assign new_n18674 = new_n14886 & ~new_n18673 ;
  assign new_n18675 = ~new_n18670 & ~new_n18674 ;
  assign new_n18676 = lo0527 & ~new_n14960 ;
  assign new_n18677 = ~new_n3723 & ~new_n14963 ;
  assign new_n18678 = ~new_n14005 & new_n14963 ;
  assign new_n18679 = ~new_n18677 & ~new_n18678 ;
  assign new_n18680 = new_n14960 & ~new_n18679 ;
  assign new_n18681 = ~new_n18676 & ~new_n18680 ;
  assign new_n18682 = lo0528 & ~new_n15033 ;
  assign new_n18683 = ~new_n3723 & ~new_n15036 ;
  assign new_n18684 = ~new_n14005 & new_n15036 ;
  assign new_n18685 = ~new_n18683 & ~new_n18684 ;
  assign new_n18686 = new_n15033 & ~new_n18685 ;
  assign new_n18687 = ~new_n18682 & ~new_n18686 ;
  assign new_n18688 = lo0529 & ~new_n15107 ;
  assign new_n18689 = ~new_n3723 & ~new_n15110 ;
  assign new_n18690 = ~new_n14005 & new_n15110 ;
  assign new_n18691 = ~new_n18689 & ~new_n18690 ;
  assign new_n18692 = new_n15107 & ~new_n18691 ;
  assign new_n18693 = ~new_n18688 & ~new_n18692 ;
  assign new_n18694 = lo0530 & ~new_n14977 ;
  assign new_n18695 = ~new_n3723 & ~new_n14980 ;
  assign new_n18696 = ~new_n14005 & new_n14980 ;
  assign new_n18697 = ~new_n18695 & ~new_n18696 ;
  assign new_n18698 = new_n14977 & ~new_n18697 ;
  assign new_n18699 = ~new_n18694 & ~new_n18698 ;
  assign new_n18700 = lo0531 & ~new_n14903 ;
  assign new_n18701 = ~new_n3723 & ~new_n14906 ;
  assign new_n18702 = ~new_n14005 & new_n14906 ;
  assign new_n18703 = ~new_n18701 & ~new_n18702 ;
  assign new_n18704 = new_n14903 & ~new_n18703 ;
  assign new_n18705 = ~new_n18700 & ~new_n18704 ;
  assign new_n18706 = lo0532 & ~new_n15050 ;
  assign new_n18707 = ~new_n3723 & ~new_n15053 ;
  assign new_n18708 = ~new_n14005 & new_n15053 ;
  assign new_n18709 = ~new_n18707 & ~new_n18708 ;
  assign new_n18710 = new_n15050 & ~new_n18709 ;
  assign new_n18711 = ~new_n18706 & ~new_n18710 ;
  assign new_n18712 = lo0533 & ~new_n15124 ;
  assign new_n18713 = ~new_n3723 & ~new_n15127 ;
  assign new_n18714 = ~new_n14005 & new_n15127 ;
  assign new_n18715 = ~new_n18713 & ~new_n18714 ;
  assign new_n18716 = new_n15124 & ~new_n18715 ;
  assign new_n18717 = ~new_n18712 & ~new_n18716 ;
  assign new_n18718 = lo0534 & ~new_n15137 ;
  assign new_n18719 = new_n15137 & ~new_n16105 ;
  assign new_n18720 = ~new_n18718 & ~new_n18719 ;
  assign new_n18721 = lo0535 & new_n15454 ;
  assign new_n18722 = lo0958 & ~new_n14005 ;
  assign new_n18723 = ~lo0958 & ~new_n14012 ;
  assign new_n18724 = ~new_n18722 & ~new_n18723 ;
  assign new_n18725 = ~new_n15454 & ~new_n18724 ;
  assign new_n18726 = ~new_n18721 & ~new_n18725 ;
  assign new_n18727 = lo0536 & ~new_n15365 ;
  assign new_n18728 = lo0952 & ~new_n14005 ;
  assign new_n18729 = ~lo0952 & ~new_n3723 ;
  assign new_n18730 = ~new_n18728 & ~new_n18729 ;
  assign new_n18731 = new_n15365 & ~new_n18730 ;
  assign new_n18732 = ~new_n18727 & ~new_n18731 ;
  assign new_n18733 = lo0537 & ~new_n17223 ;
  assign new_n18734 = ~new_n14005 & new_n17223 ;
  assign new_n18735 = ~new_n18733 & ~new_n18734 ;
  assign new_n18736 = lo0538 & ~new_n17223 ;
  assign new_n18737 = ~new_n14472 & new_n17223 ;
  assign new_n18738 = ~new_n18736 & ~new_n18737 ;
  assign new_n18739 = lo0539 & ~new_n14924 ;
  assign new_n18740 = new_n5549 & ~new_n14927 ;
  assign new_n18741 = ~new_n14036 & new_n14927 ;
  assign new_n18742 = ~new_n18740 & ~new_n18741 ;
  assign new_n18743 = new_n14924 & ~new_n18742 ;
  assign new_n18744 = ~new_n18739 & ~new_n18743 ;
  assign new_n18745 = lo0540 & ~new_n14869 ;
  assign new_n18746 = new_n5549 & ~new_n14872 ;
  assign new_n18747 = ~new_n14036 & new_n14872 ;
  assign new_n18748 = ~new_n18746 & ~new_n18747 ;
  assign new_n18749 = new_n14869 & ~new_n18748 ;
  assign new_n18750 = ~new_n18745 & ~new_n18749 ;
  assign new_n18751 = lo0541 & ~new_n15016 ;
  assign new_n18752 = new_n5549 & ~new_n15019 ;
  assign new_n18753 = ~new_n14036 & new_n15019 ;
  assign new_n18754 = ~new_n18752 & ~new_n18753 ;
  assign new_n18755 = new_n15016 & ~new_n18754 ;
  assign new_n18756 = ~new_n18751 & ~new_n18755 ;
  assign new_n18757 = lo0542 & ~new_n15071 ;
  assign new_n18758 = new_n5549 & ~new_n15074 ;
  assign new_n18759 = ~new_n14036 & new_n15074 ;
  assign new_n18760 = ~new_n18758 & ~new_n18759 ;
  assign new_n18761 = new_n15071 & ~new_n18760 ;
  assign new_n18762 = ~new_n18757 & ~new_n18761 ;
  assign new_n18763 = lo0543 & ~new_n14848 ;
  assign new_n18764 = new_n5549 & ~new_n14853 ;
  assign new_n18765 = ~new_n14036 & new_n14853 ;
  assign new_n18766 = ~new_n18764 & ~new_n18765 ;
  assign new_n18767 = new_n14848 & ~new_n18766 ;
  assign new_n18768 = ~new_n18763 & ~new_n18767 ;
  assign new_n18769 = lo0544 & ~new_n14943 ;
  assign new_n18770 = new_n5549 & ~new_n14946 ;
  assign new_n18771 = ~new_n14036 & new_n14946 ;
  assign new_n18772 = ~new_n18770 & ~new_n18771 ;
  assign new_n18773 = new_n14943 & ~new_n18772 ;
  assign new_n18774 = ~new_n18769 & ~new_n18773 ;
  assign new_n18775 = lo0545 & ~new_n14997 ;
  assign new_n18776 = new_n5549 & ~new_n15000 ;
  assign new_n18777 = ~new_n14036 & new_n15000 ;
  assign new_n18778 = ~new_n18776 & ~new_n18777 ;
  assign new_n18779 = new_n14997 & ~new_n18778 ;
  assign new_n18780 = ~new_n18775 & ~new_n18779 ;
  assign new_n18781 = lo0546 & ~new_n15090 ;
  assign new_n18782 = new_n5549 & ~new_n15093 ;
  assign new_n18783 = ~new_n14036 & new_n15093 ;
  assign new_n18784 = ~new_n18782 & ~new_n18783 ;
  assign new_n18785 = new_n15090 & ~new_n18784 ;
  assign new_n18786 = ~new_n18781 & ~new_n18785 ;
  assign new_n18787 = lo0547 & ~new_n14886 ;
  assign new_n18788 = new_n5549 & ~new_n14889 ;
  assign new_n18789 = ~new_n14036 & new_n14889 ;
  assign new_n18790 = ~new_n18788 & ~new_n18789 ;
  assign new_n18791 = new_n14886 & ~new_n18790 ;
  assign new_n18792 = ~new_n18787 & ~new_n18791 ;
  assign new_n18793 = lo0548 & ~new_n14960 ;
  assign new_n18794 = new_n5549 & ~new_n14963 ;
  assign new_n18795 = ~new_n14036 & new_n14963 ;
  assign new_n18796 = ~new_n18794 & ~new_n18795 ;
  assign new_n18797 = new_n14960 & ~new_n18796 ;
  assign new_n18798 = ~new_n18793 & ~new_n18797 ;
  assign new_n18799 = lo0549 & ~new_n15033 ;
  assign new_n18800 = new_n5549 & ~new_n15036 ;
  assign new_n18801 = ~new_n14036 & new_n15036 ;
  assign new_n18802 = ~new_n18800 & ~new_n18801 ;
  assign new_n18803 = new_n15033 & ~new_n18802 ;
  assign new_n18804 = ~new_n18799 & ~new_n18803 ;
  assign new_n18805 = lo0550 & ~new_n15107 ;
  assign new_n18806 = new_n5549 & ~new_n15110 ;
  assign new_n18807 = ~new_n14036 & new_n15110 ;
  assign new_n18808 = ~new_n18806 & ~new_n18807 ;
  assign new_n18809 = new_n15107 & ~new_n18808 ;
  assign new_n18810 = ~new_n18805 & ~new_n18809 ;
  assign new_n18811 = lo0551 & ~new_n14977 ;
  assign new_n18812 = new_n5549 & ~new_n14980 ;
  assign new_n18813 = ~new_n14036 & new_n14980 ;
  assign new_n18814 = ~new_n18812 & ~new_n18813 ;
  assign new_n18815 = new_n14977 & ~new_n18814 ;
  assign new_n18816 = ~new_n18811 & ~new_n18815 ;
  assign new_n18817 = lo0552 & ~new_n14903 ;
  assign new_n18818 = new_n5549 & ~new_n14906 ;
  assign new_n18819 = ~new_n14036 & new_n14906 ;
  assign new_n18820 = ~new_n18818 & ~new_n18819 ;
  assign new_n18821 = new_n14903 & ~new_n18820 ;
  assign new_n18822 = ~new_n18817 & ~new_n18821 ;
  assign new_n18823 = lo0553 & ~new_n15050 ;
  assign new_n18824 = new_n5549 & ~new_n15053 ;
  assign new_n18825 = ~new_n14036 & new_n15053 ;
  assign new_n18826 = ~new_n18824 & ~new_n18825 ;
  assign new_n18827 = new_n15050 & ~new_n18826 ;
  assign new_n18828 = ~new_n18823 & ~new_n18827 ;
  assign new_n18829 = lo0554 & ~new_n15124 ;
  assign new_n18830 = new_n5549 & ~new_n15127 ;
  assign new_n18831 = ~new_n14036 & new_n15127 ;
  assign new_n18832 = ~new_n18830 & ~new_n18831 ;
  assign new_n18833 = new_n15124 & ~new_n18832 ;
  assign new_n18834 = ~new_n18829 & ~new_n18833 ;
  assign new_n18835 = lo0555 & ~new_n15137 ;
  assign new_n18836 = new_n15137 & ~new_n16470 ;
  assign new_n18837 = ~new_n18835 & ~new_n18836 ;
  assign new_n18838 = lo0556 & new_n15454 ;
  assign new_n18839 = lo0958 & ~new_n14036 ;
  assign new_n18840 = ~lo0958 & ~new_n14043 ;
  assign new_n18841 = ~new_n18839 & ~new_n18840 ;
  assign new_n18842 = ~new_n15454 & ~new_n18841 ;
  assign new_n18843 = ~new_n18838 & ~new_n18842 ;
  assign new_n18844 = lo0557 & ~new_n15365 ;
  assign new_n18845 = lo0952 & ~new_n14036 ;
  assign new_n18846 = ~lo0952 & new_n5549 ;
  assign new_n18847 = ~new_n18845 & ~new_n18846 ;
  assign new_n18848 = new_n15365 & ~new_n18847 ;
  assign new_n18849 = ~new_n18844 & ~new_n18848 ;
  assign new_n18850 = lo0558 & ~new_n17223 ;
  assign new_n18851 = ~new_n14036 & new_n17223 ;
  assign new_n18852 = ~new_n18850 & ~new_n18851 ;
  assign new_n18853 = lo0559 & ~new_n17223 ;
  assign new_n18854 = ~new_n16677 & new_n17223 ;
  assign new_n18855 = ~new_n18853 & ~new_n18854 ;
  assign new_n18856 = lo0560 & ~new_n14943 ;
  assign new_n18857 = new_n6667 & ~new_n14946 ;
  assign new_n18858 = lo0954 & new_n11792 ;
  assign new_n18859 = new_n11792 & ~new_n18858 ;
  assign new_n18860 = ~new_n8936 & ~new_n18859 ;
  assign new_n18861 = ~lo0954 & new_n8936 ;
  assign new_n18862 = ~new_n11792 & new_n18861 ;
  assign new_n18863 = ~new_n18860 & ~new_n18862 ;
  assign new_n18864 = new_n14946 & ~new_n18863 ;
  assign new_n18865 = ~new_n18857 & ~new_n18864 ;
  assign new_n18866 = new_n14943 & ~new_n18865 ;
  assign new_n18867 = ~new_n18856 & ~new_n18866 ;
  assign new_n18868 = lo0561 & ~new_n14848 ;
  assign new_n18869 = new_n6667 & ~new_n14853 ;
  assign new_n18870 = new_n14853 & ~new_n18863 ;
  assign new_n18871 = ~new_n18869 & ~new_n18870 ;
  assign new_n18872 = new_n14848 & ~new_n18871 ;
  assign new_n18873 = ~new_n18868 & ~new_n18872 ;
  assign new_n18874 = lo0562 & ~new_n14997 ;
  assign new_n18875 = new_n6667 & ~new_n15000 ;
  assign new_n18876 = new_n15000 & ~new_n18863 ;
  assign new_n18877 = ~new_n18875 & ~new_n18876 ;
  assign new_n18878 = new_n14997 & ~new_n18877 ;
  assign new_n18879 = ~new_n18874 & ~new_n18878 ;
  assign new_n18880 = lo0563 & ~new_n15090 ;
  assign new_n18881 = new_n6667 & ~new_n15093 ;
  assign new_n18882 = new_n15093 & ~new_n18863 ;
  assign new_n18883 = ~new_n18881 & ~new_n18882 ;
  assign new_n18884 = new_n15090 & ~new_n18883 ;
  assign new_n18885 = ~new_n18880 & ~new_n18884 ;
  assign new_n18886 = lo0564 & ~new_n14869 ;
  assign new_n18887 = new_n6667 & ~new_n14872 ;
  assign new_n18888 = new_n14872 & ~new_n18863 ;
  assign new_n18889 = ~new_n18887 & ~new_n18888 ;
  assign new_n18890 = new_n14869 & ~new_n18889 ;
  assign new_n18891 = ~new_n18886 & ~new_n18890 ;
  assign new_n18892 = lo0565 & ~new_n14924 ;
  assign new_n18893 = new_n6667 & ~new_n14927 ;
  assign new_n18894 = new_n14927 & ~new_n18863 ;
  assign new_n18895 = ~new_n18893 & ~new_n18894 ;
  assign new_n18896 = new_n14924 & ~new_n18895 ;
  assign new_n18897 = ~new_n18892 & ~new_n18896 ;
  assign new_n18898 = lo0566 & ~new_n15016 ;
  assign new_n18899 = new_n6667 & ~new_n15019 ;
  assign new_n18900 = new_n15019 & ~new_n18863 ;
  assign new_n18901 = ~new_n18899 & ~new_n18900 ;
  assign new_n18902 = new_n15016 & ~new_n18901 ;
  assign new_n18903 = ~new_n18898 & ~new_n18902 ;
  assign new_n18904 = lo0567 & ~new_n15071 ;
  assign new_n18905 = new_n6667 & ~new_n15074 ;
  assign new_n18906 = new_n15074 & ~new_n18863 ;
  assign new_n18907 = ~new_n18905 & ~new_n18906 ;
  assign new_n18908 = new_n15071 & ~new_n18907 ;
  assign new_n18909 = ~new_n18904 & ~new_n18908 ;
  assign new_n18910 = lo0568 & ~new_n14960 ;
  assign new_n18911 = new_n6667 & ~new_n14963 ;
  assign new_n18912 = new_n14963 & ~new_n18863 ;
  assign new_n18913 = ~new_n18911 & ~new_n18912 ;
  assign new_n18914 = new_n14960 & ~new_n18913 ;
  assign new_n18915 = ~new_n18910 & ~new_n18914 ;
  assign new_n18916 = lo0569 & ~new_n14886 ;
  assign new_n18917 = new_n6667 & ~new_n14889 ;
  assign new_n18918 = new_n14889 & ~new_n18863 ;
  assign new_n18919 = ~new_n18917 & ~new_n18918 ;
  assign new_n18920 = new_n14886 & ~new_n18919 ;
  assign new_n18921 = ~new_n18916 & ~new_n18920 ;
  assign new_n18922 = lo0570 & ~new_n15033 ;
  assign new_n18923 = new_n6667 & ~new_n15036 ;
  assign new_n18924 = new_n15036 & ~new_n18863 ;
  assign new_n18925 = ~new_n18923 & ~new_n18924 ;
  assign new_n18926 = new_n15033 & ~new_n18925 ;
  assign new_n18927 = ~new_n18922 & ~new_n18926 ;
  assign new_n18928 = lo0571 & ~new_n15107 ;
  assign new_n18929 = new_n6667 & ~new_n15110 ;
  assign new_n18930 = new_n15110 & ~new_n18863 ;
  assign new_n18931 = ~new_n18929 & ~new_n18930 ;
  assign new_n18932 = new_n15107 & ~new_n18931 ;
  assign new_n18933 = ~new_n18928 & ~new_n18932 ;
  assign new_n18934 = lo0572 & ~new_n14903 ;
  assign new_n18935 = new_n6667 & ~new_n14906 ;
  assign new_n18936 = new_n14906 & ~new_n18863 ;
  assign new_n18937 = ~new_n18935 & ~new_n18936 ;
  assign new_n18938 = new_n14903 & ~new_n18937 ;
  assign new_n18939 = ~new_n18934 & ~new_n18938 ;
  assign new_n18940 = lo0573 & ~new_n14977 ;
  assign new_n18941 = new_n6667 & ~new_n14980 ;
  assign new_n18942 = new_n14980 & ~new_n18863 ;
  assign new_n18943 = ~new_n18941 & ~new_n18942 ;
  assign new_n18944 = new_n14977 & ~new_n18943 ;
  assign new_n18945 = ~new_n18940 & ~new_n18944 ;
  assign new_n18946 = lo0574 & ~new_n15050 ;
  assign new_n18947 = new_n6667 & ~new_n15053 ;
  assign new_n18948 = new_n15053 & ~new_n18863 ;
  assign new_n18949 = ~new_n18947 & ~new_n18948 ;
  assign new_n18950 = new_n15050 & ~new_n18949 ;
  assign new_n18951 = ~new_n18946 & ~new_n18950 ;
  assign new_n18952 = lo0575 & ~new_n15124 ;
  assign new_n18953 = new_n6667 & ~new_n15127 ;
  assign new_n18954 = new_n15127 & ~new_n18863 ;
  assign new_n18955 = ~new_n18953 & ~new_n18954 ;
  assign new_n18956 = new_n15124 & ~new_n18955 ;
  assign new_n18957 = ~new_n18952 & ~new_n18956 ;
  assign new_n18958 = lo0576 & ~new_n15137 ;
  assign new_n18959 = new_n15137 & ~new_n15880 ;
  assign new_n18960 = ~new_n18958 & ~new_n18959 ;
  assign new_n18961 = lo0577 & ~new_n15137 ;
  assign new_n18962 = new_n15137 & ~new_n15858 ;
  assign new_n18963 = ~new_n18961 & ~new_n18962 ;
  assign new_n18964 = lo0578 & ~new_n15137 ;
  assign new_n18965 = new_n15137 & ~new_n15696 ;
  assign new_n18966 = ~new_n18964 & ~new_n18965 ;
  assign new_n18967 = lo0579 & new_n2252 ;
  assign new_n18968 = ~new_n2252 & ~new_n12441 ;
  assign new_n18969 = ~new_n18967 & ~new_n18968 ;
  assign new_n18970 = lo0580 & new_n15454 ;
  assign new_n18971 = lo0958 & ~new_n18863 ;
  assign new_n18972 = lo0580 & ~new_n13944 ;
  assign new_n18973 = ~lo0580 & new_n13944 ;
  assign new_n18974 = ~new_n18972 & ~new_n18973 ;
  assign new_n18975 = ~lo0958 & ~new_n18974 ;
  assign new_n18976 = ~new_n18971 & ~new_n18975 ;
  assign new_n18977 = ~new_n15454 & ~new_n18976 ;
  assign new_n18978 = ~new_n18970 & ~new_n18977 ;
  assign new_n18979 = lo0581 & ~new_n17223 ;
  assign new_n18980 = new_n17223 & ~new_n18863 ;
  assign new_n18981 = ~new_n18979 & ~new_n18980 ;
  assign new_n18982 = lo0582 & ~new_n15365 ;
  assign new_n18983 = lo0952 & ~new_n18863 ;
  assign new_n18984 = ~lo0952 & new_n6667 ;
  assign new_n18985 = ~new_n18983 & ~new_n18984 ;
  assign new_n18986 = new_n15365 & ~new_n18985 ;
  assign new_n18987 = ~new_n18982 & ~new_n18986 ;
  assign new_n18988 = lo0583 & ~new_n14924 ;
  assign new_n18989 = new_n6202 & ~new_n14927 ;
  assign new_n18990 = new_n14927 & ~new_n16716 ;
  assign new_n18991 = ~new_n18989 & ~new_n18990 ;
  assign new_n18992 = new_n14924 & ~new_n18991 ;
  assign new_n18993 = ~new_n18988 & ~new_n18992 ;
  assign new_n18994 = lo0584 & ~new_n14869 ;
  assign new_n18995 = new_n6202 & ~new_n14872 ;
  assign new_n18996 = new_n14872 & ~new_n16716 ;
  assign new_n18997 = ~new_n18995 & ~new_n18996 ;
  assign new_n18998 = new_n14869 & ~new_n18997 ;
  assign new_n18999 = ~new_n18994 & ~new_n18998 ;
  assign new_n19000 = lo0585 & ~new_n15016 ;
  assign new_n19001 = new_n6202 & ~new_n15019 ;
  assign new_n19002 = new_n15019 & ~new_n16716 ;
  assign new_n19003 = ~new_n19001 & ~new_n19002 ;
  assign new_n19004 = new_n15016 & ~new_n19003 ;
  assign new_n19005 = ~new_n19000 & ~new_n19004 ;
  assign new_n19006 = lo0586 & ~new_n15071 ;
  assign new_n19007 = new_n6202 & ~new_n15074 ;
  assign new_n19008 = new_n15074 & ~new_n16716 ;
  assign new_n19009 = ~new_n19007 & ~new_n19008 ;
  assign new_n19010 = new_n15071 & ~new_n19009 ;
  assign new_n19011 = ~new_n19006 & ~new_n19010 ;
  assign new_n19012 = lo0587 & ~new_n14848 ;
  assign new_n19013 = new_n6202 & ~new_n14853 ;
  assign new_n19014 = new_n14853 & ~new_n16716 ;
  assign new_n19015 = ~new_n19013 & ~new_n19014 ;
  assign new_n19016 = new_n14848 & ~new_n19015 ;
  assign new_n19017 = ~new_n19012 & ~new_n19016 ;
  assign new_n19018 = lo0588 & ~new_n14943 ;
  assign new_n19019 = new_n6202 & ~new_n14946 ;
  assign new_n19020 = new_n14946 & ~new_n16716 ;
  assign new_n19021 = ~new_n19019 & ~new_n19020 ;
  assign new_n19022 = new_n14943 & ~new_n19021 ;
  assign new_n19023 = ~new_n19018 & ~new_n19022 ;
  assign new_n19024 = lo0589 & ~new_n14997 ;
  assign new_n19025 = new_n6202 & ~new_n15000 ;
  assign new_n19026 = new_n15000 & ~new_n16716 ;
  assign new_n19027 = ~new_n19025 & ~new_n19026 ;
  assign new_n19028 = new_n14997 & ~new_n19027 ;
  assign new_n19029 = ~new_n19024 & ~new_n19028 ;
  assign new_n19030 = lo0590 & ~new_n15090 ;
  assign new_n19031 = new_n6202 & ~new_n15093 ;
  assign new_n19032 = new_n15093 & ~new_n16716 ;
  assign new_n19033 = ~new_n19031 & ~new_n19032 ;
  assign new_n19034 = new_n15090 & ~new_n19033 ;
  assign new_n19035 = ~new_n19030 & ~new_n19034 ;
  assign new_n19036 = lo0591 & ~new_n14886 ;
  assign new_n19037 = new_n6202 & ~new_n14889 ;
  assign new_n19038 = new_n14889 & ~new_n16716 ;
  assign new_n19039 = ~new_n19037 & ~new_n19038 ;
  assign new_n19040 = new_n14886 & ~new_n19039 ;
  assign new_n19041 = ~new_n19036 & ~new_n19040 ;
  assign new_n19042 = lo0592 & ~new_n14960 ;
  assign new_n19043 = new_n6202 & ~new_n14963 ;
  assign new_n19044 = new_n14963 & ~new_n16716 ;
  assign new_n19045 = ~new_n19043 & ~new_n19044 ;
  assign new_n19046 = new_n14960 & ~new_n19045 ;
  assign new_n19047 = ~new_n19042 & ~new_n19046 ;
  assign new_n19048 = lo0593 & ~new_n15033 ;
  assign new_n19049 = new_n6202 & ~new_n15036 ;
  assign new_n19050 = new_n15036 & ~new_n16716 ;
  assign new_n19051 = ~new_n19049 & ~new_n19050 ;
  assign new_n19052 = new_n15033 & ~new_n19051 ;
  assign new_n19053 = ~new_n19048 & ~new_n19052 ;
  assign new_n19054 = lo0594 & ~new_n15107 ;
  assign new_n19055 = new_n6202 & ~new_n15110 ;
  assign new_n19056 = new_n15110 & ~new_n16716 ;
  assign new_n19057 = ~new_n19055 & ~new_n19056 ;
  assign new_n19058 = new_n15107 & ~new_n19057 ;
  assign new_n19059 = ~new_n19054 & ~new_n19058 ;
  assign new_n19060 = lo0595 & ~new_n14977 ;
  assign new_n19061 = new_n6202 & ~new_n14980 ;
  assign new_n19062 = new_n14980 & ~new_n16716 ;
  assign new_n19063 = ~new_n19061 & ~new_n19062 ;
  assign new_n19064 = new_n14977 & ~new_n19063 ;
  assign new_n19065 = ~new_n19060 & ~new_n19064 ;
  assign new_n19066 = lo0596 & ~new_n14903 ;
  assign new_n19067 = new_n6202 & ~new_n14906 ;
  assign new_n19068 = new_n14906 & ~new_n16716 ;
  assign new_n19069 = ~new_n19067 & ~new_n19068 ;
  assign new_n19070 = new_n14903 & ~new_n19069 ;
  assign new_n19071 = ~new_n19066 & ~new_n19070 ;
  assign new_n19072 = lo0597 & ~new_n15050 ;
  assign new_n19073 = new_n6202 & ~new_n15053 ;
  assign new_n19074 = new_n15053 & ~new_n16716 ;
  assign new_n19075 = ~new_n19073 & ~new_n19074 ;
  assign new_n19076 = new_n15050 & ~new_n19075 ;
  assign new_n19077 = ~new_n19072 & ~new_n19076 ;
  assign new_n19078 = lo0598 & ~new_n15124 ;
  assign new_n19079 = new_n6202 & ~new_n15127 ;
  assign new_n19080 = new_n15127 & ~new_n16716 ;
  assign new_n19081 = ~new_n19079 & ~new_n19080 ;
  assign new_n19082 = new_n15124 & ~new_n19081 ;
  assign new_n19083 = ~new_n19078 & ~new_n19082 ;
  assign new_n19084 = lo0599 & ~new_n15137 ;
  assign new_n19085 = new_n15137 & ~new_n15973 ;
  assign new_n19086 = ~new_n19084 & ~new_n19085 ;
  assign new_n19087 = lo0600 & new_n15454 ;
  assign new_n19088 = lo0958 & ~new_n16716 ;
  assign new_n19089 = lo0600 & ~new_n13946 ;
  assign new_n19090 = ~lo0600 & new_n13946 ;
  assign new_n19091 = ~new_n19089 & ~new_n19090 ;
  assign new_n19092 = ~lo0958 & ~new_n19091 ;
  assign new_n19093 = ~new_n19088 & ~new_n19092 ;
  assign new_n19094 = ~new_n15454 & ~new_n19093 ;
  assign new_n19095 = ~new_n19087 & ~new_n19094 ;
  assign new_n19096 = lo0601 & ~new_n17223 ;
  assign new_n19097 = ~new_n16716 & new_n17223 ;
  assign new_n19098 = ~new_n19096 & ~new_n19097 ;
  assign new_n19099 = lo0602 & ~new_n15365 ;
  assign new_n19100 = lo0952 & ~new_n16716 ;
  assign new_n19101 = ~lo0952 & new_n6202 ;
  assign new_n19102 = ~new_n19100 & ~new_n19101 ;
  assign new_n19103 = new_n15365 & ~new_n19102 ;
  assign new_n19104 = ~new_n19099 & ~new_n19103 ;
  assign new_n19105 = lo0603 & ~new_n14848 ;
  assign new_n19106 = new_n2813 & ~new_n14853 ;
  assign new_n19107 = ~new_n14287 & new_n14853 ;
  assign new_n19108 = ~new_n19106 & ~new_n19107 ;
  assign new_n19109 = new_n14848 & ~new_n19108 ;
  assign new_n19110 = ~new_n19105 & ~new_n19109 ;
  assign new_n19111 = lo0604 & ~new_n14869 ;
  assign new_n19112 = new_n2813 & ~new_n14872 ;
  assign new_n19113 = ~new_n14287 & new_n14872 ;
  assign new_n19114 = ~new_n19112 & ~new_n19113 ;
  assign new_n19115 = new_n14869 & ~new_n19114 ;
  assign new_n19116 = ~new_n19111 & ~new_n19115 ;
  assign new_n19117 = lo0605 & ~new_n14886 ;
  assign new_n19118 = new_n2813 & ~new_n14889 ;
  assign new_n19119 = ~new_n14287 & new_n14889 ;
  assign new_n19120 = ~new_n19118 & ~new_n19119 ;
  assign new_n19121 = new_n14886 & ~new_n19120 ;
  assign new_n19122 = ~new_n19117 & ~new_n19121 ;
  assign new_n19123 = lo0606 & ~new_n14903 ;
  assign new_n19124 = new_n2813 & ~new_n14906 ;
  assign new_n19125 = ~new_n14287 & new_n14906 ;
  assign new_n19126 = ~new_n19124 & ~new_n19125 ;
  assign new_n19127 = new_n14903 & ~new_n19126 ;
  assign new_n19128 = ~new_n19123 & ~new_n19127 ;
  assign new_n19129 = lo0607 & ~new_n14924 ;
  assign new_n19130 = new_n2813 & ~new_n14927 ;
  assign new_n19131 = ~new_n14287 & new_n14927 ;
  assign new_n19132 = ~new_n19130 & ~new_n19131 ;
  assign new_n19133 = new_n14924 & ~new_n19132 ;
  assign new_n19134 = ~new_n19129 & ~new_n19133 ;
  assign new_n19135 = lo0608 & ~new_n14943 ;
  assign new_n19136 = new_n2813 & ~new_n14946 ;
  assign new_n19137 = ~new_n14287 & new_n14946 ;
  assign new_n19138 = ~new_n19136 & ~new_n19137 ;
  assign new_n19139 = new_n14943 & ~new_n19138 ;
  assign new_n19140 = ~new_n19135 & ~new_n19139 ;
  assign new_n19141 = lo0609 & ~new_n14960 ;
  assign new_n19142 = new_n2813 & ~new_n14963 ;
  assign new_n19143 = ~new_n14287 & new_n14963 ;
  assign new_n19144 = ~new_n19142 & ~new_n19143 ;
  assign new_n19145 = new_n14960 & ~new_n19144 ;
  assign new_n19146 = ~new_n19141 & ~new_n19145 ;
  assign new_n19147 = lo0610 & ~new_n14977 ;
  assign new_n19148 = new_n2813 & ~new_n14980 ;
  assign new_n19149 = ~new_n14287 & new_n14980 ;
  assign new_n19150 = ~new_n19148 & ~new_n19149 ;
  assign new_n19151 = new_n14977 & ~new_n19150 ;
  assign new_n19152 = ~new_n19147 & ~new_n19151 ;
  assign new_n19153 = lo0611 & ~new_n14997 ;
  assign new_n19154 = new_n2813 & ~new_n15000 ;
  assign new_n19155 = ~new_n14287 & new_n15000 ;
  assign new_n19156 = ~new_n19154 & ~new_n19155 ;
  assign new_n19157 = new_n14997 & ~new_n19156 ;
  assign new_n19158 = ~new_n19153 & ~new_n19157 ;
  assign new_n19159 = lo0612 & ~new_n15016 ;
  assign new_n19160 = new_n2813 & ~new_n15019 ;
  assign new_n19161 = ~new_n14287 & new_n15019 ;
  assign new_n19162 = ~new_n19160 & ~new_n19161 ;
  assign new_n19163 = new_n15016 & ~new_n19162 ;
  assign new_n19164 = ~new_n19159 & ~new_n19163 ;
  assign new_n19165 = lo0613 & ~new_n15033 ;
  assign new_n19166 = new_n2813 & ~new_n15036 ;
  assign new_n19167 = ~new_n14287 & new_n15036 ;
  assign new_n19168 = ~new_n19166 & ~new_n19167 ;
  assign new_n19169 = new_n15033 & ~new_n19168 ;
  assign new_n19170 = ~new_n19165 & ~new_n19169 ;
  assign new_n19171 = lo0614 & ~new_n15050 ;
  assign new_n19172 = new_n2813 & ~new_n15053 ;
  assign new_n19173 = ~new_n14287 & new_n15053 ;
  assign new_n19174 = ~new_n19172 & ~new_n19173 ;
  assign new_n19175 = new_n15050 & ~new_n19174 ;
  assign new_n19176 = ~new_n19171 & ~new_n19175 ;
  assign new_n19177 = lo0615 & ~new_n15071 ;
  assign new_n19178 = new_n2813 & ~new_n15074 ;
  assign new_n19179 = ~new_n14287 & new_n15074 ;
  assign new_n19180 = ~new_n19178 & ~new_n19179 ;
  assign new_n19181 = new_n15071 & ~new_n19180 ;
  assign new_n19182 = ~new_n19177 & ~new_n19181 ;
  assign new_n19183 = lo0616 & ~new_n15090 ;
  assign new_n19184 = new_n2813 & ~new_n15093 ;
  assign new_n19185 = ~new_n14287 & new_n15093 ;
  assign new_n19186 = ~new_n19184 & ~new_n19185 ;
  assign new_n19187 = new_n15090 & ~new_n19186 ;
  assign new_n19188 = ~new_n19183 & ~new_n19187 ;
  assign new_n19189 = lo0617 & ~new_n15107 ;
  assign new_n19190 = new_n2813 & ~new_n15110 ;
  assign new_n19191 = ~new_n14287 & new_n15110 ;
  assign new_n19192 = ~new_n19190 & ~new_n19191 ;
  assign new_n19193 = new_n15107 & ~new_n19192 ;
  assign new_n19194 = ~new_n19189 & ~new_n19193 ;
  assign new_n19195 = lo0618 & ~new_n15124 ;
  assign new_n19196 = new_n2813 & ~new_n15127 ;
  assign new_n19197 = ~new_n14287 & new_n15127 ;
  assign new_n19198 = ~new_n19196 & ~new_n19197 ;
  assign new_n19199 = new_n15124 & ~new_n19198 ;
  assign new_n19200 = ~new_n19195 & ~new_n19199 ;
  assign new_n19201 = lo0619 & new_n15454 ;
  assign new_n19202 = lo0958 & ~new_n14287 ;
  assign new_n19203 = ~lo0958 & ~new_n14291 ;
  assign new_n19204 = ~new_n19202 & ~new_n19203 ;
  assign new_n19205 = ~new_n15454 & ~new_n19204 ;
  assign new_n19206 = ~new_n19201 & ~new_n19205 ;
  assign new_n19207 = lo0620 & ~new_n15365 ;
  assign new_n19208 = lo0952 & ~new_n14287 ;
  assign new_n19209 = ~lo0952 & new_n2813 ;
  assign new_n19210 = ~new_n19208 & ~new_n19209 ;
  assign new_n19211 = new_n15365 & ~new_n19210 ;
  assign new_n19212 = ~new_n19207 & ~new_n19211 ;
  assign new_n19213 = lo0621 & ~new_n17223 ;
  assign new_n19214 = ~new_n14287 & new_n17223 ;
  assign new_n19215 = ~new_n19213 & ~new_n19214 ;
  assign new_n19216 = lo0622 & ~new_n14943 ;
  assign new_n19217 = new_n6899 & ~new_n14946 ;
  assign new_n19218 = lo0954 & new_n11892 ;
  assign new_n19219 = new_n11892 & ~new_n19218 ;
  assign new_n19220 = ~new_n9056 & ~new_n19219 ;
  assign new_n19221 = ~lo0954 & new_n9056 ;
  assign new_n19222 = ~new_n11892 & new_n19221 ;
  assign new_n19223 = ~new_n19220 & ~new_n19222 ;
  assign new_n19224 = new_n14946 & ~new_n19223 ;
  assign new_n19225 = ~new_n19217 & ~new_n19224 ;
  assign new_n19226 = new_n14943 & ~new_n19225 ;
  assign new_n19227 = ~new_n19216 & ~new_n19226 ;
  assign new_n19228 = lo0623 & ~new_n14924 ;
  assign new_n19229 = new_n6899 & ~new_n14927 ;
  assign new_n19230 = new_n14927 & ~new_n19223 ;
  assign new_n19231 = ~new_n19229 & ~new_n19230 ;
  assign new_n19232 = new_n14924 & ~new_n19231 ;
  assign new_n19233 = ~new_n19228 & ~new_n19232 ;
  assign new_n19234 = lo0624 & ~new_n14960 ;
  assign new_n19235 = new_n6899 & ~new_n14963 ;
  assign new_n19236 = new_n14963 & ~new_n19223 ;
  assign new_n19237 = ~new_n19235 & ~new_n19236 ;
  assign new_n19238 = new_n14960 & ~new_n19237 ;
  assign new_n19239 = ~new_n19234 & ~new_n19238 ;
  assign new_n19240 = lo0625 & ~new_n14977 ;
  assign new_n19241 = new_n6899 & ~new_n14980 ;
  assign new_n19242 = new_n14980 & ~new_n19223 ;
  assign new_n19243 = ~new_n19241 & ~new_n19242 ;
  assign new_n19244 = new_n14977 & ~new_n19243 ;
  assign new_n19245 = ~new_n19240 & ~new_n19244 ;
  assign new_n19246 = lo0626 & ~new_n14869 ;
  assign new_n19247 = new_n6899 & ~new_n14872 ;
  assign new_n19248 = new_n14872 & ~new_n19223 ;
  assign new_n19249 = ~new_n19247 & ~new_n19248 ;
  assign new_n19250 = new_n14869 & ~new_n19249 ;
  assign new_n19251 = ~new_n19246 & ~new_n19250 ;
  assign new_n19252 = lo0627 & ~new_n14848 ;
  assign new_n19253 = new_n6899 & ~new_n14853 ;
  assign new_n19254 = new_n14853 & ~new_n19223 ;
  assign new_n19255 = ~new_n19253 & ~new_n19254 ;
  assign new_n19256 = new_n14848 & ~new_n19255 ;
  assign new_n19257 = ~new_n19252 & ~new_n19256 ;
  assign new_n19258 = lo0628 & ~new_n14886 ;
  assign new_n19259 = new_n6899 & ~new_n14889 ;
  assign new_n19260 = new_n14889 & ~new_n19223 ;
  assign new_n19261 = ~new_n19259 & ~new_n19260 ;
  assign new_n19262 = new_n14886 & ~new_n19261 ;
  assign new_n19263 = ~new_n19258 & ~new_n19262 ;
  assign new_n19264 = lo0629 & ~new_n14903 ;
  assign new_n19265 = new_n6899 & ~new_n14906 ;
  assign new_n19266 = new_n14906 & ~new_n19223 ;
  assign new_n19267 = ~new_n19265 & ~new_n19266 ;
  assign new_n19268 = new_n14903 & ~new_n19267 ;
  assign new_n19269 = ~new_n19264 & ~new_n19268 ;
  assign new_n19270 = lo0630 & ~new_n15016 ;
  assign new_n19271 = new_n6899 & ~new_n15019 ;
  assign new_n19272 = new_n15019 & ~new_n19223 ;
  assign new_n19273 = ~new_n19271 & ~new_n19272 ;
  assign new_n19274 = new_n15016 & ~new_n19273 ;
  assign new_n19275 = ~new_n19270 & ~new_n19274 ;
  assign new_n19276 = lo0631 & ~new_n14997 ;
  assign new_n19277 = new_n6899 & ~new_n15000 ;
  assign new_n19278 = new_n15000 & ~new_n19223 ;
  assign new_n19279 = ~new_n19277 & ~new_n19278 ;
  assign new_n19280 = new_n14997 & ~new_n19279 ;
  assign new_n19281 = ~new_n19276 & ~new_n19280 ;
  assign new_n19282 = lo0632 & ~new_n15033 ;
  assign new_n19283 = new_n6899 & ~new_n15036 ;
  assign new_n19284 = new_n15036 & ~new_n19223 ;
  assign new_n19285 = ~new_n19283 & ~new_n19284 ;
  assign new_n19286 = new_n15033 & ~new_n19285 ;
  assign new_n19287 = ~new_n19282 & ~new_n19286 ;
  assign new_n19288 = lo0633 & ~new_n15050 ;
  assign new_n19289 = new_n6899 & ~new_n15053 ;
  assign new_n19290 = new_n15053 & ~new_n19223 ;
  assign new_n19291 = ~new_n19289 & ~new_n19290 ;
  assign new_n19292 = new_n15050 & ~new_n19291 ;
  assign new_n19293 = ~new_n19288 & ~new_n19292 ;
  assign new_n19294 = lo0634 & ~new_n15090 ;
  assign new_n19295 = new_n6899 & ~new_n15093 ;
  assign new_n19296 = new_n15093 & ~new_n19223 ;
  assign new_n19297 = ~new_n19295 & ~new_n19296 ;
  assign new_n19298 = new_n15090 & ~new_n19297 ;
  assign new_n19299 = ~new_n19294 & ~new_n19298 ;
  assign new_n19300 = lo0635 & ~new_n15071 ;
  assign new_n19301 = new_n6899 & ~new_n15074 ;
  assign new_n19302 = new_n15074 & ~new_n19223 ;
  assign new_n19303 = ~new_n19301 & ~new_n19302 ;
  assign new_n19304 = new_n15071 & ~new_n19303 ;
  assign new_n19305 = ~new_n19300 & ~new_n19304 ;
  assign new_n19306 = lo0636 & ~new_n15107 ;
  assign new_n19307 = new_n6899 & ~new_n15110 ;
  assign new_n19308 = new_n15110 & ~new_n19223 ;
  assign new_n19309 = ~new_n19307 & ~new_n19308 ;
  assign new_n19310 = new_n15107 & ~new_n19309 ;
  assign new_n19311 = ~new_n19306 & ~new_n19310 ;
  assign new_n19312 = lo0637 & ~new_n15124 ;
  assign new_n19313 = new_n6899 & ~new_n15127 ;
  assign new_n19314 = new_n15127 & ~new_n19223 ;
  assign new_n19315 = ~new_n19313 & ~new_n19314 ;
  assign new_n19316 = new_n15124 & ~new_n19315 ;
  assign new_n19317 = ~new_n19312 & ~new_n19316 ;
  assign new_n19318 = lo0638 & ~new_n15137 ;
  assign new_n19319 = new_n15137 & ~new_n15928 ;
  assign new_n19320 = ~new_n19318 & ~new_n19319 ;
  assign new_n19321 = lo0639 & ~new_n15137 ;
  assign new_n19322 = new_n15137 & ~new_n15906 ;
  assign new_n19323 = ~new_n19321 & ~new_n19322 ;
  assign new_n19324 = lo0640 & ~new_n15137 ;
  assign new_n19325 = new_n15137 & ~new_n16052 ;
  assign new_n19326 = ~new_n19324 & ~new_n19325 ;
  assign new_n19327 = lo0641 & new_n2252 ;
  assign new_n19328 = ~new_n2252 & ~new_n12429 ;
  assign new_n19329 = ~new_n19327 & ~new_n19328 ;
  assign new_n19330 = lo0642 & new_n15454 ;
  assign new_n19331 = lo0958 & ~new_n19223 ;
  assign new_n19332 = lo0642 & ~lo0803 ;
  assign new_n19333 = ~lo0642 & lo0803 ;
  assign new_n19334 = ~new_n19332 & ~new_n19333 ;
  assign new_n19335 = ~lo0958 & ~new_n19334 ;
  assign new_n19336 = ~new_n19331 & ~new_n19335 ;
  assign new_n19337 = ~new_n15454 & ~new_n19336 ;
  assign new_n19338 = ~new_n19330 & ~new_n19337 ;
  assign new_n19339 = lo0643 & ~new_n17223 ;
  assign new_n19340 = new_n17223 & ~new_n19223 ;
  assign new_n19341 = ~new_n19339 & ~new_n19340 ;
  assign new_n19342 = lo0644 & ~new_n15365 ;
  assign new_n19343 = lo0952 & ~new_n19223 ;
  assign new_n19344 = ~lo0952 & new_n6899 ;
  assign new_n19345 = ~new_n19343 & ~new_n19344 ;
  assign new_n19346 = new_n15365 & ~new_n19345 ;
  assign new_n19347 = ~new_n19342 & ~new_n19346 ;
  assign new_n19348 = lo0645 & ~new_n14848 ;
  assign new_n19349 = new_n3806 & ~new_n14853 ;
  assign new_n19350 = ~new_n14181 & new_n14853 ;
  assign new_n19351 = ~new_n19349 & ~new_n19350 ;
  assign new_n19352 = new_n14848 & ~new_n19351 ;
  assign new_n19353 = ~new_n19348 & ~new_n19352 ;
  assign new_n19354 = lo0646 & ~new_n14869 ;
  assign new_n19355 = new_n3806 & ~new_n14872 ;
  assign new_n19356 = ~new_n14181 & new_n14872 ;
  assign new_n19357 = ~new_n19355 & ~new_n19356 ;
  assign new_n19358 = new_n14869 & ~new_n19357 ;
  assign new_n19359 = ~new_n19354 & ~new_n19358 ;
  assign new_n19360 = lo0647 & ~new_n14886 ;
  assign new_n19361 = new_n3806 & ~new_n14889 ;
  assign new_n19362 = ~new_n14181 & new_n14889 ;
  assign new_n19363 = ~new_n19361 & ~new_n19362 ;
  assign new_n19364 = new_n14886 & ~new_n19363 ;
  assign new_n19365 = ~new_n19360 & ~new_n19364 ;
  assign new_n19366 = lo0648 & ~new_n14903 ;
  assign new_n19367 = new_n3806 & ~new_n14906 ;
  assign new_n19368 = ~new_n14181 & new_n14906 ;
  assign new_n19369 = ~new_n19367 & ~new_n19368 ;
  assign new_n19370 = new_n14903 & ~new_n19369 ;
  assign new_n19371 = ~new_n19366 & ~new_n19370 ;
  assign new_n19372 = lo0649 & ~new_n14924 ;
  assign new_n19373 = new_n3806 & ~new_n14927 ;
  assign new_n19374 = ~new_n14181 & new_n14927 ;
  assign new_n19375 = ~new_n19373 & ~new_n19374 ;
  assign new_n19376 = new_n14924 & ~new_n19375 ;
  assign new_n19377 = ~new_n19372 & ~new_n19376 ;
  assign new_n19378 = lo0650 & ~new_n14943 ;
  assign new_n19379 = new_n3806 & ~new_n14946 ;
  assign new_n19380 = ~new_n14181 & new_n14946 ;
  assign new_n19381 = ~new_n19379 & ~new_n19380 ;
  assign new_n19382 = new_n14943 & ~new_n19381 ;
  assign new_n19383 = ~new_n19378 & ~new_n19382 ;
  assign new_n19384 = lo0651 & ~new_n14960 ;
  assign new_n19385 = new_n3806 & ~new_n14963 ;
  assign new_n19386 = ~new_n14181 & new_n14963 ;
  assign new_n19387 = ~new_n19385 & ~new_n19386 ;
  assign new_n19388 = new_n14960 & ~new_n19387 ;
  assign new_n19389 = ~new_n19384 & ~new_n19388 ;
  assign new_n19390 = lo0652 & ~new_n14977 ;
  assign new_n19391 = new_n3806 & ~new_n14980 ;
  assign new_n19392 = ~new_n14181 & new_n14980 ;
  assign new_n19393 = ~new_n19391 & ~new_n19392 ;
  assign new_n19394 = new_n14977 & ~new_n19393 ;
  assign new_n19395 = ~new_n19390 & ~new_n19394 ;
  assign new_n19396 = lo0653 & ~new_n14997 ;
  assign new_n19397 = new_n3806 & ~new_n15000 ;
  assign new_n19398 = ~new_n14181 & new_n15000 ;
  assign new_n19399 = ~new_n19397 & ~new_n19398 ;
  assign new_n19400 = new_n14997 & ~new_n19399 ;
  assign new_n19401 = ~new_n19396 & ~new_n19400 ;
  assign new_n19402 = lo0654 & ~new_n15016 ;
  assign new_n19403 = new_n3806 & ~new_n15019 ;
  assign new_n19404 = ~new_n14181 & new_n15019 ;
  assign new_n19405 = ~new_n19403 & ~new_n19404 ;
  assign new_n19406 = new_n15016 & ~new_n19405 ;
  assign new_n19407 = ~new_n19402 & ~new_n19406 ;
  assign new_n19408 = lo0655 & ~new_n15033 ;
  assign new_n19409 = new_n3806 & ~new_n15036 ;
  assign new_n19410 = ~new_n14181 & new_n15036 ;
  assign new_n19411 = ~new_n19409 & ~new_n19410 ;
  assign new_n19412 = new_n15033 & ~new_n19411 ;
  assign new_n19413 = ~new_n19408 & ~new_n19412 ;
  assign new_n19414 = lo0656 & ~new_n15050 ;
  assign new_n19415 = new_n3806 & ~new_n15053 ;
  assign new_n19416 = ~new_n14181 & new_n15053 ;
  assign new_n19417 = ~new_n19415 & ~new_n19416 ;
  assign new_n19418 = new_n15050 & ~new_n19417 ;
  assign new_n19419 = ~new_n19414 & ~new_n19418 ;
  assign new_n19420 = lo0657 & ~new_n15071 ;
  assign new_n19421 = new_n3806 & ~new_n15074 ;
  assign new_n19422 = ~new_n14181 & new_n15074 ;
  assign new_n19423 = ~new_n19421 & ~new_n19422 ;
  assign new_n19424 = new_n15071 & ~new_n19423 ;
  assign new_n19425 = ~new_n19420 & ~new_n19424 ;
  assign new_n19426 = lo0658 & ~new_n15090 ;
  assign new_n19427 = new_n3806 & ~new_n15093 ;
  assign new_n19428 = ~new_n14181 & new_n15093 ;
  assign new_n19429 = ~new_n19427 & ~new_n19428 ;
  assign new_n19430 = new_n15090 & ~new_n19429 ;
  assign new_n19431 = ~new_n19426 & ~new_n19430 ;
  assign new_n19432 = lo0659 & ~new_n15107 ;
  assign new_n19433 = new_n3806 & ~new_n15110 ;
  assign new_n19434 = ~new_n14181 & new_n15110 ;
  assign new_n19435 = ~new_n19433 & ~new_n19434 ;
  assign new_n19436 = new_n15107 & ~new_n19435 ;
  assign new_n19437 = ~new_n19432 & ~new_n19436 ;
  assign new_n19438 = lo0660 & ~new_n15124 ;
  assign new_n19439 = new_n3806 & ~new_n15127 ;
  assign new_n19440 = ~new_n14181 & new_n15127 ;
  assign new_n19441 = ~new_n19439 & ~new_n19440 ;
  assign new_n19442 = new_n15124 & ~new_n19441 ;
  assign new_n19443 = ~new_n19438 & ~new_n19442 ;
  assign new_n19444 = lo0661 & new_n15454 ;
  assign new_n19445 = lo0958 & ~new_n14181 ;
  assign new_n19446 = ~lo0958 & ~new_n14185 ;
  assign new_n19447 = ~new_n19445 & ~new_n19446 ;
  assign new_n19448 = ~new_n15454 & ~new_n19447 ;
  assign new_n19449 = ~new_n19444 & ~new_n19448 ;
  assign new_n19450 = lo0662 & ~new_n15365 ;
  assign new_n19451 = lo0952 & ~new_n14181 ;
  assign new_n19452 = ~lo0952 & new_n3806 ;
  assign new_n19453 = ~new_n19451 & ~new_n19452 ;
  assign new_n19454 = new_n15365 & ~new_n19453 ;
  assign new_n19455 = ~new_n19450 & ~new_n19454 ;
  assign new_n19456 = lo0663 & ~new_n17223 ;
  assign new_n19457 = ~new_n14181 & new_n17223 ;
  assign new_n19458 = ~new_n19456 & ~new_n19457 ;
  assign new_n19459 = lo0664 & ~new_n14943 ;
  assign new_n19460 = new_n4086 & ~new_n14946 ;
  assign new_n19461 = ~new_n14207 & new_n14946 ;
  assign new_n19462 = ~new_n19460 & ~new_n19461 ;
  assign new_n19463 = new_n14943 & ~new_n19462 ;
  assign new_n19464 = ~new_n19459 & ~new_n19463 ;
  assign new_n19465 = lo0665 & ~new_n14848 ;
  assign new_n19466 = new_n4086 & ~new_n14853 ;
  assign new_n19467 = ~new_n14207 & new_n14853 ;
  assign new_n19468 = ~new_n19466 & ~new_n19467 ;
  assign new_n19469 = new_n14848 & ~new_n19468 ;
  assign new_n19470 = ~new_n19465 & ~new_n19469 ;
  assign new_n19471 = lo0666 & ~new_n14997 ;
  assign new_n19472 = new_n4086 & ~new_n15000 ;
  assign new_n19473 = ~new_n14207 & new_n15000 ;
  assign new_n19474 = ~new_n19472 & ~new_n19473 ;
  assign new_n19475 = new_n14997 & ~new_n19474 ;
  assign new_n19476 = ~new_n19471 & ~new_n19475 ;
  assign new_n19477 = lo0667 & ~new_n15090 ;
  assign new_n19478 = new_n4086 & ~new_n15093 ;
  assign new_n19479 = ~new_n14207 & new_n15093 ;
  assign new_n19480 = ~new_n19478 & ~new_n19479 ;
  assign new_n19481 = new_n15090 & ~new_n19480 ;
  assign new_n19482 = ~new_n19477 & ~new_n19481 ;
  assign new_n19483 = lo0668 & ~new_n14869 ;
  assign new_n19484 = new_n4086 & ~new_n14872 ;
  assign new_n19485 = ~new_n14207 & new_n14872 ;
  assign new_n19486 = ~new_n19484 & ~new_n19485 ;
  assign new_n19487 = new_n14869 & ~new_n19486 ;
  assign new_n19488 = ~new_n19483 & ~new_n19487 ;
  assign new_n19489 = lo0669 & ~new_n14924 ;
  assign new_n19490 = new_n4086 & ~new_n14927 ;
  assign new_n19491 = ~new_n14207 & new_n14927 ;
  assign new_n19492 = ~new_n19490 & ~new_n19491 ;
  assign new_n19493 = new_n14924 & ~new_n19492 ;
  assign new_n19494 = ~new_n19489 & ~new_n19493 ;
  assign new_n19495 = lo0670 & ~new_n15016 ;
  assign new_n19496 = new_n4086 & ~new_n15019 ;
  assign new_n19497 = ~new_n14207 & new_n15019 ;
  assign new_n19498 = ~new_n19496 & ~new_n19497 ;
  assign new_n19499 = new_n15016 & ~new_n19498 ;
  assign new_n19500 = ~new_n19495 & ~new_n19499 ;
  assign new_n19501 = lo0671 & ~new_n15071 ;
  assign new_n19502 = new_n4086 & ~new_n15074 ;
  assign new_n19503 = ~new_n14207 & new_n15074 ;
  assign new_n19504 = ~new_n19502 & ~new_n19503 ;
  assign new_n19505 = new_n15071 & ~new_n19504 ;
  assign new_n19506 = ~new_n19501 & ~new_n19505 ;
  assign new_n19507 = lo0672 & ~new_n14960 ;
  assign new_n19508 = new_n4086 & ~new_n14963 ;
  assign new_n19509 = ~new_n14207 & new_n14963 ;
  assign new_n19510 = ~new_n19508 & ~new_n19509 ;
  assign new_n19511 = new_n14960 & ~new_n19510 ;
  assign new_n19512 = ~new_n19507 & ~new_n19511 ;
  assign new_n19513 = lo0673 & ~new_n14886 ;
  assign new_n19514 = new_n4086 & ~new_n14889 ;
  assign new_n19515 = ~new_n14207 & new_n14889 ;
  assign new_n19516 = ~new_n19514 & ~new_n19515 ;
  assign new_n19517 = new_n14886 & ~new_n19516 ;
  assign new_n19518 = ~new_n19513 & ~new_n19517 ;
  assign new_n19519 = lo0674 & ~new_n15033 ;
  assign new_n19520 = new_n4086 & ~new_n15036 ;
  assign new_n19521 = ~new_n14207 & new_n15036 ;
  assign new_n19522 = ~new_n19520 & ~new_n19521 ;
  assign new_n19523 = new_n15033 & ~new_n19522 ;
  assign new_n19524 = ~new_n19519 & ~new_n19523 ;
  assign new_n19525 = lo0675 & ~new_n15107 ;
  assign new_n19526 = new_n4086 & ~new_n15110 ;
  assign new_n19527 = ~new_n14207 & new_n15110 ;
  assign new_n19528 = ~new_n19526 & ~new_n19527 ;
  assign new_n19529 = new_n15107 & ~new_n19528 ;
  assign new_n19530 = ~new_n19525 & ~new_n19529 ;
  assign new_n19531 = lo0676 & ~new_n14903 ;
  assign new_n19532 = new_n4086 & ~new_n14906 ;
  assign new_n19533 = ~new_n14207 & new_n14906 ;
  assign new_n19534 = ~new_n19532 & ~new_n19533 ;
  assign new_n19535 = new_n14903 & ~new_n19534 ;
  assign new_n19536 = ~new_n19531 & ~new_n19535 ;
  assign new_n19537 = lo0677 & ~new_n14977 ;
  assign new_n19538 = new_n4086 & ~new_n14980 ;
  assign new_n19539 = ~new_n14207 & new_n14980 ;
  assign new_n19540 = ~new_n19538 & ~new_n19539 ;
  assign new_n19541 = new_n14977 & ~new_n19540 ;
  assign new_n19542 = ~new_n19537 & ~new_n19541 ;
  assign new_n19543 = lo0678 & ~new_n15050 ;
  assign new_n19544 = new_n4086 & ~new_n15053 ;
  assign new_n19545 = ~new_n14207 & new_n15053 ;
  assign new_n19546 = ~new_n19544 & ~new_n19545 ;
  assign new_n19547 = new_n15050 & ~new_n19546 ;
  assign new_n19548 = ~new_n19543 & ~new_n19547 ;
  assign new_n19549 = lo0679 & ~new_n15124 ;
  assign new_n19550 = new_n4086 & ~new_n15127 ;
  assign new_n19551 = ~new_n14207 & new_n15127 ;
  assign new_n19552 = ~new_n19550 & ~new_n19551 ;
  assign new_n19553 = new_n15124 & ~new_n19552 ;
  assign new_n19554 = ~new_n19549 & ~new_n19553 ;
  assign new_n19555 = lo0680 & new_n15454 ;
  assign new_n19556 = lo0958 & ~new_n14207 ;
  assign new_n19557 = ~lo0958 & ~new_n14210 ;
  assign new_n19558 = ~new_n19556 & ~new_n19557 ;
  assign new_n19559 = ~new_n15454 & ~new_n19558 ;
  assign new_n19560 = ~new_n19555 & ~new_n19559 ;
  assign new_n19561 = lo0681 & ~new_n15365 ;
  assign new_n19562 = lo0952 & ~new_n14207 ;
  assign new_n19563 = ~lo0952 & new_n4086 ;
  assign new_n19564 = ~new_n19562 & ~new_n19563 ;
  assign new_n19565 = new_n15365 & ~new_n19564 ;
  assign new_n19566 = ~new_n19561 & ~new_n19565 ;
  assign new_n19567 = lo0682 & ~new_n17223 ;
  assign new_n19568 = ~new_n14207 & new_n17223 ;
  assign new_n19569 = ~new_n19567 & ~new_n19568 ;
  assign new_n19570 = lo0683 & ~new_n14943 ;
  assign new_n19571 = ~new_n4889 & ~new_n14946 ;
  assign new_n19572 = ~new_n14525 & new_n14946 ;
  assign new_n19573 = ~new_n19571 & ~new_n19572 ;
  assign new_n19574 = new_n14943 & ~new_n19573 ;
  assign new_n19575 = ~new_n19570 & ~new_n19574 ;
  assign new_n19576 = lo0684 & ~new_n14924 ;
  assign new_n19577 = ~new_n4889 & ~new_n14927 ;
  assign new_n19578 = ~new_n14525 & new_n14927 ;
  assign new_n19579 = ~new_n19577 & ~new_n19578 ;
  assign new_n19580 = new_n14924 & ~new_n19579 ;
  assign new_n19581 = ~new_n19576 & ~new_n19580 ;
  assign new_n19582 = lo0685 & ~new_n14960 ;
  assign new_n19583 = ~new_n4889 & ~new_n14963 ;
  assign new_n19584 = ~new_n14525 & new_n14963 ;
  assign new_n19585 = ~new_n19583 & ~new_n19584 ;
  assign new_n19586 = new_n14960 & ~new_n19585 ;
  assign new_n19587 = ~new_n19582 & ~new_n19586 ;
  assign new_n19588 = lo0686 & ~new_n14977 ;
  assign new_n19589 = ~new_n4889 & ~new_n14980 ;
  assign new_n19590 = ~new_n14525 & new_n14980 ;
  assign new_n19591 = ~new_n19589 & ~new_n19590 ;
  assign new_n19592 = new_n14977 & ~new_n19591 ;
  assign new_n19593 = ~new_n19588 & ~new_n19592 ;
  assign new_n19594 = lo0687 & ~new_n14869 ;
  assign new_n19595 = ~new_n4889 & ~new_n14872 ;
  assign new_n19596 = ~new_n14525 & new_n14872 ;
  assign new_n19597 = ~new_n19595 & ~new_n19596 ;
  assign new_n19598 = new_n14869 & ~new_n19597 ;
  assign new_n19599 = ~new_n19594 & ~new_n19598 ;
  assign new_n19600 = lo0688 & ~new_n14848 ;
  assign new_n19601 = ~new_n4889 & ~new_n14853 ;
  assign new_n19602 = ~new_n14525 & new_n14853 ;
  assign new_n19603 = ~new_n19601 & ~new_n19602 ;
  assign new_n19604 = new_n14848 & ~new_n19603 ;
  assign new_n19605 = ~new_n19600 & ~new_n19604 ;
  assign new_n19606 = lo0689 & ~new_n14886 ;
  assign new_n19607 = ~new_n4889 & ~new_n14889 ;
  assign new_n19608 = ~new_n14525 & new_n14889 ;
  assign new_n19609 = ~new_n19607 & ~new_n19608 ;
  assign new_n19610 = new_n14886 & ~new_n19609 ;
  assign new_n19611 = ~new_n19606 & ~new_n19610 ;
  assign new_n19612 = lo0690 & ~new_n14903 ;
  assign new_n19613 = ~new_n4889 & ~new_n14906 ;
  assign new_n19614 = ~new_n14525 & new_n14906 ;
  assign new_n19615 = ~new_n19613 & ~new_n19614 ;
  assign new_n19616 = new_n14903 & ~new_n19615 ;
  assign new_n19617 = ~new_n19612 & ~new_n19616 ;
  assign new_n19618 = lo0691 & ~new_n15016 ;
  assign new_n19619 = ~new_n4889 & ~new_n15019 ;
  assign new_n19620 = ~new_n14525 & new_n15019 ;
  assign new_n19621 = ~new_n19619 & ~new_n19620 ;
  assign new_n19622 = new_n15016 & ~new_n19621 ;
  assign new_n19623 = ~new_n19618 & ~new_n19622 ;
  assign new_n19624 = lo0692 & ~new_n14997 ;
  assign new_n19625 = ~new_n4889 & ~new_n15000 ;
  assign new_n19626 = ~new_n14525 & new_n15000 ;
  assign new_n19627 = ~new_n19625 & ~new_n19626 ;
  assign new_n19628 = new_n14997 & ~new_n19627 ;
  assign new_n19629 = ~new_n19624 & ~new_n19628 ;
  assign new_n19630 = lo0693 & ~new_n15050 ;
  assign new_n19631 = ~new_n4889 & ~new_n15053 ;
  assign new_n19632 = ~new_n14525 & new_n15053 ;
  assign new_n19633 = ~new_n19631 & ~new_n19632 ;
  assign new_n19634 = new_n15050 & ~new_n19633 ;
  assign new_n19635 = ~new_n19630 & ~new_n19634 ;
  assign new_n19636 = lo0694 & ~new_n15090 ;
  assign new_n19637 = ~new_n4889 & ~new_n15093 ;
  assign new_n19638 = ~new_n14525 & new_n15093 ;
  assign new_n19639 = ~new_n19637 & ~new_n19638 ;
  assign new_n19640 = new_n15090 & ~new_n19639 ;
  assign new_n19641 = ~new_n19636 & ~new_n19640 ;
  assign new_n19642 = lo0695 & ~new_n15071 ;
  assign new_n19643 = ~new_n4889 & ~new_n15074 ;
  assign new_n19644 = ~new_n14525 & new_n15074 ;
  assign new_n19645 = ~new_n19643 & ~new_n19644 ;
  assign new_n19646 = new_n15071 & ~new_n19645 ;
  assign new_n19647 = ~new_n19642 & ~new_n19646 ;
  assign new_n19648 = lo0696 & ~new_n15107 ;
  assign new_n19649 = ~new_n4889 & ~new_n15110 ;
  assign new_n19650 = ~new_n14525 & new_n15110 ;
  assign new_n19651 = ~new_n19649 & ~new_n19650 ;
  assign new_n19652 = new_n15107 & ~new_n19651 ;
  assign new_n19653 = ~new_n19648 & ~new_n19652 ;
  assign new_n19654 = lo0697 & ~new_n15124 ;
  assign new_n19655 = ~new_n4889 & ~new_n15127 ;
  assign new_n19656 = ~new_n14525 & new_n15127 ;
  assign new_n19657 = ~new_n19655 & ~new_n19656 ;
  assign new_n19658 = new_n15124 & ~new_n19657 ;
  assign new_n19659 = ~new_n19654 & ~new_n19658 ;
  assign new_n19660 = lo0698 & new_n2252 ;
  assign new_n19661 = ~new_n2252 & ~new_n2465 ;
  assign new_n19662 = ~new_n19660 & ~new_n19661 ;
  assign new_n19663 = lo0699 & new_n15454 ;
  assign new_n19664 = lo0958 & ~new_n14525 ;
  assign new_n19665 = ~lo0958 & ~new_n14528 ;
  assign new_n19666 = ~new_n19664 & ~new_n19665 ;
  assign new_n19667 = ~new_n15454 & ~new_n19666 ;
  assign new_n19668 = ~new_n19663 & ~new_n19667 ;
  assign new_n19669 = lo0700 & ~new_n17706 ;
  assign new_n19670 = lo0955 & ~new_n14525 ;
  assign new_n19671 = ~lo0955 & ~new_n4889 ;
  assign new_n19672 = ~new_n19670 & ~new_n19671 ;
  assign new_n19673 = new_n17706 & ~new_n19672 ;
  assign new_n19674 = ~new_n19669 & ~new_n19673 ;
  assign new_n19675 = lo0701 & ~new_n17223 ;
  assign new_n19676 = ~new_n14525 & new_n17223 ;
  assign new_n19677 = ~new_n19675 & ~new_n19676 ;
  assign new_n19678 = lo0702 & ~new_n15365 ;
  assign new_n19679 = lo0952 & ~new_n14525 ;
  assign new_n19680 = ~lo0952 & ~new_n4889 ;
  assign new_n19681 = ~new_n19679 & ~new_n19680 ;
  assign new_n19682 = new_n15365 & ~new_n19681 ;
  assign new_n19683 = ~new_n19678 & ~new_n19682 ;
  assign new_n19684 = lo0703 & ~new_n14943 ;
  assign new_n19685 = ~new_n4446 & ~new_n14946 ;
  assign new_n19686 = ~new_n14578 & new_n14946 ;
  assign new_n19687 = ~new_n19685 & ~new_n19686 ;
  assign new_n19688 = new_n14943 & ~new_n19687 ;
  assign new_n19689 = ~new_n19684 & ~new_n19688 ;
  assign new_n19690 = lo0704 & ~new_n14848 ;
  assign new_n19691 = ~new_n4446 & ~new_n14853 ;
  assign new_n19692 = ~new_n14578 & new_n14853 ;
  assign new_n19693 = ~new_n19691 & ~new_n19692 ;
  assign new_n19694 = new_n14848 & ~new_n19693 ;
  assign new_n19695 = ~new_n19690 & ~new_n19694 ;
  assign new_n19696 = lo0705 & ~new_n14997 ;
  assign new_n19697 = ~new_n4446 & ~new_n15000 ;
  assign new_n19698 = ~new_n14578 & new_n15000 ;
  assign new_n19699 = ~new_n19697 & ~new_n19698 ;
  assign new_n19700 = new_n14997 & ~new_n19699 ;
  assign new_n19701 = ~new_n19696 & ~new_n19700 ;
  assign new_n19702 = lo0706 & ~new_n15090 ;
  assign new_n19703 = ~new_n4446 & ~new_n15093 ;
  assign new_n19704 = ~new_n14578 & new_n15093 ;
  assign new_n19705 = ~new_n19703 & ~new_n19704 ;
  assign new_n19706 = new_n15090 & ~new_n19705 ;
  assign new_n19707 = ~new_n19702 & ~new_n19706 ;
  assign new_n19708 = lo0707 & ~new_n14869 ;
  assign new_n19709 = ~new_n4446 & ~new_n14872 ;
  assign new_n19710 = ~new_n14578 & new_n14872 ;
  assign new_n19711 = ~new_n19709 & ~new_n19710 ;
  assign new_n19712 = new_n14869 & ~new_n19711 ;
  assign new_n19713 = ~new_n19708 & ~new_n19712 ;
  assign new_n19714 = lo0708 & ~new_n14924 ;
  assign new_n19715 = ~new_n4446 & ~new_n14927 ;
  assign new_n19716 = ~new_n14578 & new_n14927 ;
  assign new_n19717 = ~new_n19715 & ~new_n19716 ;
  assign new_n19718 = new_n14924 & ~new_n19717 ;
  assign new_n19719 = ~new_n19714 & ~new_n19718 ;
  assign new_n19720 = lo0709 & ~new_n15016 ;
  assign new_n19721 = ~new_n4446 & ~new_n15019 ;
  assign new_n19722 = ~new_n14578 & new_n15019 ;
  assign new_n19723 = ~new_n19721 & ~new_n19722 ;
  assign new_n19724 = new_n15016 & ~new_n19723 ;
  assign new_n19725 = ~new_n19720 & ~new_n19724 ;
  assign new_n19726 = lo0710 & ~new_n15071 ;
  assign new_n19727 = ~new_n4446 & ~new_n15074 ;
  assign new_n19728 = ~new_n14578 & new_n15074 ;
  assign new_n19729 = ~new_n19727 & ~new_n19728 ;
  assign new_n19730 = new_n15071 & ~new_n19729 ;
  assign new_n19731 = ~new_n19726 & ~new_n19730 ;
  assign new_n19732 = lo0711 & ~new_n14960 ;
  assign new_n19733 = ~new_n4446 & ~new_n14963 ;
  assign new_n19734 = ~new_n14578 & new_n14963 ;
  assign new_n19735 = ~new_n19733 & ~new_n19734 ;
  assign new_n19736 = new_n14960 & ~new_n19735 ;
  assign new_n19737 = ~new_n19732 & ~new_n19736 ;
  assign new_n19738 = lo0712 & ~new_n14886 ;
  assign new_n19739 = ~new_n4446 & ~new_n14889 ;
  assign new_n19740 = ~new_n14578 & new_n14889 ;
  assign new_n19741 = ~new_n19739 & ~new_n19740 ;
  assign new_n19742 = new_n14886 & ~new_n19741 ;
  assign new_n19743 = ~new_n19738 & ~new_n19742 ;
  assign new_n19744 = lo0713 & ~new_n15033 ;
  assign new_n19745 = ~new_n4446 & ~new_n15036 ;
  assign new_n19746 = ~new_n14578 & new_n15036 ;
  assign new_n19747 = ~new_n19745 & ~new_n19746 ;
  assign new_n19748 = new_n15033 & ~new_n19747 ;
  assign new_n19749 = ~new_n19744 & ~new_n19748 ;
  assign new_n19750 = lo0714 & ~new_n15107 ;
  assign new_n19751 = ~new_n4446 & ~new_n15110 ;
  assign new_n19752 = ~new_n14578 & new_n15110 ;
  assign new_n19753 = ~new_n19751 & ~new_n19752 ;
  assign new_n19754 = new_n15107 & ~new_n19753 ;
  assign new_n19755 = ~new_n19750 & ~new_n19754 ;
  assign new_n19756 = lo0715 & ~new_n14903 ;
  assign new_n19757 = ~new_n4446 & ~new_n14906 ;
  assign new_n19758 = ~new_n14578 & new_n14906 ;
  assign new_n19759 = ~new_n19757 & ~new_n19758 ;
  assign new_n19760 = new_n14903 & ~new_n19759 ;
  assign new_n19761 = ~new_n19756 & ~new_n19760 ;
  assign new_n19762 = lo0716 & ~new_n14977 ;
  assign new_n19763 = ~new_n4446 & ~new_n14980 ;
  assign new_n19764 = ~new_n14578 & new_n14980 ;
  assign new_n19765 = ~new_n19763 & ~new_n19764 ;
  assign new_n19766 = new_n14977 & ~new_n19765 ;
  assign new_n19767 = ~new_n19762 & ~new_n19766 ;
  assign new_n19768 = lo0717 & ~new_n15050 ;
  assign new_n19769 = ~new_n4446 & ~new_n15053 ;
  assign new_n19770 = ~new_n14578 & new_n15053 ;
  assign new_n19771 = ~new_n19769 & ~new_n19770 ;
  assign new_n19772 = new_n15050 & ~new_n19771 ;
  assign new_n19773 = ~new_n19768 & ~new_n19772 ;
  assign new_n19774 = lo0718 & ~new_n15124 ;
  assign new_n19775 = ~new_n4446 & ~new_n15127 ;
  assign new_n19776 = ~new_n14578 & new_n15127 ;
  assign new_n19777 = ~new_n19775 & ~new_n19776 ;
  assign new_n19778 = new_n15124 & ~new_n19777 ;
  assign new_n19779 = ~new_n19774 & ~new_n19778 ;
  assign new_n19780 = lo0719 & new_n2252 ;
  assign new_n19781 = ~new_n2252 & ~new_n12325 ;
  assign new_n19782 = ~new_n19780 & ~new_n19781 ;
  assign new_n19783 = lo0720 & new_n15454 ;
  assign new_n19784 = lo0958 & ~new_n14578 ;
  assign new_n19785 = ~lo0958 & ~new_n14581 ;
  assign new_n19786 = ~new_n19784 & ~new_n19785 ;
  assign new_n19787 = ~new_n15454 & ~new_n19786 ;
  assign new_n19788 = ~new_n19783 & ~new_n19787 ;
  assign new_n19789 = lo0721 & ~new_n17223 ;
  assign new_n19790 = ~new_n14578 & new_n17223 ;
  assign new_n19791 = ~new_n19789 & ~new_n19790 ;
  assign new_n19792 = lo0722 & ~new_n15365 ;
  assign new_n19793 = lo0952 & ~new_n14578 ;
  assign new_n19794 = ~lo0952 & ~new_n4446 ;
  assign new_n19795 = ~new_n19793 & ~new_n19794 ;
  assign new_n19796 = new_n15365 & ~new_n19795 ;
  assign new_n19797 = ~new_n19792 & ~new_n19796 ;
  assign new_n19798 = lo0723 & ~new_n14924 ;
  assign new_n19799 = new_n4807 & ~new_n14927 ;
  assign new_n19800 = ~new_n14260 & new_n14927 ;
  assign new_n19801 = ~new_n19799 & ~new_n19800 ;
  assign new_n19802 = new_n14924 & ~new_n19801 ;
  assign new_n19803 = ~new_n19798 & ~new_n19802 ;
  assign new_n19804 = lo0724 & ~new_n14869 ;
  assign new_n19805 = new_n4807 & ~new_n14872 ;
  assign new_n19806 = ~new_n14260 & new_n14872 ;
  assign new_n19807 = ~new_n19805 & ~new_n19806 ;
  assign new_n19808 = new_n14869 & ~new_n19807 ;
  assign new_n19809 = ~new_n19804 & ~new_n19808 ;
  assign new_n19810 = lo0725 & ~new_n15016 ;
  assign new_n19811 = new_n4807 & ~new_n15019 ;
  assign new_n19812 = ~new_n14260 & new_n15019 ;
  assign new_n19813 = ~new_n19811 & ~new_n19812 ;
  assign new_n19814 = new_n15016 & ~new_n19813 ;
  assign new_n19815 = ~new_n19810 & ~new_n19814 ;
  assign new_n19816 = lo0726 & ~new_n15071 ;
  assign new_n19817 = new_n4807 & ~new_n15074 ;
  assign new_n19818 = ~new_n14260 & new_n15074 ;
  assign new_n19819 = ~new_n19817 & ~new_n19818 ;
  assign new_n19820 = new_n15071 & ~new_n19819 ;
  assign new_n19821 = ~new_n19816 & ~new_n19820 ;
  assign new_n19822 = lo0727 & ~new_n14848 ;
  assign new_n19823 = new_n4807 & ~new_n14853 ;
  assign new_n19824 = ~new_n14260 & new_n14853 ;
  assign new_n19825 = ~new_n19823 & ~new_n19824 ;
  assign new_n19826 = new_n14848 & ~new_n19825 ;
  assign new_n19827 = ~new_n19822 & ~new_n19826 ;
  assign new_n19828 = lo0728 & ~new_n14943 ;
  assign new_n19829 = new_n4807 & ~new_n14946 ;
  assign new_n19830 = ~new_n14260 & new_n14946 ;
  assign new_n19831 = ~new_n19829 & ~new_n19830 ;
  assign new_n19832 = new_n14943 & ~new_n19831 ;
  assign new_n19833 = ~new_n19828 & ~new_n19832 ;
  assign new_n19834 = lo0729 & ~new_n14997 ;
  assign new_n19835 = new_n4807 & ~new_n15000 ;
  assign new_n19836 = ~new_n14260 & new_n15000 ;
  assign new_n19837 = ~new_n19835 & ~new_n19836 ;
  assign new_n19838 = new_n14997 & ~new_n19837 ;
  assign new_n19839 = ~new_n19834 & ~new_n19838 ;
  assign new_n19840 = lo0730 & ~new_n15090 ;
  assign new_n19841 = new_n4807 & ~new_n15093 ;
  assign new_n19842 = ~new_n14260 & new_n15093 ;
  assign new_n19843 = ~new_n19841 & ~new_n19842 ;
  assign new_n19844 = new_n15090 & ~new_n19843 ;
  assign new_n19845 = ~new_n19840 & ~new_n19844 ;
  assign new_n19846 = lo0731 & ~new_n14886 ;
  assign new_n19847 = new_n4807 & ~new_n14889 ;
  assign new_n19848 = ~new_n14260 & new_n14889 ;
  assign new_n19849 = ~new_n19847 & ~new_n19848 ;
  assign new_n19850 = new_n14886 & ~new_n19849 ;
  assign new_n19851 = ~new_n19846 & ~new_n19850 ;
  assign new_n19852 = lo0732 & ~new_n14960 ;
  assign new_n19853 = new_n4807 & ~new_n14963 ;
  assign new_n19854 = ~new_n14260 & new_n14963 ;
  assign new_n19855 = ~new_n19853 & ~new_n19854 ;
  assign new_n19856 = new_n14960 & ~new_n19855 ;
  assign new_n19857 = ~new_n19852 & ~new_n19856 ;
  assign new_n19858 = lo0733 & ~new_n15033 ;
  assign new_n19859 = new_n4807 & ~new_n15036 ;
  assign new_n19860 = ~new_n14260 & new_n15036 ;
  assign new_n19861 = ~new_n19859 & ~new_n19860 ;
  assign new_n19862 = new_n15033 & ~new_n19861 ;
  assign new_n19863 = ~new_n19858 & ~new_n19862 ;
  assign new_n19864 = lo0734 & ~new_n15107 ;
  assign new_n19865 = new_n4807 & ~new_n15110 ;
  assign new_n19866 = ~new_n14260 & new_n15110 ;
  assign new_n19867 = ~new_n19865 & ~new_n19866 ;
  assign new_n19868 = new_n15107 & ~new_n19867 ;
  assign new_n19869 = ~new_n19864 & ~new_n19868 ;
  assign new_n19870 = lo0735 & ~new_n14977 ;
  assign new_n19871 = new_n4807 & ~new_n14980 ;
  assign new_n19872 = ~new_n14260 & new_n14980 ;
  assign new_n19873 = ~new_n19871 & ~new_n19872 ;
  assign new_n19874 = new_n14977 & ~new_n19873 ;
  assign new_n19875 = ~new_n19870 & ~new_n19874 ;
  assign new_n19876 = lo0736 & ~new_n14903 ;
  assign new_n19877 = new_n4807 & ~new_n14906 ;
  assign new_n19878 = ~new_n14260 & new_n14906 ;
  assign new_n19879 = ~new_n19877 & ~new_n19878 ;
  assign new_n19880 = new_n14903 & ~new_n19879 ;
  assign new_n19881 = ~new_n19876 & ~new_n19880 ;
  assign new_n19882 = lo0737 & ~new_n15050 ;
  assign new_n19883 = new_n4807 & ~new_n15053 ;
  assign new_n19884 = ~new_n14260 & new_n15053 ;
  assign new_n19885 = ~new_n19883 & ~new_n19884 ;
  assign new_n19886 = new_n15050 & ~new_n19885 ;
  assign new_n19887 = ~new_n19882 & ~new_n19886 ;
  assign new_n19888 = lo0738 & ~new_n15124 ;
  assign new_n19889 = new_n4807 & ~new_n15127 ;
  assign new_n19890 = ~new_n14260 & new_n15127 ;
  assign new_n19891 = ~new_n19889 & ~new_n19890 ;
  assign new_n19892 = new_n15124 & ~new_n19891 ;
  assign new_n19893 = ~new_n19888 & ~new_n19892 ;
  assign new_n19894 = lo0739 & new_n15454 ;
  assign new_n19895 = lo0958 & ~new_n14260 ;
  assign new_n19896 = ~lo0958 & ~new_n14263 ;
  assign new_n19897 = ~new_n19895 & ~new_n19896 ;
  assign new_n19898 = ~new_n15454 & ~new_n19897 ;
  assign new_n19899 = ~new_n19894 & ~new_n19898 ;
  assign new_n19900 = lo0740 & ~new_n15365 ;
  assign new_n19901 = lo0952 & ~new_n14260 ;
  assign new_n19902 = ~lo0952 & new_n4807 ;
  assign new_n19903 = ~new_n19901 & ~new_n19902 ;
  assign new_n19904 = new_n15365 & ~new_n19903 ;
  assign new_n19905 = ~new_n19900 & ~new_n19904 ;
  assign new_n19906 = lo0741 & ~new_n17223 ;
  assign new_n19907 = ~new_n14260 & new_n17223 ;
  assign new_n19908 = ~new_n19906 & ~new_n19907 ;
  assign new_n19909 = lo0742 & ~new_n15033 ;
  assign new_n19910 = new_n2586 & ~new_n15036 ;
  assign new_n19911 = ~new_n10308 & new_n15036 ;
  assign new_n19912 = ~new_n19910 & ~new_n19911 ;
  assign new_n19913 = new_n15033 & ~new_n19912 ;
  assign new_n19914 = ~new_n19909 & ~new_n19913 ;
  assign new_n19915 = lo0743 & ~new_n14848 ;
  assign new_n19916 = new_n2586 & ~new_n14853 ;
  assign new_n19917 = ~new_n10308 & new_n14853 ;
  assign new_n19918 = ~new_n19916 & ~new_n19917 ;
  assign new_n19919 = new_n14848 & ~new_n19918 ;
  assign new_n19920 = ~new_n19915 & ~new_n19919 ;
  assign new_n19921 = lo0744 & ~new_n14869 ;
  assign new_n19922 = new_n2586 & ~new_n14872 ;
  assign new_n19923 = ~new_n10308 & new_n14872 ;
  assign new_n19924 = ~new_n19922 & ~new_n19923 ;
  assign new_n19925 = new_n14869 & ~new_n19924 ;
  assign new_n19926 = ~new_n19921 & ~new_n19925 ;
  assign new_n19927 = lo0745 & ~new_n14886 ;
  assign new_n19928 = new_n2586 & ~new_n14889 ;
  assign new_n19929 = ~new_n10308 & new_n14889 ;
  assign new_n19930 = ~new_n19928 & ~new_n19929 ;
  assign new_n19931 = new_n14886 & ~new_n19930 ;
  assign new_n19932 = ~new_n19927 & ~new_n19931 ;
  assign new_n19933 = lo0746 & ~new_n14903 ;
  assign new_n19934 = new_n2586 & ~new_n14906 ;
  assign new_n19935 = ~new_n10308 & new_n14906 ;
  assign new_n19936 = ~new_n19934 & ~new_n19935 ;
  assign new_n19937 = new_n14903 & ~new_n19936 ;
  assign new_n19938 = ~new_n19933 & ~new_n19937 ;
  assign new_n19939 = lo0747 & ~new_n14924 ;
  assign new_n19940 = new_n2586 & ~new_n14927 ;
  assign new_n19941 = ~new_n10308 & new_n14927 ;
  assign new_n19942 = ~new_n19940 & ~new_n19941 ;
  assign new_n19943 = new_n14924 & ~new_n19942 ;
  assign new_n19944 = ~new_n19939 & ~new_n19943 ;
  assign new_n19945 = lo0748 & ~new_n14943 ;
  assign new_n19946 = new_n2586 & ~new_n14946 ;
  assign new_n19947 = ~new_n10308 & new_n14946 ;
  assign new_n19948 = ~new_n19946 & ~new_n19947 ;
  assign new_n19949 = new_n14943 & ~new_n19948 ;
  assign new_n19950 = ~new_n19945 & ~new_n19949 ;
  assign new_n19951 = lo0749 & ~new_n14960 ;
  assign new_n19952 = new_n2586 & ~new_n14963 ;
  assign new_n19953 = ~new_n10308 & new_n14963 ;
  assign new_n19954 = ~new_n19952 & ~new_n19953 ;
  assign new_n19955 = new_n14960 & ~new_n19954 ;
  assign new_n19956 = ~new_n19951 & ~new_n19955 ;
  assign new_n19957 = lo0750 & ~new_n14977 ;
  assign new_n19958 = new_n2586 & ~new_n14980 ;
  assign new_n19959 = ~new_n10308 & new_n14980 ;
  assign new_n19960 = ~new_n19958 & ~new_n19959 ;
  assign new_n19961 = new_n14977 & ~new_n19960 ;
  assign new_n19962 = ~new_n19957 & ~new_n19961 ;
  assign new_n19963 = lo0751 & ~new_n14997 ;
  assign new_n19964 = new_n2586 & ~new_n15000 ;
  assign new_n19965 = ~new_n10308 & new_n15000 ;
  assign new_n19966 = ~new_n19964 & ~new_n19965 ;
  assign new_n19967 = new_n14997 & ~new_n19966 ;
  assign new_n19968 = ~new_n19963 & ~new_n19967 ;
  assign new_n19969 = lo0752 & ~new_n15016 ;
  assign new_n19970 = new_n2586 & ~new_n15019 ;
  assign new_n19971 = ~new_n10308 & new_n15019 ;
  assign new_n19972 = ~new_n19970 & ~new_n19971 ;
  assign new_n19973 = new_n15016 & ~new_n19972 ;
  assign new_n19974 = ~new_n19969 & ~new_n19973 ;
  assign new_n19975 = lo0753 & ~new_n15050 ;
  assign new_n19976 = new_n2586 & ~new_n15053 ;
  assign new_n19977 = ~new_n10308 & new_n15053 ;
  assign new_n19978 = ~new_n19976 & ~new_n19977 ;
  assign new_n19979 = new_n15050 & ~new_n19978 ;
  assign new_n19980 = ~new_n19975 & ~new_n19979 ;
  assign new_n19981 = lo0754 & ~new_n15071 ;
  assign new_n19982 = new_n2586 & ~new_n15074 ;
  assign new_n19983 = ~new_n10308 & new_n15074 ;
  assign new_n19984 = ~new_n19982 & ~new_n19983 ;
  assign new_n19985 = new_n15071 & ~new_n19984 ;
  assign new_n19986 = ~new_n19981 & ~new_n19985 ;
  assign new_n19987 = lo0755 & ~new_n15090 ;
  assign new_n19988 = new_n2586 & ~new_n15093 ;
  assign new_n19989 = ~new_n10308 & new_n15093 ;
  assign new_n19990 = ~new_n19988 & ~new_n19989 ;
  assign new_n19991 = new_n15090 & ~new_n19990 ;
  assign new_n19992 = ~new_n19987 & ~new_n19991 ;
  assign new_n19993 = lo0756 & ~new_n15107 ;
  assign new_n19994 = new_n2586 & ~new_n15110 ;
  assign new_n19995 = ~new_n10308 & new_n15110 ;
  assign new_n19996 = ~new_n19994 & ~new_n19995 ;
  assign new_n19997 = new_n15107 & ~new_n19996 ;
  assign new_n19998 = ~new_n19993 & ~new_n19997 ;
  assign new_n19999 = lo0757 & ~new_n15124 ;
  assign new_n20000 = new_n2586 & ~new_n15127 ;
  assign new_n20001 = ~new_n10308 & new_n15127 ;
  assign new_n20002 = ~new_n20000 & ~new_n20001 ;
  assign new_n20003 = new_n15124 & ~new_n20002 ;
  assign new_n20004 = ~new_n19999 & ~new_n20003 ;
  assign new_n20005 = lo0758 & ~new_n15137 ;
  assign new_n20006 = new_n15137 & ~new_n16443 ;
  assign new_n20007 = ~new_n20005 & ~new_n20006 ;
  assign new_n20008 = ~new_n10308 & new_n15393 ;
  assign new_n20009 = lo0759 & ~new_n15393 ;
  assign new_n20010 = ~new_n20008 & ~new_n20009 ;
  assign new_n20011 = lo0760 & ~new_n15376 ;
  assign new_n20012 = ~new_n12313 & new_n15376 ;
  assign new_n20013 = ~new_n20011 & ~new_n20012 ;
  assign new_n20014 = lo0761 & ~new_n15365 ;
  assign new_n20015 = lo0952 & ~new_n10308 ;
  assign new_n20016 = ~lo0952 & new_n2586 ;
  assign new_n20017 = ~new_n20015 & ~new_n20016 ;
  assign new_n20018 = new_n15365 & ~new_n20017 ;
  assign new_n20019 = ~new_n20014 & ~new_n20018 ;
  assign new_n20020 = lo0762 & ~new_n17223 ;
  assign new_n20021 = ~new_n10308 & new_n17223 ;
  assign new_n20022 = ~new_n20020 & ~new_n20021 ;
  assign new_n20023 = lo0763 & ~new_n17223 ;
  assign new_n20024 = ~new_n13936 & new_n17223 ;
  assign new_n20025 = ~new_n20023 & ~new_n20024 ;
  assign new_n20026 = lo0764 & ~new_n14943 ;
  assign new_n20027 = new_n5265 & ~new_n14946 ;
  assign new_n20028 = ~new_n14446 & new_n14946 ;
  assign new_n20029 = ~new_n20027 & ~new_n20028 ;
  assign new_n20030 = new_n14943 & ~new_n20029 ;
  assign new_n20031 = ~new_n20026 & ~new_n20030 ;
  assign new_n20032 = lo0765 & ~new_n14924 ;
  assign new_n20033 = new_n5265 & ~new_n14927 ;
  assign new_n20034 = ~new_n14446 & new_n14927 ;
  assign new_n20035 = ~new_n20033 & ~new_n20034 ;
  assign new_n20036 = new_n14924 & ~new_n20035 ;
  assign new_n20037 = ~new_n20032 & ~new_n20036 ;
  assign new_n20038 = lo0766 & ~new_n14960 ;
  assign new_n20039 = new_n5265 & ~new_n14963 ;
  assign new_n20040 = ~new_n14446 & new_n14963 ;
  assign new_n20041 = ~new_n20039 & ~new_n20040 ;
  assign new_n20042 = new_n14960 & ~new_n20041 ;
  assign new_n20043 = ~new_n20038 & ~new_n20042 ;
  assign new_n20044 = lo0767 & ~new_n14977 ;
  assign new_n20045 = new_n5265 & ~new_n14980 ;
  assign new_n20046 = ~new_n14446 & new_n14980 ;
  assign new_n20047 = ~new_n20045 & ~new_n20046 ;
  assign new_n20048 = new_n14977 & ~new_n20047 ;
  assign new_n20049 = ~new_n20044 & ~new_n20048 ;
  assign new_n20050 = lo0768 & ~new_n14869 ;
  assign new_n20051 = new_n5265 & ~new_n14872 ;
  assign new_n20052 = ~new_n14446 & new_n14872 ;
  assign new_n20053 = ~new_n20051 & ~new_n20052 ;
  assign new_n20054 = new_n14869 & ~new_n20053 ;
  assign new_n20055 = ~new_n20050 & ~new_n20054 ;
  assign new_n20056 = lo0769 & ~new_n14848 ;
  assign new_n20057 = new_n5265 & ~new_n14853 ;
  assign new_n20058 = ~new_n14446 & new_n14853 ;
  assign new_n20059 = ~new_n20057 & ~new_n20058 ;
  assign new_n20060 = new_n14848 & ~new_n20059 ;
  assign new_n20061 = ~new_n20056 & ~new_n20060 ;
  assign new_n20062 = lo0770 & ~new_n14886 ;
  assign new_n20063 = new_n5265 & ~new_n14889 ;
  assign new_n20064 = ~new_n14446 & new_n14889 ;
  assign new_n20065 = ~new_n20063 & ~new_n20064 ;
  assign new_n20066 = new_n14886 & ~new_n20065 ;
  assign new_n20067 = ~new_n20062 & ~new_n20066 ;
  assign new_n20068 = lo0771 & ~new_n14903 ;
  assign new_n20069 = new_n5265 & ~new_n14906 ;
  assign new_n20070 = ~new_n14446 & new_n14906 ;
  assign new_n20071 = ~new_n20069 & ~new_n20070 ;
  assign new_n20072 = new_n14903 & ~new_n20071 ;
  assign new_n20073 = ~new_n20068 & ~new_n20072 ;
  assign new_n20074 = lo0772 & ~new_n15016 ;
  assign new_n20075 = new_n5265 & ~new_n15019 ;
  assign new_n20076 = ~new_n14446 & new_n15019 ;
  assign new_n20077 = ~new_n20075 & ~new_n20076 ;
  assign new_n20078 = new_n15016 & ~new_n20077 ;
  assign new_n20079 = ~new_n20074 & ~new_n20078 ;
  assign new_n20080 = lo0773 & ~new_n14997 ;
  assign new_n20081 = new_n5265 & ~new_n15000 ;
  assign new_n20082 = ~new_n14446 & new_n15000 ;
  assign new_n20083 = ~new_n20081 & ~new_n20082 ;
  assign new_n20084 = new_n14997 & ~new_n20083 ;
  assign new_n20085 = ~new_n20080 & ~new_n20084 ;
  assign new_n20086 = lo0774 & ~new_n15033 ;
  assign new_n20087 = new_n5265 & ~new_n15036 ;
  assign new_n20088 = ~new_n14446 & new_n15036 ;
  assign new_n20089 = ~new_n20087 & ~new_n20088 ;
  assign new_n20090 = new_n15033 & ~new_n20089 ;
  assign new_n20091 = ~new_n20086 & ~new_n20090 ;
  assign new_n20092 = lo0775 & ~new_n15050 ;
  assign new_n20093 = new_n5265 & ~new_n15053 ;
  assign new_n20094 = ~new_n14446 & new_n15053 ;
  assign new_n20095 = ~new_n20093 & ~new_n20094 ;
  assign new_n20096 = new_n15050 & ~new_n20095 ;
  assign new_n20097 = ~new_n20092 & ~new_n20096 ;
  assign new_n20098 = lo0776 & ~new_n15090 ;
  assign new_n20099 = new_n5265 & ~new_n15093 ;
  assign new_n20100 = ~new_n14446 & new_n15093 ;
  assign new_n20101 = ~new_n20099 & ~new_n20100 ;
  assign new_n20102 = new_n15090 & ~new_n20101 ;
  assign new_n20103 = ~new_n20098 & ~new_n20102 ;
  assign new_n20104 = lo0777 & ~new_n15071 ;
  assign new_n20105 = new_n5265 & ~new_n15074 ;
  assign new_n20106 = ~new_n14446 & new_n15074 ;
  assign new_n20107 = ~new_n20105 & ~new_n20106 ;
  assign new_n20108 = new_n15071 & ~new_n20107 ;
  assign new_n20109 = ~new_n20104 & ~new_n20108 ;
  assign new_n20110 = lo0778 & ~new_n15107 ;
  assign new_n20111 = new_n5265 & ~new_n15110 ;
  assign new_n20112 = ~new_n14446 & new_n15110 ;
  assign new_n20113 = ~new_n20111 & ~new_n20112 ;
  assign new_n20114 = new_n15107 & ~new_n20113 ;
  assign new_n20115 = ~new_n20110 & ~new_n20114 ;
  assign new_n20116 = lo0779 & ~new_n15124 ;
  assign new_n20117 = new_n5265 & ~new_n15127 ;
  assign new_n20118 = ~new_n14446 & new_n15127 ;
  assign new_n20119 = ~new_n20117 & ~new_n20118 ;
  assign new_n20120 = new_n15124 & ~new_n20119 ;
  assign new_n20121 = ~new_n20116 & ~new_n20120 ;
  assign new_n20122 = lo0780 & ~new_n15137 ;
  assign new_n20123 = new_n15137 & ~new_n16326 ;
  assign new_n20124 = ~new_n20122 & ~new_n20123 ;
  assign new_n20125 = lo0781 & new_n15454 ;
  assign new_n20126 = lo0958 & ~new_n14446 ;
  assign new_n20127 = ~lo0958 & ~new_n14450 ;
  assign new_n20128 = ~new_n20126 & ~new_n20127 ;
  assign new_n20129 = ~new_n15454 & ~new_n20128 ;
  assign new_n20130 = ~new_n20125 & ~new_n20129 ;
  assign new_n20131 = lo0782 & ~new_n15365 ;
  assign new_n20132 = lo0952 & ~new_n14446 ;
  assign new_n20133 = ~lo0952 & new_n5265 ;
  assign new_n20134 = ~new_n20132 & ~new_n20133 ;
  assign new_n20135 = new_n15365 & ~new_n20134 ;
  assign new_n20136 = ~new_n20131 & ~new_n20135 ;
  assign new_n20137 = lo0783 & ~new_n17223 ;
  assign new_n20138 = ~new_n14446 & new_n17223 ;
  assign new_n20139 = ~new_n20137 & ~new_n20138 ;
  assign new_n20140 = lo0784 & ~new_n14924 ;
  assign new_n20141 = new_n7122 & ~new_n14927 ;
  assign new_n20142 = ~new_n13907 & new_n14927 ;
  assign new_n20143 = ~new_n20141 & ~new_n20142 ;
  assign new_n20144 = new_n14924 & ~new_n20143 ;
  assign new_n20145 = ~new_n20140 & ~new_n20144 ;
  assign new_n20146 = lo0785 & ~new_n14869 ;
  assign new_n20147 = new_n7122 & ~new_n14872 ;
  assign new_n20148 = ~new_n13907 & new_n14872 ;
  assign new_n20149 = ~new_n20147 & ~new_n20148 ;
  assign new_n20150 = new_n14869 & ~new_n20149 ;
  assign new_n20151 = ~new_n20146 & ~new_n20150 ;
  assign new_n20152 = lo0786 & ~new_n15016 ;
  assign new_n20153 = new_n7122 & ~new_n15019 ;
  assign new_n20154 = ~new_n13907 & new_n15019 ;
  assign new_n20155 = ~new_n20153 & ~new_n20154 ;
  assign new_n20156 = new_n15016 & ~new_n20155 ;
  assign new_n20157 = ~new_n20152 & ~new_n20156 ;
  assign new_n20158 = lo0787 & ~new_n15071 ;
  assign new_n20159 = new_n7122 & ~new_n15074 ;
  assign new_n20160 = ~new_n13907 & new_n15074 ;
  assign new_n20161 = ~new_n20159 & ~new_n20160 ;
  assign new_n20162 = new_n15071 & ~new_n20161 ;
  assign new_n20163 = ~new_n20158 & ~new_n20162 ;
  assign new_n20164 = lo0788 & ~new_n14848 ;
  assign new_n20165 = new_n7122 & ~new_n14853 ;
  assign new_n20166 = ~new_n13907 & new_n14853 ;
  assign new_n20167 = ~new_n20165 & ~new_n20166 ;
  assign new_n20168 = new_n14848 & ~new_n20167 ;
  assign new_n20169 = ~new_n20164 & ~new_n20168 ;
  assign new_n20170 = lo0789 & ~new_n14943 ;
  assign new_n20171 = new_n7122 & ~new_n14946 ;
  assign new_n20172 = ~new_n13907 & new_n14946 ;
  assign new_n20173 = ~new_n20171 & ~new_n20172 ;
  assign new_n20174 = new_n14943 & ~new_n20173 ;
  assign new_n20175 = ~new_n20170 & ~new_n20174 ;
  assign new_n20176 = lo0790 & ~new_n14997 ;
  assign new_n20177 = new_n7122 & ~new_n15000 ;
  assign new_n20178 = ~new_n13907 & new_n15000 ;
  assign new_n20179 = ~new_n20177 & ~new_n20178 ;
  assign new_n20180 = new_n14997 & ~new_n20179 ;
  assign new_n20181 = ~new_n20176 & ~new_n20180 ;
  assign new_n20182 = lo0791 & ~new_n15090 ;
  assign new_n20183 = new_n7122 & ~new_n15093 ;
  assign new_n20184 = ~new_n13907 & new_n15093 ;
  assign new_n20185 = ~new_n20183 & ~new_n20184 ;
  assign new_n20186 = new_n15090 & ~new_n20185 ;
  assign new_n20187 = ~new_n20182 & ~new_n20186 ;
  assign new_n20188 = lo0792 & ~new_n14886 ;
  assign new_n20189 = new_n7122 & ~new_n14889 ;
  assign new_n20190 = ~new_n13907 & new_n14889 ;
  assign new_n20191 = ~new_n20189 & ~new_n20190 ;
  assign new_n20192 = new_n14886 & ~new_n20191 ;
  assign new_n20193 = ~new_n20188 & ~new_n20192 ;
  assign new_n20194 = lo0793 & ~new_n14960 ;
  assign new_n20195 = new_n7122 & ~new_n14963 ;
  assign new_n20196 = ~new_n13907 & new_n14963 ;
  assign new_n20197 = ~new_n20195 & ~new_n20196 ;
  assign new_n20198 = new_n14960 & ~new_n20197 ;
  assign new_n20199 = ~new_n20194 & ~new_n20198 ;
  assign new_n20200 = lo0794 & ~new_n15033 ;
  assign new_n20201 = new_n7122 & ~new_n15036 ;
  assign new_n20202 = ~new_n13907 & new_n15036 ;
  assign new_n20203 = ~new_n20201 & ~new_n20202 ;
  assign new_n20204 = new_n15033 & ~new_n20203 ;
  assign new_n20205 = ~new_n20200 & ~new_n20204 ;
  assign new_n20206 = lo0795 & ~new_n15107 ;
  assign new_n20207 = new_n7122 & ~new_n15110 ;
  assign new_n20208 = ~new_n13907 & new_n15110 ;
  assign new_n20209 = ~new_n20207 & ~new_n20208 ;
  assign new_n20210 = new_n15107 & ~new_n20209 ;
  assign new_n20211 = ~new_n20206 & ~new_n20210 ;
  assign new_n20212 = lo0796 & ~new_n14977 ;
  assign new_n20213 = new_n7122 & ~new_n14980 ;
  assign new_n20214 = ~new_n13907 & new_n14980 ;
  assign new_n20215 = ~new_n20213 & ~new_n20214 ;
  assign new_n20216 = new_n14977 & ~new_n20215 ;
  assign new_n20217 = ~new_n20212 & ~new_n20216 ;
  assign new_n20218 = lo0797 & ~new_n14903 ;
  assign new_n20219 = new_n7122 & ~new_n14906 ;
  assign new_n20220 = ~new_n13907 & new_n14906 ;
  assign new_n20221 = ~new_n20219 & ~new_n20220 ;
  assign new_n20222 = new_n14903 & ~new_n20221 ;
  assign new_n20223 = ~new_n20218 & ~new_n20222 ;
  assign new_n20224 = lo0798 & ~new_n15050 ;
  assign new_n20225 = new_n7122 & ~new_n15053 ;
  assign new_n20226 = ~new_n13907 & new_n15053 ;
  assign new_n20227 = ~new_n20225 & ~new_n20226 ;
  assign new_n20228 = new_n15050 & ~new_n20227 ;
  assign new_n20229 = ~new_n20224 & ~new_n20228 ;
  assign new_n20230 = lo0799 & ~new_n15124 ;
  assign new_n20231 = new_n7122 & ~new_n15127 ;
  assign new_n20232 = ~new_n13907 & new_n15127 ;
  assign new_n20233 = ~new_n20231 & ~new_n20232 ;
  assign new_n20234 = new_n15124 & ~new_n20233 ;
  assign new_n20235 = ~new_n20230 & ~new_n20234 ;
  assign new_n20236 = lo0800 & ~new_n15137 ;
  assign new_n20237 = new_n15137 & ~new_n15832 ;
  assign new_n20238 = ~new_n20236 & ~new_n20237 ;
  assign new_n20239 = lo0801 & ~new_n15137 ;
  assign new_n20240 = new_n15137 & ~new_n15807 ;
  assign new_n20241 = ~new_n20239 & ~new_n20240 ;
  assign new_n20242 = lo0802 & ~new_n15137 ;
  assign new_n20243 = new_n15137 & ~new_n16299 ;
  assign new_n20244 = ~new_n20242 & ~new_n20243 ;
  assign new_n20245 = lo0803 & new_n15454 ;
  assign new_n20246 = lo0958 & ~new_n13907 ;
  assign new_n20247 = ~lo0803 & ~lo0958 ;
  assign new_n20248 = ~new_n20246 & ~new_n20247 ;
  assign new_n20249 = ~new_n15454 & ~new_n20248 ;
  assign new_n20250 = ~new_n20245 & ~new_n20249 ;
  assign new_n20251 = lo0804 & ~new_n17223 ;
  assign new_n20252 = ~new_n13907 & new_n17223 ;
  assign new_n20253 = ~new_n20251 & ~new_n20252 ;
  assign new_n20254 = lo0805 & ~new_n15365 ;
  assign new_n20255 = lo0952 & ~new_n13907 ;
  assign new_n20256 = ~lo0952 & new_n7122 ;
  assign new_n20257 = ~new_n20255 & ~new_n20256 ;
  assign new_n20258 = new_n15365 & ~new_n20257 ;
  assign new_n20259 = ~new_n20254 & ~new_n20258 ;
  assign new_n20260 = lo0806 & ~new_n14924 ;
  assign new_n20261 = ~new_n5170 & ~new_n14927 ;
  assign new_n20262 = ~new_n13977 & new_n14927 ;
  assign new_n20263 = ~new_n20261 & ~new_n20262 ;
  assign new_n20264 = new_n14924 & ~new_n20263 ;
  assign new_n20265 = ~new_n20260 & ~new_n20264 ;
  assign new_n20266 = lo0807 & ~new_n14869 ;
  assign new_n20267 = ~new_n5170 & ~new_n14872 ;
  assign new_n20268 = ~new_n13977 & new_n14872 ;
  assign new_n20269 = ~new_n20267 & ~new_n20268 ;
  assign new_n20270 = new_n14869 & ~new_n20269 ;
  assign new_n20271 = ~new_n20266 & ~new_n20270 ;
  assign new_n20272 = lo0808 & ~new_n15016 ;
  assign new_n20273 = ~new_n5170 & ~new_n15019 ;
  assign new_n20274 = ~new_n13977 & new_n15019 ;
  assign new_n20275 = ~new_n20273 & ~new_n20274 ;
  assign new_n20276 = new_n15016 & ~new_n20275 ;
  assign new_n20277 = ~new_n20272 & ~new_n20276 ;
  assign new_n20278 = lo0809 & ~new_n15071 ;
  assign new_n20279 = ~new_n5170 & ~new_n15074 ;
  assign new_n20280 = ~new_n13977 & new_n15074 ;
  assign new_n20281 = ~new_n20279 & ~new_n20280 ;
  assign new_n20282 = new_n15071 & ~new_n20281 ;
  assign new_n20283 = ~new_n20278 & ~new_n20282 ;
  assign new_n20284 = lo0810 & ~new_n14848 ;
  assign new_n20285 = ~new_n5170 & ~new_n14853 ;
  assign new_n20286 = ~new_n13977 & new_n14853 ;
  assign new_n20287 = ~new_n20285 & ~new_n20286 ;
  assign new_n20288 = new_n14848 & ~new_n20287 ;
  assign new_n20289 = ~new_n20284 & ~new_n20288 ;
  assign new_n20290 = lo0811 & ~new_n14943 ;
  assign new_n20291 = ~new_n5170 & ~new_n14946 ;
  assign new_n20292 = ~new_n13977 & new_n14946 ;
  assign new_n20293 = ~new_n20291 & ~new_n20292 ;
  assign new_n20294 = new_n14943 & ~new_n20293 ;
  assign new_n20295 = ~new_n20290 & ~new_n20294 ;
  assign new_n20296 = lo0812 & ~new_n14997 ;
  assign new_n20297 = ~new_n5170 & ~new_n15000 ;
  assign new_n20298 = ~new_n13977 & new_n15000 ;
  assign new_n20299 = ~new_n20297 & ~new_n20298 ;
  assign new_n20300 = new_n14997 & ~new_n20299 ;
  assign new_n20301 = ~new_n20296 & ~new_n20300 ;
  assign new_n20302 = lo0813 & ~new_n15090 ;
  assign new_n20303 = ~new_n5170 & ~new_n15093 ;
  assign new_n20304 = ~new_n13977 & new_n15093 ;
  assign new_n20305 = ~new_n20303 & ~new_n20304 ;
  assign new_n20306 = new_n15090 & ~new_n20305 ;
  assign new_n20307 = ~new_n20302 & ~new_n20306 ;
  assign new_n20308 = lo0814 & ~new_n14886 ;
  assign new_n20309 = ~new_n5170 & ~new_n14889 ;
  assign new_n20310 = ~new_n13977 & new_n14889 ;
  assign new_n20311 = ~new_n20309 & ~new_n20310 ;
  assign new_n20312 = new_n14886 & ~new_n20311 ;
  assign new_n20313 = ~new_n20308 & ~new_n20312 ;
  assign new_n20314 = lo0815 & ~new_n14960 ;
  assign new_n20315 = ~new_n5170 & ~new_n14963 ;
  assign new_n20316 = ~new_n13977 & new_n14963 ;
  assign new_n20317 = ~new_n20315 & ~new_n20316 ;
  assign new_n20318 = new_n14960 & ~new_n20317 ;
  assign new_n20319 = ~new_n20314 & ~new_n20318 ;
  assign new_n20320 = lo0816 & ~new_n15033 ;
  assign new_n20321 = ~new_n5170 & ~new_n15036 ;
  assign new_n20322 = ~new_n13977 & new_n15036 ;
  assign new_n20323 = ~new_n20321 & ~new_n20322 ;
  assign new_n20324 = new_n15033 & ~new_n20323 ;
  assign new_n20325 = ~new_n20320 & ~new_n20324 ;
  assign new_n20326 = lo0817 & ~new_n15107 ;
  assign new_n20327 = ~new_n5170 & ~new_n15110 ;
  assign new_n20328 = ~new_n13977 & new_n15110 ;
  assign new_n20329 = ~new_n20327 & ~new_n20328 ;
  assign new_n20330 = new_n15107 & ~new_n20329 ;
  assign new_n20331 = ~new_n20326 & ~new_n20330 ;
  assign new_n20332 = lo0818 & ~new_n14977 ;
  assign new_n20333 = ~new_n5170 & ~new_n14980 ;
  assign new_n20334 = ~new_n13977 & new_n14980 ;
  assign new_n20335 = ~new_n20333 & ~new_n20334 ;
  assign new_n20336 = new_n14977 & ~new_n20335 ;
  assign new_n20337 = ~new_n20332 & ~new_n20336 ;
  assign new_n20338 = lo0819 & ~new_n14903 ;
  assign new_n20339 = ~new_n5170 & ~new_n14906 ;
  assign new_n20340 = ~new_n13977 & new_n14906 ;
  assign new_n20341 = ~new_n20339 & ~new_n20340 ;
  assign new_n20342 = new_n14903 & ~new_n20341 ;
  assign new_n20343 = ~new_n20338 & ~new_n20342 ;
  assign new_n20344 = lo0820 & ~new_n15050 ;
  assign new_n20345 = ~new_n5170 & ~new_n15053 ;
  assign new_n20346 = ~new_n13977 & new_n15053 ;
  assign new_n20347 = ~new_n20345 & ~new_n20346 ;
  assign new_n20348 = new_n15050 & ~new_n20347 ;
  assign new_n20349 = ~new_n20344 & ~new_n20348 ;
  assign new_n20350 = lo0821 & ~new_n15124 ;
  assign new_n20351 = ~new_n5170 & ~new_n15127 ;
  assign new_n20352 = ~new_n13977 & new_n15127 ;
  assign new_n20353 = ~new_n20351 & ~new_n20352 ;
  assign new_n20354 = new_n15124 & ~new_n20353 ;
  assign new_n20355 = ~new_n20350 & ~new_n20354 ;
  assign new_n20356 = lo0822 & new_n2252 ;
  assign new_n20357 = ~new_n15357 & ~new_n20356 ;
  assign new_n20358 = lo0823 & ~new_n17223 ;
  assign new_n20359 = ~new_n13977 & new_n17223 ;
  assign new_n20360 = ~new_n20358 & ~new_n20359 ;
  assign new_n20361 = lo0824 & ~new_n15365 ;
  assign new_n20362 = lo0952 & ~new_n13977 ;
  assign new_n20363 = ~lo0952 & ~new_n5170 ;
  assign new_n20364 = ~new_n20362 & ~new_n20363 ;
  assign new_n20365 = new_n15365 & ~new_n20364 ;
  assign new_n20366 = ~new_n20361 & ~new_n20365 ;
  assign new_n20367 = lo0825 & new_n15454 ;
  assign new_n20368 = lo0958 & ~new_n13977 ;
  assign new_n20369 = ~lo0958 & ~new_n13983 ;
  assign new_n20370 = ~new_n20368 & ~new_n20369 ;
  assign new_n20371 = ~new_n15454 & ~new_n20370 ;
  assign new_n20372 = ~new_n20367 & ~new_n20371 ;
  assign new_n20373 = lo0826 & ~new_n15376 ;
  assign new_n20374 = lo0855 & ~new_n3281 ;
  assign new_n20375 = lo0858 & ~new_n5170 ;
  assign new_n20376 = lo0859 & ~new_n13977 ;
  assign new_n20377 = lo0826 & ~lo0859 ;
  assign new_n20378 = ~new_n20376 & ~new_n20377 ;
  assign new_n20379 = ~lo0858 & ~new_n20378 ;
  assign new_n20380 = ~new_n20375 & ~new_n20379 ;
  assign new_n20381 = new_n15380 & ~new_n20380 ;
  assign new_n20382 = ~new_n20374 & ~new_n20381 ;
  assign new_n20383 = new_n15376 & ~new_n20382 ;
  assign new_n20384 = ~new_n20373 & ~new_n20383 ;
  assign new_n20385 = lo0827 & ~new_n14943 ;
  assign new_n20386 = new_n4530 & ~new_n14946 ;
  assign new_n20387 = ~new_n14234 & new_n14946 ;
  assign new_n20388 = ~new_n20386 & ~new_n20387 ;
  assign new_n20389 = new_n14943 & ~new_n20388 ;
  assign new_n20390 = ~new_n20385 & ~new_n20389 ;
  assign new_n20391 = lo0828 & ~new_n14924 ;
  assign new_n20392 = new_n4530 & ~new_n14927 ;
  assign new_n20393 = ~new_n14234 & new_n14927 ;
  assign new_n20394 = ~new_n20392 & ~new_n20393 ;
  assign new_n20395 = new_n14924 & ~new_n20394 ;
  assign new_n20396 = ~new_n20391 & ~new_n20395 ;
  assign new_n20397 = lo0829 & ~new_n14960 ;
  assign new_n20398 = new_n4530 & ~new_n14963 ;
  assign new_n20399 = ~new_n14234 & new_n14963 ;
  assign new_n20400 = ~new_n20398 & ~new_n20399 ;
  assign new_n20401 = new_n14960 & ~new_n20400 ;
  assign new_n20402 = ~new_n20397 & ~new_n20401 ;
  assign new_n20403 = lo0830 & ~new_n14977 ;
  assign new_n20404 = new_n4530 & ~new_n14980 ;
  assign new_n20405 = ~new_n14234 & new_n14980 ;
  assign new_n20406 = ~new_n20404 & ~new_n20405 ;
  assign new_n20407 = new_n14977 & ~new_n20406 ;
  assign new_n20408 = ~new_n20403 & ~new_n20407 ;
  assign new_n20409 = lo0831 & ~new_n14869 ;
  assign new_n20410 = new_n4530 & ~new_n14872 ;
  assign new_n20411 = ~new_n14234 & new_n14872 ;
  assign new_n20412 = ~new_n20410 & ~new_n20411 ;
  assign new_n20413 = new_n14869 & ~new_n20412 ;
  assign new_n20414 = ~new_n20409 & ~new_n20413 ;
  assign new_n20415 = lo0832 & ~new_n14848 ;
  assign new_n20416 = new_n4530 & ~new_n14853 ;
  assign new_n20417 = ~new_n14234 & new_n14853 ;
  assign new_n20418 = ~new_n20416 & ~new_n20417 ;
  assign new_n20419 = new_n14848 & ~new_n20418 ;
  assign new_n20420 = ~new_n20415 & ~new_n20419 ;
  assign new_n20421 = lo0833 & ~new_n14886 ;
  assign new_n20422 = new_n4530 & ~new_n14889 ;
  assign new_n20423 = ~new_n14234 & new_n14889 ;
  assign new_n20424 = ~new_n20422 & ~new_n20423 ;
  assign new_n20425 = new_n14886 & ~new_n20424 ;
  assign new_n20426 = ~new_n20421 & ~new_n20425 ;
  assign new_n20427 = lo0834 & ~new_n14903 ;
  assign new_n20428 = new_n4530 & ~new_n14906 ;
  assign new_n20429 = ~new_n14234 & new_n14906 ;
  assign new_n20430 = ~new_n20428 & ~new_n20429 ;
  assign new_n20431 = new_n14903 & ~new_n20430 ;
  assign new_n20432 = ~new_n20427 & ~new_n20431 ;
  assign new_n20433 = lo0835 & ~new_n15016 ;
  assign new_n20434 = new_n4530 & ~new_n15019 ;
  assign new_n20435 = ~new_n14234 & new_n15019 ;
  assign new_n20436 = ~new_n20434 & ~new_n20435 ;
  assign new_n20437 = new_n15016 & ~new_n20436 ;
  assign new_n20438 = ~new_n20433 & ~new_n20437 ;
  assign new_n20439 = lo0836 & ~new_n14997 ;
  assign new_n20440 = new_n4530 & ~new_n15000 ;
  assign new_n20441 = ~new_n14234 & new_n15000 ;
  assign new_n20442 = ~new_n20440 & ~new_n20441 ;
  assign new_n20443 = new_n14997 & ~new_n20442 ;
  assign new_n20444 = ~new_n20439 & ~new_n20443 ;
  assign new_n20445 = lo0837 & ~new_n15033 ;
  assign new_n20446 = new_n4530 & ~new_n15036 ;
  assign new_n20447 = ~new_n14234 & new_n15036 ;
  assign new_n20448 = ~new_n20446 & ~new_n20447 ;
  assign new_n20449 = new_n15033 & ~new_n20448 ;
  assign new_n20450 = ~new_n20445 & ~new_n20449 ;
  assign new_n20451 = lo0838 & ~new_n15050 ;
  assign new_n20452 = new_n4530 & ~new_n15053 ;
  assign new_n20453 = ~new_n14234 & new_n15053 ;
  assign new_n20454 = ~new_n20452 & ~new_n20453 ;
  assign new_n20455 = new_n15050 & ~new_n20454 ;
  assign new_n20456 = ~new_n20451 & ~new_n20455 ;
  assign new_n20457 = lo0839 & ~new_n15090 ;
  assign new_n20458 = new_n4530 & ~new_n15093 ;
  assign new_n20459 = ~new_n14234 & new_n15093 ;
  assign new_n20460 = ~new_n20458 & ~new_n20459 ;
  assign new_n20461 = new_n15090 & ~new_n20460 ;
  assign new_n20462 = ~new_n20457 & ~new_n20461 ;
  assign new_n20463 = lo0840 & ~new_n15071 ;
  assign new_n20464 = new_n4530 & ~new_n15074 ;
  assign new_n20465 = ~new_n14234 & new_n15074 ;
  assign new_n20466 = ~new_n20464 & ~new_n20465 ;
  assign new_n20467 = new_n15071 & ~new_n20466 ;
  assign new_n20468 = ~new_n20463 & ~new_n20467 ;
  assign new_n20469 = lo0841 & ~new_n15107 ;
  assign new_n20470 = new_n4530 & ~new_n15110 ;
  assign new_n20471 = ~new_n14234 & new_n15110 ;
  assign new_n20472 = ~new_n20470 & ~new_n20471 ;
  assign new_n20473 = new_n15107 & ~new_n20472 ;
  assign new_n20474 = ~new_n20469 & ~new_n20473 ;
  assign new_n20475 = lo0842 & ~new_n15124 ;
  assign new_n20476 = new_n4530 & ~new_n15127 ;
  assign new_n20477 = ~new_n14234 & new_n15127 ;
  assign new_n20478 = ~new_n20476 & ~new_n20477 ;
  assign new_n20479 = new_n15124 & ~new_n20478 ;
  assign new_n20480 = ~new_n20475 & ~new_n20479 ;
  assign new_n20481 = lo0843 & new_n15454 ;
  assign new_n20482 = lo0958 & ~new_n14234 ;
  assign new_n20483 = ~lo0958 & ~new_n14238 ;
  assign new_n20484 = ~new_n20482 & ~new_n20483 ;
  assign new_n20485 = ~new_n15454 & ~new_n20484 ;
  assign new_n20486 = ~new_n20481 & ~new_n20485 ;
  assign new_n20487 = lo0844 & ~new_n15365 ;
  assign new_n20488 = lo0952 & ~new_n14234 ;
  assign new_n20489 = ~lo0952 & new_n4530 ;
  assign new_n20490 = ~new_n20488 & ~new_n20489 ;
  assign new_n20491 = new_n15365 & ~new_n20490 ;
  assign new_n20492 = ~new_n20487 & ~new_n20491 ;
  assign new_n20493 = lo0845 & ~new_n17223 ;
  assign new_n20494 = ~new_n14234 & new_n17223 ;
  assign new_n20495 = ~new_n20493 & ~new_n20494 ;
  assign new_n20496 = lo0846 & ~new_n14699 ;
  assign new_n20497 = new_n2450 & new_n12460 ;
  assign new_n20498 = ~new_n17359 & ~new_n20497 ;
  assign new_n20499 = new_n12553 & new_n14699 ;
  assign new_n20500 = ~new_n20498 & new_n20499 ;
  assign new_n20501 = new_n17356 & new_n20500 ;
  assign new_n20502 = ~new_n20496 & ~new_n20501 ;
  assign new_n20503 = lo0847 & new_n2252 ;
  assign new_n20504 = ~new_n2450 & new_n12508 ;
  assign new_n20505 = new_n12524 & new_n20504 ;
  assign new_n20506 = new_n12509 & new_n20505 ;
  assign new_n20507 = ~new_n2446 & new_n13286 ;
  assign new_n20508 = new_n12796 & new_n20507 ;
  assign new_n20509 = new_n2446 & new_n12851 ;
  assign new_n20510 = ~new_n20508 & ~new_n20509 ;
  assign new_n20511 = new_n12768 & ~new_n20510 ;
  assign new_n20512 = ~new_n20506 & ~new_n20511 ;
  assign new_n20513 = ~new_n2252 & new_n2454 ;
  assign new_n20514 = ~new_n20512 & new_n20513 ;
  assign new_n20515 = new_n15451 & new_n20514 ;
  assign new_n20516 = ~new_n20503 & ~new_n20515 ;
  assign new_n20517 = lo0848 & new_n2252 ;
  assign new_n20518 = new_n2446 & new_n15451 ;
  assign new_n20519 = ~new_n12329 & ~new_n12933 ;
  assign new_n20520 = ~new_n2252 & ~new_n2450 ;
  assign new_n20521 = new_n13819 & new_n20520 ;
  assign new_n20522 = ~new_n13513 & new_n20521 ;
  assign new_n20523 = ~new_n20519 & new_n20522 ;
  assign new_n20524 = new_n20518 & new_n20523 ;
  assign new_n20525 = ~new_n20517 & ~new_n20524 ;
  assign new_n20526 = lo0849 & new_n2252 ;
  assign new_n20527 = new_n12524 & new_n12720 ;
  assign new_n20528 = new_n2454 & new_n20527 ;
  assign new_n20529 = new_n12441 & ~new_n12933 ;
  assign new_n20530 = ~new_n2454 & new_n12420 ;
  assign new_n20531 = ~new_n20529 & new_n20530 ;
  assign new_n20532 = ~new_n20528 & ~new_n20531 ;
  assign new_n20533 = new_n20504 & ~new_n20532 ;
  assign new_n20534 = new_n12523 & new_n12549 ;
  assign new_n20535 = ~new_n12329 & new_n12420 ;
  assign new_n20536 = new_n2446 & new_n20535 ;
  assign new_n20537 = new_n20534 & new_n20536 ;
  assign new_n20538 = ~new_n16898 & ~new_n20537 ;
  assign new_n20539 = new_n2455 & ~new_n20538 ;
  assign new_n20540 = ~new_n20533 & ~new_n20539 ;
  assign new_n20541 = ~new_n2252 & ~new_n20540 ;
  assign new_n20542 = new_n15451 & new_n20541 ;
  assign new_n20543 = ~new_n20526 & ~new_n20542 ;
  assign new_n20544 = lo0850 & ~new_n14699 ;
  assign new_n20545 = new_n2455 & new_n12420 ;
  assign new_n20546 = new_n20534 & new_n20545 ;
  assign new_n20547 = new_n2454 & ~new_n20527 ;
  assign new_n20548 = ~new_n2450 & ~new_n20547 ;
  assign new_n20549 = ~new_n20546 & ~new_n20548 ;
  assign new_n20550 = new_n2454 & ~new_n16901 ;
  assign new_n20551 = ~new_n13512 & ~new_n20550 ;
  assign new_n20552 = ~new_n20549 & ~new_n20551 ;
  assign new_n20553 = new_n20518 & new_n20552 ;
  assign new_n20554 = ~new_n2454 & ~new_n12513 ;
  assign new_n20555 = new_n20553 & ~new_n20554 ;
  assign new_n20556 = ~new_n12452 & new_n14699 ;
  assign new_n20557 = new_n20555 & new_n20556 ;
  assign new_n20558 = ~new_n20544 & ~new_n20557 ;
  assign new_n20559 = lo0851 & ~new_n14699 ;
  assign new_n20560 = ~new_n12429 & new_n14699 ;
  assign new_n20561 = new_n20555 & new_n20560 ;
  assign new_n20562 = ~new_n20559 & ~new_n20561 ;
  assign new_n20563 = lo0852 & ~new_n14699 ;
  assign new_n20564 = ~new_n2454 & ~new_n12420 ;
  assign new_n20565 = ~new_n12441 & new_n14699 ;
  assign new_n20566 = ~new_n20564 & new_n20565 ;
  assign new_n20567 = new_n20553 & new_n20566 ;
  assign new_n20568 = ~new_n20563 & ~new_n20567 ;
  assign new_n20569 = lo0853 & new_n2252 ;
  assign new_n20570 = ~new_n2252 & new_n12460 ;
  assign new_n20571 = new_n12848 & new_n20570 ;
  assign new_n20572 = new_n17339 & new_n20571 ;
  assign new_n20573 = ~new_n20569 & ~new_n20572 ;
  assign new_n20574 = lo0854 & new_n2252 ;
  assign new_n20575 = new_n12698 & new_n15361 ;
  assign new_n20576 = new_n12569 & new_n20575 ;
  assign new_n20577 = new_n20518 & new_n20576 ;
  assign new_n20578 = ~new_n20574 & ~new_n20577 ;
  assign new_n20579 = lo0855 & new_n2252 ;
  assign new_n20580 = ~new_n2252 & new_n13424 ;
  assign new_n20581 = new_n12721 & new_n20580 ;
  assign new_n20582 = new_n20518 & new_n20581 ;
  assign new_n20583 = ~new_n20579 & ~new_n20582 ;
  assign new_n20584 = lo0856 & new_n2252 ;
  assign new_n20585 = new_n2455 & new_n20518 ;
  assign new_n20586 = new_n13046 & new_n20585 ;
  assign new_n20587 = ~new_n12429 & new_n12460 ;
  assign new_n20588 = new_n12429 & ~new_n12460 ;
  assign new_n20589 = ~new_n2252 & new_n12441 ;
  assign new_n20590 = new_n12467 & new_n20589 ;
  assign new_n20591 = ~new_n20588 & new_n20590 ;
  assign new_n20592 = ~new_n20587 & new_n20591 ;
  assign new_n20593 = new_n20586 & new_n20592 ;
  assign new_n20594 = ~new_n20584 & ~new_n20593 ;
  assign new_n20595 = lo0857 & new_n2252 ;
  assign new_n20596 = ~new_n2252 & new_n12525 ;
  assign new_n20597 = new_n20586 & new_n20596 ;
  assign new_n20598 = ~new_n20595 & ~new_n20597 ;
  assign new_n20599 = lo0858 & new_n2252 ;
  assign new_n20600 = lo1067 & ~new_n2252 ;
  assign new_n20601 = ~new_n20599 & ~new_n20600 ;
  assign new_n20602 = lo0859 & new_n2252 ;
  assign new_n20603 = new_n12550 & new_n12720 ;
  assign new_n20604 = new_n17339 & new_n20603 ;
  assign new_n20605 = new_n14806 & new_n20604 ;
  assign new_n20606 = ~new_n20602 & ~new_n20605 ;
  assign new_n20607 = lo0860 & ~new_n16687 ;
  assign new_n20608 = lo1424 & new_n16687 ;
  assign new_n20609 = ~new_n20607 & ~new_n20608 ;
  assign new_n20610 = lo0861 & ~new_n15612 ;
  assign new_n20611 = ~new_n12417 & new_n15612 ;
  assign new_n20612 = ~new_n20610 & ~new_n20611 ;
  assign new_n20613 = lo0862 & ~new_n16687 ;
  assign new_n20614 = lo1421 & new_n16687 ;
  assign new_n20615 = ~new_n20613 & ~new_n20614 ;
  assign new_n20616 = lo0863 & ~new_n15612 ;
  assign new_n20617 = ~new_n12426 & new_n15612 ;
  assign new_n20618 = ~new_n20616 & ~new_n20617 ;
  assign new_n20619 = lo0864 & ~new_n16687 ;
  assign new_n20620 = lo1422 & new_n16687 ;
  assign new_n20621 = ~new_n20619 & ~new_n20620 ;
  assign new_n20622 = lo0865 & ~new_n15612 ;
  assign new_n20623 = ~new_n12438 & new_n15612 ;
  assign new_n20624 = ~new_n20622 & ~new_n20623 ;
  assign new_n20625 = lo0866 & ~new_n16687 ;
  assign new_n20626 = lo1423 & new_n16687 ;
  assign new_n20627 = ~new_n20625 & ~new_n20626 ;
  assign new_n20628 = lo0867 & ~new_n15612 ;
  assign new_n20629 = ~new_n12449 & new_n15612 ;
  assign new_n20630 = ~new_n20628 & ~new_n20629 ;
  assign new_n20631 = lo0868 & ~new_n15612 ;
  assign new_n20632 = new_n12458 & new_n15612 ;
  assign new_n20633 = ~new_n20631 & ~new_n20632 ;
  assign new_n20634 = lo0869 & ~new_n16687 ;
  assign new_n20635 = lo1280 & new_n16687 ;
  assign new_n20636 = ~new_n20634 & ~new_n20635 ;
  assign new_n20637 = lo0870 & ~new_n15612 ;
  assign new_n20638 = new_n12465 & new_n15612 ;
  assign new_n20639 = ~new_n20637 & ~new_n20638 ;
  assign new_n20640 = lo0871 & ~new_n16687 ;
  assign new_n20641 = lo1281 & new_n16687 ;
  assign new_n20642 = ~new_n20640 & ~new_n20641 ;
  assign new_n20643 = lo0872 & new_n2252 ;
  assign new_n20644 = ~new_n12442 & new_n12508 ;
  assign new_n20645 = new_n12720 & new_n20644 ;
  assign new_n20646 = ~new_n12329 & ~new_n12368 ;
  assign new_n20647 = ~new_n13558 & ~new_n20646 ;
  assign new_n20648 = ~new_n2446 & new_n13781 ;
  assign new_n20649 = ~new_n20647 & new_n20648 ;
  assign new_n20650 = ~new_n20645 & ~new_n20649 ;
  assign new_n20651 = new_n2455 & ~new_n20650 ;
  assign new_n20652 = new_n12405 & new_n20535 ;
  assign new_n20653 = new_n13403 & new_n20652 ;
  assign new_n20654 = ~new_n12402 & ~new_n20653 ;
  assign new_n20655 = ~new_n20651 & new_n20654 ;
  assign new_n20656 = new_n2454 & ~new_n20655 ;
  assign new_n20657 = ~new_n2454 & new_n20655 ;
  assign new_n20658 = ~new_n20656 & ~new_n20657 ;
  assign new_n20659 = ~new_n12508 & ~new_n20658 ;
  assign new_n20660 = new_n12508 & new_n20656 ;
  assign new_n20661 = ~new_n2446 & new_n12472 ;
  assign new_n20662 = new_n17100 & new_n20661 ;
  assign new_n20663 = ~new_n2454 & new_n20662 ;
  assign new_n20664 = ~new_n20655 & new_n20663 ;
  assign new_n20665 = ~new_n20660 & ~new_n20664 ;
  assign new_n20666 = ~new_n20659 & new_n20665 ;
  assign new_n20667 = ~new_n2252 & ~new_n20666 ;
  assign new_n20668 = new_n15451 & new_n20667 ;
  assign new_n20669 = ~new_n20643 & ~new_n20668 ;
  assign new_n20670 = lo0873 & ~new_n14699 ;
  assign new_n20671 = ~new_n2454 & ~new_n12404 ;
  assign new_n20672 = ~new_n2446 & new_n12404 ;
  assign new_n20673 = ~new_n20671 & ~new_n20672 ;
  assign new_n20674 = ~new_n12404 & new_n20673 ;
  assign new_n20675 = new_n13098 & new_n20674 ;
  assign new_n20676 = ~new_n12404 & ~new_n20673 ;
  assign new_n20677 = new_n12404 & new_n13144 ;
  assign new_n20678 = new_n20673 & new_n20677 ;
  assign new_n20679 = ~new_n20676 & ~new_n20678 ;
  assign new_n20680 = ~new_n20675 & new_n20679 ;
  assign new_n20681 = new_n20673 & ~new_n20680 ;
  assign new_n20682 = ~new_n20673 & new_n20680 ;
  assign new_n20683 = ~new_n20681 & ~new_n20682 ;
  assign new_n20684 = ~new_n12357 & ~new_n20683 ;
  assign new_n20685 = new_n12357 & new_n20681 ;
  assign new_n20686 = new_n20662 & ~new_n20673 ;
  assign new_n20687 = ~new_n20680 & new_n20686 ;
  assign new_n20688 = ~new_n20685 & ~new_n20687 ;
  assign new_n20689 = ~new_n20684 & new_n20688 ;
  assign new_n20690 = new_n2450 & ~new_n13030 ;
  assign new_n20691 = ~new_n2450 & ~new_n20535 ;
  assign new_n20692 = new_n2446 & ~new_n20691 ;
  assign new_n20693 = ~new_n20690 & new_n20692 ;
  assign new_n20694 = new_n20674 & ~new_n20693 ;
  assign new_n20695 = new_n14699 & ~new_n20694 ;
  assign new_n20696 = ~new_n20689 & new_n20695 ;
  assign new_n20697 = ~new_n20670 & ~new_n20696 ;
  assign new_n20698 = lo0874 & ~new_n14699 ;
  assign new_n20699 = new_n12325 & ~new_n12404 ;
  assign new_n20700 = new_n12325 & ~new_n20699 ;
  assign new_n20701 = ~new_n20673 & ~new_n20700 ;
  assign new_n20702 = ~new_n12329 & new_n20673 ;
  assign new_n20703 = ~new_n12325 & new_n12404 ;
  assign new_n20704 = new_n20702 & new_n20703 ;
  assign new_n20705 = ~new_n20701 & ~new_n20704 ;
  assign new_n20706 = new_n12404 & ~new_n20705 ;
  assign new_n20707 = ~new_n12404 & new_n20705 ;
  assign new_n20708 = ~new_n20706 & ~new_n20707 ;
  assign new_n20709 = new_n13317 & ~new_n20708 ;
  assign new_n20710 = ~new_n13317 & new_n20706 ;
  assign new_n20711 = ~new_n12404 & new_n20662 ;
  assign new_n20712 = ~new_n20705 & new_n20711 ;
  assign new_n20713 = ~new_n20710 & ~new_n20712 ;
  assign new_n20714 = ~new_n20709 & new_n20713 ;
  assign new_n20715 = new_n20695 & ~new_n20714 ;
  assign new_n20716 = ~new_n20698 & ~new_n20715 ;
  assign new_n20717 = lo0875 & ~new_n14699 ;
  assign new_n20718 = new_n13179 & new_n20674 ;
  assign new_n20719 = new_n12404 & new_n13218 ;
  assign new_n20720 = new_n20673 & new_n20719 ;
  assign new_n20721 = ~new_n20676 & ~new_n20720 ;
  assign new_n20722 = ~new_n20718 & new_n20721 ;
  assign new_n20723 = new_n20673 & ~new_n20722 ;
  assign new_n20724 = ~new_n20673 & new_n20722 ;
  assign new_n20725 = ~new_n20723 & ~new_n20724 ;
  assign new_n20726 = ~new_n2465 & ~new_n20725 ;
  assign new_n20727 = new_n2465 & new_n20723 ;
  assign new_n20728 = new_n20686 & ~new_n20722 ;
  assign new_n20729 = ~new_n20727 & ~new_n20728 ;
  assign new_n20730 = ~new_n20726 & new_n20729 ;
  assign new_n20731 = new_n20695 & ~new_n20730 ;
  assign new_n20732 = ~new_n20717 & ~new_n20731 ;
  assign new_n20733 = lo0876 & ~new_n14699 ;
  assign new_n20734 = new_n12367 & ~new_n12404 ;
  assign new_n20735 = new_n12367 & ~new_n20734 ;
  assign new_n20736 = ~new_n20673 & ~new_n20735 ;
  assign new_n20737 = ~new_n12367 & new_n12404 ;
  assign new_n20738 = new_n20702 & new_n20737 ;
  assign new_n20739 = ~new_n20736 & ~new_n20738 ;
  assign new_n20740 = new_n12404 & ~new_n20739 ;
  assign new_n20741 = ~new_n12404 & new_n20739 ;
  assign new_n20742 = ~new_n20740 & ~new_n20741 ;
  assign new_n20743 = new_n12939 & ~new_n20742 ;
  assign new_n20744 = ~new_n12939 & new_n20740 ;
  assign new_n20745 = new_n20711 & ~new_n20739 ;
  assign new_n20746 = ~new_n20744 & ~new_n20745 ;
  assign new_n20747 = ~new_n20743 & new_n20746 ;
  assign new_n20748 = new_n20695 & ~new_n20747 ;
  assign new_n20749 = ~new_n20733 & ~new_n20748 ;
  assign new_n20750 = lo0877 & ~new_n15612 ;
  assign new_n20751 = new_n13103 & new_n15612 ;
  assign new_n20752 = ~new_n20750 & ~new_n20751 ;
  assign new_n20753 = lo0878 & ~new_n16687 ;
  assign new_n20754 = lo1283 & new_n16687 ;
  assign new_n20755 = ~new_n20753 & ~new_n20754 ;
  assign new_n20756 = lo0879 & ~new_n15612 ;
  assign new_n20757 = new_n13322 & new_n15612 ;
  assign new_n20758 = ~new_n20756 & ~new_n20757 ;
  assign new_n20759 = lo0880 & ~new_n16687 ;
  assign new_n20760 = lo1282 & new_n16687 ;
  assign new_n20761 = ~new_n20759 & ~new_n20760 ;
  assign new_n20762 = lo0881 & new_n2252 ;
  assign new_n20763 = new_n12553 & new_n17339 ;
  assign new_n20764 = new_n12550 & new_n20763 ;
  assign new_n20765 = new_n17927 & new_n20764 ;
  assign new_n20766 = ~new_n20762 & ~new_n20765 ;
  assign new_n20767 = lo0882 & new_n2252 ;
  assign new_n20768 = new_n2455 & new_n12721 ;
  assign new_n20769 = ~new_n13824 & ~new_n20768 ;
  assign new_n20770 = new_n12329 & ~new_n20769 ;
  assign new_n20771 = new_n20518 & new_n20770 ;
  assign new_n20772 = ~new_n2252 & new_n20771 ;
  assign new_n20773 = ~new_n20767 & ~new_n20772 ;
  assign new_n20774 = lo0883 & new_n2252 ;
  assign new_n20775 = lo0884 & ~new_n2252 ;
  assign new_n20776 = ~new_n20774 & ~new_n20775 ;
  assign new_n20777 = lo0884 & new_n2252 ;
  assign new_n20778 = lo0885 & ~new_n2252 ;
  assign new_n20779 = ~new_n20777 & ~new_n20778 ;
  assign new_n20780 = lo0885 & new_n2252 ;
  assign new_n20781 = new_n13826 & new_n20535 ;
  assign new_n20782 = new_n15451 & new_n20781 ;
  assign new_n20783 = ~new_n12420 & new_n12443 ;
  assign new_n20784 = ~new_n12329 & ~new_n20783 ;
  assign new_n20785 = new_n12383 & ~new_n20784 ;
  assign new_n20786 = ~new_n20782 & ~new_n20785 ;
  assign new_n20787 = new_n12442 & new_n13030 ;
  assign new_n20788 = ~new_n12479 & ~new_n20787 ;
  assign new_n20789 = new_n13807 & ~new_n20788 ;
  assign new_n20790 = ~new_n2252 & new_n20789 ;
  assign new_n20791 = ~new_n20786 & new_n20790 ;
  assign new_n20792 = ~new_n20780 & ~new_n20791 ;
  assign new_n20793 = ~lo0945 & lo0946 ;
  assign new_n20794 = lo0942 & ~new_n2252 ;
  assign new_n20795 = lo0943 & new_n20794 ;
  assign new_n20796 = new_n13842 & new_n20795 ;
  assign new_n20797 = new_n20793 & new_n20796 ;
  assign new_n20798 = lo0944 & new_n20797 ;
  assign new_n20799 = ~lo0947 & lo0948 ;
  assign new_n20800 = lo0959 & new_n20799 ;
  assign new_n20801 = new_n20798 & new_n20800 ;
  assign new_n20802 = ~lo1068 & new_n20801 ;
  assign new_n20803 = lo0948 & ~lo0959 ;
  assign new_n20804 = ~lo0947 & new_n20803 ;
  assign new_n20805 = ~lo0944 & new_n20804 ;
  assign new_n20806 = new_n20797 & new_n20805 ;
  assign new_n20807 = ~lo0946 & lo0947 ;
  assign new_n20808 = lo0945 & new_n20807 ;
  assign new_n20809 = new_n20803 & new_n20808 ;
  assign new_n20810 = new_n20796 & new_n20809 ;
  assign new_n20811 = ~lo0944 & new_n20810 ;
  assign new_n20812 = lo0944 & new_n20810 ;
  assign new_n20813 = new_n20798 & new_n20804 ;
  assign new_n20814 = lo1068 & new_n20813 ;
  assign new_n20815 = ~lo1068 & new_n20813 ;
  assign new_n20816 = lo0892 & ~new_n13928 ;
  assign new_n20817 = ~new_n10308 & ~new_n13940 ;
  assign new_n20818 = lo0759 & new_n2261 ;
  assign new_n20819 = ~new_n2261 & ~new_n14616 ;
  assign new_n20820 = ~new_n20818 & ~new_n20819 ;
  assign new_n20821 = new_n13940 & ~new_n20820 ;
  assign new_n20822 = ~new_n20817 & ~new_n20821 ;
  assign new_n20823 = new_n13928 & ~new_n20822 ;
  assign new_n20824 = ~new_n20816 & ~new_n20823 ;
  assign new_n20825 = lo0893 & ~new_n13928 ;
  assign new_n20826 = ~new_n13907 & ~new_n13940 ;
  assign new_n20827 = ~lo0803 & new_n2261 ;
  assign new_n20828 = ~new_n2261 & ~new_n14605 ;
  assign new_n20829 = ~new_n20827 & ~new_n20828 ;
  assign new_n20830 = new_n13940 & ~new_n20829 ;
  assign new_n20831 = ~new_n20826 & ~new_n20830 ;
  assign new_n20832 = new_n13928 & ~new_n20831 ;
  assign new_n20833 = ~new_n20825 & ~new_n20832 ;
  assign new_n20834 = lo0895 & new_n2252 ;
  assign new_n20835 = new_n12329 & new_n12591 ;
  assign new_n20836 = new_n2264 & ~new_n12357 ;
  assign new_n20837 = ~new_n12863 & ~new_n20836 ;
  assign new_n20838 = ~new_n12325 & ~new_n20837 ;
  assign new_n20839 = ~new_n15591 & ~new_n20838 ;
  assign new_n20840 = ~new_n12329 & ~new_n20839 ;
  assign new_n20841 = ~new_n20835 & ~new_n20840 ;
  assign new_n20842 = ~new_n2446 & ~new_n20841 ;
  assign new_n20843 = new_n12329 & new_n12840 ;
  assign new_n20844 = new_n2264 & new_n12523 ;
  assign new_n20845 = new_n12443 & new_n20844 ;
  assign new_n20846 = ~new_n12605 & ~new_n20845 ;
  assign new_n20847 = new_n12486 & ~new_n20846 ;
  assign new_n20848 = ~new_n20843 & ~new_n20847 ;
  assign new_n20849 = new_n2446 & ~new_n20848 ;
  assign new_n20850 = new_n2454 & ~new_n20849 ;
  assign new_n20851 = ~new_n20842 & new_n20850 ;
  assign new_n20852 = new_n2450 & ~new_n20851 ;
  assign new_n20853 = new_n12420 & ~new_n13829 ;
  assign new_n20854 = new_n12329 & ~new_n20853 ;
  assign new_n20855 = new_n12646 & ~new_n13296 ;
  assign new_n20856 = ~new_n20854 & new_n20855 ;
  assign new_n20857 = ~new_n15537 & ~new_n20856 ;
  assign new_n20858 = ~new_n20852 & new_n20857 ;
  assign new_n20859 = ~new_n2252 & ~new_n20858 ;
  assign new_n20860 = new_n15451 & new_n20859 ;
  assign new_n20861 = ~new_n20834 & ~new_n20860 ;
  assign new_n20862 = ~lo0048 & ~lo0897 ;
  assign new_n20863 = lo0050 & ~new_n20862 ;
  assign new_n20864 = lo0896 & ~new_n20863 ;
  assign new_n20865 = lo1069 & ~new_n14656 ;
  assign new_n20866 = ~lo0977 & lo1072 ;
  assign new_n20867 = ~lo0980 & new_n20866 ;
  assign new_n20868 = lo0977 & lo0980 ;
  assign new_n20869 = ~lo0977 & lo1071 ;
  assign new_n20870 = lo0980 & new_n20869 ;
  assign new_n20871 = ~new_n20868 & ~new_n20870 ;
  assign new_n20872 = ~new_n20867 & new_n20871 ;
  assign new_n20873 = ~lo0977 & ~new_n20872 ;
  assign new_n20874 = lo0977 & new_n20872 ;
  assign new_n20875 = ~new_n20873 & ~new_n20874 ;
  assign new_n20876 = lo1070 & ~new_n20875 ;
  assign new_n20877 = ~lo1070 & new_n20873 ;
  assign new_n20878 = lo0977 & lo1073 ;
  assign new_n20879 = ~new_n20872 & new_n20878 ;
  assign new_n20880 = ~new_n20877 & ~new_n20879 ;
  assign new_n20881 = ~new_n20876 & new_n20880 ;
  assign new_n20882 = new_n14656 & ~new_n20881 ;
  assign new_n20883 = ~new_n20865 & ~new_n20882 ;
  assign new_n20884 = new_n20863 & ~new_n20883 ;
  assign new_n20885 = ~new_n20864 & ~new_n20884 ;
  assign new_n20886 = ~lo0048 & ~lo1447 ;
  assign new_n20887 = ~pi015 & new_n20886 ;
  assign new_n20888 = ~lo1450 & lo1451 ;
  assign new_n20889 = lo1448 & ~lo1449 ;
  assign new_n20890 = new_n20888 & new_n20889 ;
  assign new_n20891 = lo0902 & new_n2252 ;
  assign new_n20892 = lo0872 & ~new_n2252 ;
  assign new_n20893 = ~new_n20891 & ~new_n20892 ;
  assign new_n20894 = lo0903 & ~new_n14699 ;
  assign new_n20895 = lo0874 & new_n14699 ;
  assign new_n20896 = ~new_n20894 & ~new_n20895 ;
  assign new_n20897 = lo0904 & ~new_n14699 ;
  assign new_n20898 = lo0873 & new_n14699 ;
  assign new_n20899 = ~new_n20897 & ~new_n20898 ;
  assign new_n20900 = lo0905 & ~new_n14699 ;
  assign new_n20901 = lo0876 & new_n14699 ;
  assign new_n20902 = ~new_n20900 & ~new_n20901 ;
  assign new_n20903 = lo0906 & ~new_n14699 ;
  assign new_n20904 = lo0875 & new_n14699 ;
  assign new_n20905 = ~new_n20903 & ~new_n20904 ;
  assign new_n20906 = lo0907 & new_n2252 ;
  assign new_n20907 = lo0881 & ~new_n2252 ;
  assign new_n20908 = ~new_n20906 & ~new_n20907 ;
  assign new_n20909 = lo0908 & new_n2252 ;
  assign new_n20910 = ~new_n2252 & ~new_n13312 ;
  assign new_n20911 = new_n15451 & new_n20910 ;
  assign new_n20912 = ~new_n20909 & ~new_n20911 ;
  assign new_n20913 = lo0909 & ~new_n14699 ;
  assign new_n20914 = ~new_n13094 & new_n14699 ;
  assign new_n20915 = ~new_n20913 & ~new_n20914 ;
  assign new_n20916 = lo0910 & ~new_n14699 ;
  assign new_n20917 = ~new_n13246 & new_n14699 ;
  assign new_n20918 = ~new_n20916 & ~new_n20917 ;
  assign new_n20919 = lo0911 & ~new_n14699 ;
  assign new_n20920 = ~new_n13390 & new_n14699 ;
  assign new_n20921 = ~new_n20919 & ~new_n20920 ;
  assign new_n20922 = lo0912 & ~new_n14699 ;
  assign new_n20923 = ~new_n13172 & new_n14699 ;
  assign new_n20924 = ~new_n20922 & ~new_n20923 ;
  assign new_n20925 = lo0913 & new_n2252 ;
  assign new_n20926 = lo1076 & ~new_n2252 ;
  assign new_n20927 = ~new_n20925 & ~new_n20926 ;
  assign new_n20928 = lo0914 & ~new_n13928 ;
  assign new_n20929 = lo0113 & new_n13928 ;
  assign new_n20930 = ~new_n20928 & ~new_n20929 ;
  assign new_n20931 = lo0915 & ~new_n13928 ;
  assign new_n20932 = lo0114 & new_n13928 ;
  assign new_n20933 = ~new_n20931 & ~new_n20932 ;
  assign new_n20934 = new_n1942 & new_n14668 ;
  assign new_n20935 = lo0916 & ~new_n20934 ;
  assign new_n20936 = lo1444 & new_n20934 ;
  assign new_n20937 = ~new_n20935 & ~new_n20936 ;
  assign new_n20938 = lo0917 & ~new_n13928 ;
  assign new_n20939 = new_n13978 & ~new_n19223 ;
  assign new_n20940 = ~new_n13937 & ~new_n19334 ;
  assign new_n20941 = new_n13943 & new_n20940 ;
  assign new_n20942 = ~new_n13955 & ~new_n20941 ;
  assign new_n20943 = ~new_n20939 & new_n20942 ;
  assign new_n20944 = ~new_n13937 & ~new_n20943 ;
  assign new_n20945 = new_n13937 & new_n20943 ;
  assign new_n20946 = ~new_n20944 & ~new_n20945 ;
  assign new_n20947 = ~new_n6917 & ~new_n20946 ;
  assign new_n20948 = new_n6917 & new_n20944 ;
  assign new_n20949 = lo0643 & new_n13937 ;
  assign new_n20950 = ~new_n20943 & new_n20949 ;
  assign new_n20951 = ~new_n20948 & ~new_n20950 ;
  assign new_n20952 = ~new_n20947 & new_n20951 ;
  assign new_n20953 = new_n13928 & ~new_n20952 ;
  assign new_n20954 = ~new_n20938 & ~new_n20953 ;
  assign new_n20955 = lo0044 & ~new_n2249 ;
  assign new_n20956 = new_n15207 & new_n20955 ;
  assign new_n20957 = lo0918 & ~new_n20956 ;
  assign new_n20958 = lo1444 & new_n20956 ;
  assign new_n20959 = ~new_n20957 & ~new_n20958 ;
  assign new_n20960 = lo0919 & ~new_n20956 ;
  assign new_n20961 = lo1424 & new_n20956 ;
  assign new_n20962 = ~new_n20960 & ~new_n20961 ;
  assign new_n20963 = new_n2002 & new_n14668 ;
  assign new_n20964 = lo0920 & ~new_n20963 ;
  assign new_n20965 = lo1061 & new_n20963 ;
  assign new_n20966 = ~new_n20964 & ~new_n20965 ;
  assign new_n20967 = lo0921 & ~new_n20956 ;
  assign new_n20968 = lo1061 & new_n20956 ;
  assign new_n20969 = ~new_n20967 & ~new_n20968 ;
  assign new_n20970 = lo0922 & ~new_n20956 ;
  assign new_n20971 = lo1279 & new_n20956 ;
  assign new_n20972 = ~new_n20970 & ~new_n20971 ;
  assign new_n20973 = ~lo0052 & new_n14677 ;
  assign new_n20974 = lo0053 & new_n20973 ;
  assign new_n20975 = lo0923 & ~new_n20974 ;
  assign new_n20976 = lo1077 & new_n20974 ;
  assign new_n20977 = ~new_n20975 & ~new_n20976 ;
  assign new_n20978 = lo0052 & new_n14677 ;
  assign new_n20979 = ~lo0053 & new_n20978 ;
  assign new_n20980 = lo0924 & ~new_n20979 ;
  assign new_n20981 = lo1077 & new_n20979 ;
  assign new_n20982 = ~new_n20980 & ~new_n20981 ;
  assign new_n20983 = ~lo0053 & new_n20973 ;
  assign new_n20984 = lo0925 & ~new_n20983 ;
  assign new_n20985 = lo1077 & new_n20983 ;
  assign new_n20986 = ~new_n20984 & ~new_n20985 ;
  assign new_n20987 = lo0053 & new_n20978 ;
  assign new_n20988 = lo0926 & ~new_n20987 ;
  assign new_n20989 = lo1077 & new_n20987 ;
  assign new_n20990 = ~new_n20988 & ~new_n20989 ;
  assign new_n20991 = lo0927 & ~new_n20956 ;
  assign new_n20992 = lo1269 & new_n20956 ;
  assign new_n20993 = ~new_n20991 & ~new_n20992 ;
  assign new_n20994 = lo0928 & ~new_n20963 ;
  assign new_n20995 = lo1078 & new_n20963 ;
  assign new_n20996 = ~new_n20994 & ~new_n20995 ;
  assign new_n20997 = lo0929 & ~new_n20956 ;
  assign new_n20998 = lo1078 & new_n20956 ;
  assign new_n20999 = ~new_n20997 & ~new_n20998 ;
  assign new_n21000 = lo0930 & ~new_n16687 ;
  assign new_n21001 = lo1078 & new_n16687 ;
  assign new_n21002 = ~new_n21000 & ~new_n21001 ;
  assign new_n21003 = lo0931 & new_n2252 ;
  assign new_n21004 = ~new_n2252 & new_n13812 ;
  assign new_n21005 = new_n15451 & new_n21004 ;
  assign new_n21006 = ~new_n21003 & ~new_n21005 ;
  assign new_n21007 = lo0932 & new_n2252 ;
  assign new_n21008 = new_n2264 & new_n12789 ;
  assign new_n21009 = new_n12698 & new_n21008 ;
  assign new_n21010 = new_n12509 & new_n12761 ;
  assign new_n21011 = ~new_n12329 & new_n12460 ;
  assign new_n21012 = new_n21010 & new_n21011 ;
  assign new_n21013 = new_n12329 & new_n13768 ;
  assign new_n21014 = ~new_n21012 & ~new_n21013 ;
  assign new_n21015 = new_n12467 & new_n13807 ;
  assign new_n21016 = ~new_n21014 & new_n21015 ;
  assign new_n21017 = ~new_n21009 & ~new_n21016 ;
  assign new_n21018 = ~new_n2252 & ~new_n21017 ;
  assign new_n21019 = new_n15451 & new_n21018 ;
  assign new_n21020 = ~new_n21007 & ~new_n21019 ;
  assign new_n21021 = ~lo0887 & ~lo0933 ;
  assign new_n21022 = ~new_n13842 & ~new_n21021 ;
  assign new_n21023 = ~lo0888 & ~lo0934 ;
  assign new_n21024 = ~new_n13842 & ~new_n21023 ;
  assign new_n21025 = ~lo0889 & ~lo0935 ;
  assign new_n21026 = ~new_n13842 & ~new_n21025 ;
  assign new_n21027 = ~lo0890 & ~lo0936 ;
  assign new_n21028 = ~new_n13842 & ~new_n21027 ;
  assign new_n21029 = ~lo0891 & ~lo0937 ;
  assign new_n21030 = ~new_n13842 & ~new_n21029 ;
  assign new_n21031 = lo0944 & lo0947 ;
  assign new_n21032 = new_n20793 & new_n21031 ;
  assign new_n21033 = new_n20803 & ~new_n21032 ;
  assign new_n21034 = lo0945 & lo0947 ;
  assign new_n21035 = ~lo0946 & new_n21034 ;
  assign new_n21036 = ~lo0947 & new_n20793 ;
  assign new_n21037 = ~new_n21035 & ~new_n21036 ;
  assign new_n21038 = new_n21033 & new_n21037 ;
  assign new_n21039 = lo0944 & new_n20793 ;
  assign new_n21040 = ~new_n20803 & ~new_n21039 ;
  assign new_n21041 = ~lo0947 & ~lo0948 ;
  assign new_n21042 = lo0947 & lo0959 ;
  assign new_n21043 = ~new_n21041 & ~new_n21042 ;
  assign new_n21044 = ~new_n21040 & new_n21043 ;
  assign new_n21045 = ~new_n21038 & new_n21044 ;
  assign new_n21046 = new_n20795 & new_n21045 ;
  assign new_n21047 = new_n13842 & ~new_n21046 ;
  assign new_n21048 = lo0947 & new_n20798 ;
  assign new_n21049 = ~lo0948 & ~lo0959 ;
  assign new_n21050 = new_n21048 & new_n21049 ;
  assign new_n21051 = new_n20803 & new_n21048 ;
  assign new_n21052 = lo1068 & new_n20801 ;
  assign new_n21053 = lo0942 & new_n2252 ;
  assign new_n21054 = new_n12508 & ~new_n20769 ;
  assign new_n21055 = new_n15451 & new_n21054 ;
  assign new_n21056 = ~lo1079 & ~new_n21055 ;
  assign new_n21057 = ~new_n2252 & ~new_n21056 ;
  assign new_n21058 = ~new_n21053 & ~new_n21057 ;
  assign new_n21059 = lo0943 & new_n2252 ;
  assign new_n21060 = ~new_n12452 & new_n20771 ;
  assign new_n21061 = ~lo1080 & ~new_n21060 ;
  assign new_n21062 = ~new_n2252 & ~new_n21061 ;
  assign new_n21063 = ~new_n21059 & ~new_n21062 ;
  assign new_n21064 = lo0944 & new_n2252 ;
  assign new_n21065 = ~new_n12420 & new_n20771 ;
  assign new_n21066 = ~lo1081 & ~new_n21065 ;
  assign new_n21067 = ~new_n2252 & ~new_n21066 ;
  assign new_n21068 = ~new_n21064 & ~new_n21067 ;
  assign new_n21069 = lo0945 & new_n2252 ;
  assign new_n21070 = new_n15361 & new_n20771 ;
  assign new_n21071 = ~new_n21069 & ~new_n21070 ;
  assign new_n21072 = lo0946 & new_n2252 ;
  assign new_n21073 = ~new_n12441 & new_n20771 ;
  assign new_n21074 = ~lo1082 & ~new_n21073 ;
  assign new_n21075 = ~new_n2252 & ~new_n21074 ;
  assign new_n21076 = ~new_n21072 & ~new_n21075 ;
  assign new_n21077 = lo0947 & new_n2252 ;
  assign new_n21078 = new_n20520 & new_n20771 ;
  assign new_n21079 = ~new_n21077 & ~new_n21078 ;
  assign new_n21080 = lo0948 & new_n2252 ;
  assign new_n21081 = ~new_n12429 & new_n20771 ;
  assign new_n21082 = ~lo1083 & ~new_n21081 ;
  assign new_n21083 = ~new_n2252 & ~new_n21082 ;
  assign new_n21084 = ~new_n21080 & ~new_n21083 ;
  assign new_n21085 = lo0949 & new_n2252 ;
  assign new_n21086 = lo1084 & ~new_n2252 ;
  assign new_n21087 = ~new_n21085 & ~new_n21086 ;
  assign new_n21088 = lo0950 & new_n2252 ;
  assign new_n21089 = new_n13810 & new_n17339 ;
  assign new_n21090 = new_n14732 & new_n21089 ;
  assign new_n21091 = ~new_n21088 & ~new_n21090 ;
  assign new_n21092 = lo0951 & new_n2252 ;
  assign new_n21093 = ~new_n12329 & new_n13810 ;
  assign new_n21094 = new_n12524 & new_n13046 ;
  assign new_n21095 = ~new_n21093 & ~new_n21094 ;
  assign new_n21096 = new_n20585 & ~new_n21095 ;
  assign new_n21097 = ~new_n13043 & ~new_n13740 ;
  assign new_n21098 = new_n21096 & ~new_n21097 ;
  assign new_n21099 = ~lo1085 & ~new_n21098 ;
  assign new_n21100 = ~new_n2252 & ~new_n21099 ;
  assign new_n21101 = ~new_n21092 & ~new_n21100 ;
  assign new_n21102 = lo0952 & new_n2252 ;
  assign new_n21103 = new_n14732 & new_n20604 ;
  assign new_n21104 = ~new_n21102 & ~new_n21103 ;
  assign new_n21105 = lo0953 & new_n2252 ;
  assign new_n21106 = lo1086 & ~new_n2252 ;
  assign new_n21107 = ~new_n21105 & ~new_n21106 ;
  assign new_n21108 = lo0954 & new_n2252 ;
  assign new_n21109 = new_n12420 & new_n12460 ;
  assign new_n21110 = ~new_n12509 & ~new_n21109 ;
  assign new_n21111 = ~new_n2252 & ~new_n21110 ;
  assign new_n21112 = new_n17340 & new_n21111 ;
  assign new_n21113 = ~new_n21108 & ~new_n21112 ;
  assign new_n21114 = lo0955 & new_n2252 ;
  assign new_n21115 = ~new_n12467 & new_n13807 ;
  assign new_n21116 = new_n20603 & new_n21115 ;
  assign new_n21117 = new_n12402 & new_n13862 ;
  assign new_n21118 = new_n17099 & new_n21117 ;
  assign new_n21119 = ~new_n21116 & ~new_n21118 ;
  assign new_n21120 = ~new_n2252 & ~new_n21119 ;
  assign new_n21121 = new_n17045 & new_n21120 ;
  assign new_n21122 = ~new_n21114 & ~new_n21121 ;
  assign new_n21123 = lo0956 & new_n2252 ;
  assign new_n21124 = lo1087 & ~new_n2252 ;
  assign new_n21125 = ~new_n21123 & ~new_n21124 ;
  assign new_n21126 = lo0957 & new_n2252 ;
  assign new_n21127 = ~lo0870 & ~new_n2265 ;
  assign new_n21128 = new_n2265 & ~new_n12465 ;
  assign new_n21129 = ~new_n21127 & ~new_n21128 ;
  assign new_n21130 = new_n16908 & ~new_n21129 ;
  assign new_n21131 = new_n12549 & new_n21130 ;
  assign new_n21132 = new_n20586 & new_n21131 ;
  assign new_n21133 = ~new_n21126 & ~new_n21132 ;
  assign new_n21134 = lo0958 & new_n2252 ;
  assign new_n21135 = ~new_n12316 & new_n12507 ;
  assign new_n21136 = ~new_n12420 & new_n12838 ;
  assign new_n21137 = new_n2264 & new_n12420 ;
  assign new_n21138 = ~new_n21136 & ~new_n21137 ;
  assign new_n21139 = new_n12452 & new_n12508 ;
  assign new_n21140 = new_n12442 & new_n21139 ;
  assign new_n21141 = ~new_n21138 & new_n21140 ;
  assign new_n21142 = new_n2446 & new_n21012 ;
  assign new_n21143 = ~new_n12522 & ~new_n21142 ;
  assign new_n21144 = ~new_n21141 & new_n21143 ;
  assign new_n21145 = new_n2446 & ~new_n21144 ;
  assign new_n21146 = ~new_n21135 & new_n21145 ;
  assign new_n21147 = ~new_n2446 & new_n21144 ;
  assign new_n21148 = ~new_n21145 & ~new_n21147 ;
  assign new_n21149 = new_n21135 & ~new_n21148 ;
  assign new_n21150 = ~new_n2446 & new_n12860 ;
  assign new_n21151 = new_n12369 & new_n21150 ;
  assign new_n21152 = ~new_n21144 & new_n21151 ;
  assign new_n21153 = ~new_n21149 & ~new_n21152 ;
  assign new_n21154 = ~new_n21146 & new_n21153 ;
  assign new_n21155 = new_n2455 & ~new_n21154 ;
  assign new_n21156 = new_n2454 & new_n15442 ;
  assign new_n21157 = ~lo1291 & ~lo1293 ;
  assign new_n21158 = ~new_n13430 & ~new_n21157 ;
  assign new_n21159 = ~lo1292 & lo1294 ;
  assign new_n21160 = ~lo1292 & ~new_n21159 ;
  assign new_n21161 = ~new_n21158 & ~new_n21160 ;
  assign new_n21162 = new_n12912 & ~new_n21161 ;
  assign new_n21163 = new_n12357 & ~new_n21162 ;
  assign new_n21164 = lo1292 & lo1293 ;
  assign new_n21165 = ~new_n12811 & ~new_n21164 ;
  assign new_n21166 = ~new_n12791 & ~new_n21165 ;
  assign new_n21167 = new_n12576 & ~new_n21166 ;
  assign new_n21168 = ~new_n12357 & ~new_n21167 ;
  assign new_n21169 = new_n12325 & ~new_n21168 ;
  assign new_n21170 = ~new_n21163 & new_n21169 ;
  assign new_n21171 = new_n12658 & new_n12860 ;
  assign new_n21172 = ~new_n12658 & new_n21167 ;
  assign new_n21173 = ~new_n21171 & ~new_n21172 ;
  assign new_n21174 = ~new_n12325 & ~new_n21173 ;
  assign new_n21175 = ~new_n21170 & ~new_n21174 ;
  assign new_n21176 = ~new_n12329 & ~new_n21175 ;
  assign new_n21177 = ~new_n12547 & ~new_n21176 ;
  assign new_n21178 = new_n12789 & ~new_n21177 ;
  assign new_n21179 = ~new_n21156 & ~new_n21178 ;
  assign new_n21180 = ~new_n2450 & ~new_n21179 ;
  assign new_n21181 = ~new_n21155 & ~new_n21180 ;
  assign new_n21182 = ~new_n2252 & ~new_n21181 ;
  assign new_n21183 = new_n15451 & new_n21182 ;
  assign new_n21184 = ~new_n21134 & ~new_n21183 ;
  assign new_n21185 = lo0959 & new_n2252 ;
  assign new_n21186 = lo1088 & ~new_n2252 ;
  assign new_n21187 = ~new_n21185 & ~new_n21186 ;
  assign new_n21188 = lo0960 & new_n2252 ;
  assign new_n21189 = lo1089 & ~new_n2252 ;
  assign new_n21190 = ~new_n21188 & ~new_n21189 ;
  assign new_n21191 = lo0961 & new_n2252 ;
  assign new_n21192 = new_n14806 & new_n21089 ;
  assign new_n21193 = ~new_n21191 & ~new_n21192 ;
  assign new_n21194 = lo0962 & new_n2252 ;
  assign new_n21195 = ~new_n12329 & new_n12468 ;
  assign new_n21196 = ~new_n13740 & ~new_n21195 ;
  assign new_n21197 = new_n21096 & ~new_n21196 ;
  assign new_n21198 = ~lo1090 & ~new_n21197 ;
  assign new_n21199 = ~new_n2252 & ~new_n21198 ;
  assign new_n21200 = ~new_n21194 & ~new_n21199 ;
  assign new_n21201 = ~new_n2252 & new_n13916 ;
  assign new_n21202 = lo0963 & ~new_n21201 ;
  assign new_n21203 = ~new_n15196 & new_n21201 ;
  assign new_n21204 = ~new_n21202 & ~new_n21203 ;
  assign new_n21205 = lo0964 & ~new_n21201 ;
  assign new_n21206 = ~new_n15696 & new_n21201 ;
  assign new_n21207 = ~new_n21205 & ~new_n21206 ;
  assign new_n21208 = lo0965 & ~new_n20956 ;
  assign new_n21209 = lo1275 & new_n20956 ;
  assign new_n21210 = ~new_n21208 & ~new_n21209 ;
  assign new_n21211 = lo0966 & ~new_n20974 ;
  assign new_n21212 = lo1091 & new_n20974 ;
  assign new_n21213 = ~new_n21211 & ~new_n21212 ;
  assign new_n21214 = lo0967 & ~new_n20979 ;
  assign new_n21215 = lo1091 & new_n20979 ;
  assign new_n21216 = ~new_n21214 & ~new_n21215 ;
  assign new_n21217 = lo0968 & ~new_n20983 ;
  assign new_n21218 = lo1091 & new_n20983 ;
  assign new_n21219 = ~new_n21217 & ~new_n21218 ;
  assign new_n21220 = lo0969 & ~new_n20987 ;
  assign new_n21221 = lo1091 & new_n20987 ;
  assign new_n21222 = ~new_n21220 & ~new_n21221 ;
  assign new_n21223 = lo0970 & ~new_n20956 ;
  assign new_n21224 = lo1283 & new_n20956 ;
  assign new_n21225 = ~new_n21223 & ~new_n21224 ;
  assign new_n21226 = lo0971 & ~new_n20934 ;
  assign new_n21227 = lo1283 & new_n20934 ;
  assign new_n21228 = ~new_n21226 & ~new_n21227 ;
  assign new_n21229 = lo0972 & ~new_n21201 ;
  assign new_n21230 = ~new_n15749 & new_n21201 ;
  assign new_n21231 = ~new_n21229 & ~new_n21230 ;
  assign new_n21232 = lo0973 & ~new_n20956 ;
  assign new_n21233 = lo1423 & new_n20956 ;
  assign new_n21234 = ~new_n21232 & ~new_n21233 ;
  assign new_n21235 = lo0974 & ~new_n20963 ;
  assign new_n21236 = lo1055 & new_n20963 ;
  assign new_n21237 = ~new_n21235 & ~new_n21236 ;
  assign new_n21238 = lo0975 & ~new_n20956 ;
  assign new_n21239 = lo1055 & new_n20956 ;
  assign new_n21240 = ~new_n21238 & ~new_n21239 ;
  assign new_n21241 = lo0976 & ~new_n21201 ;
  assign new_n21242 = ~new_n15807 & new_n21201 ;
  assign new_n21243 = ~new_n21241 & ~new_n21242 ;
  assign new_n21244 = lo0980 & new_n14656 ;
  assign new_n21245 = lo0977 & ~new_n21244 ;
  assign new_n21246 = ~lo0977 & new_n21244 ;
  assign new_n21247 = ~new_n21245 & ~new_n21246 ;
  assign new_n21248 = new_n2011 & new_n14668 ;
  assign new_n21249 = lo1092 & ~new_n21248 ;
  assign new_n21250 = lo0978 & ~new_n21249 ;
  assign new_n21251 = lo0978 & ~lo0979 ;
  assign new_n21252 = ~lo0978 & lo0979 ;
  assign new_n21253 = ~new_n21251 & ~new_n21252 ;
  assign new_n21254 = new_n21249 & ~new_n21253 ;
  assign new_n21255 = ~new_n21250 & ~new_n21254 ;
  assign new_n21256 = lo0979 & ~new_n21249 ;
  assign new_n21257 = ~lo0979 & new_n21249 ;
  assign new_n21258 = ~new_n21256 & ~new_n21257 ;
  assign new_n21259 = ~lo0980 & ~new_n14656 ;
  assign new_n21260 = ~new_n21244 & ~new_n21259 ;
  assign new_n21261 = lo0981 & ~new_n20956 ;
  assign new_n21262 = lo1270 & new_n20956 ;
  assign new_n21263 = ~new_n21261 & ~new_n21262 ;
  assign new_n21264 = lo0982 & ~new_n20963 ;
  assign new_n21265 = lo1093 & new_n20963 ;
  assign new_n21266 = ~new_n21264 & ~new_n21265 ;
  assign new_n21267 = lo0983 & ~new_n20956 ;
  assign new_n21268 = lo1093 & new_n20956 ;
  assign new_n21269 = ~new_n21267 & ~new_n21268 ;
  assign new_n21270 = lo0984 & ~new_n16687 ;
  assign new_n21271 = lo1093 & new_n16687 ;
  assign new_n21272 = ~new_n21270 & ~new_n21271 ;
  assign new_n21273 = lo0985 & ~new_n21201 ;
  assign new_n21274 = ~new_n15858 & new_n21201 ;
  assign new_n21275 = ~new_n21273 & ~new_n21274 ;
  assign new_n21276 = lo0986 & ~new_n20956 ;
  assign new_n21277 = lo1420 & new_n20956 ;
  assign new_n21278 = ~new_n21276 & ~new_n21277 ;
  assign new_n21279 = lo0987 & ~new_n20963 ;
  assign new_n21280 = lo1053 & new_n20963 ;
  assign new_n21281 = ~new_n21279 & ~new_n21280 ;
  assign new_n21282 = lo0988 & ~new_n20956 ;
  assign new_n21283 = lo1053 & new_n20956 ;
  assign new_n21284 = ~new_n21282 & ~new_n21283 ;
  assign new_n21285 = lo0989 & ~new_n21201 ;
  assign new_n21286 = ~new_n15906 & new_n21201 ;
  assign new_n21287 = ~new_n21285 & ~new_n21286 ;
  assign new_n21288 = lo0990 & ~new_n20956 ;
  assign new_n21289 = lo1271 & new_n20956 ;
  assign new_n21290 = ~new_n21288 & ~new_n21289 ;
  assign new_n21291 = lo0991 & ~new_n20963 ;
  assign new_n21292 = lo1094 & new_n20963 ;
  assign new_n21293 = ~new_n21291 & ~new_n21292 ;
  assign new_n21294 = lo0992 & ~new_n20956 ;
  assign new_n21295 = lo1094 & new_n20956 ;
  assign new_n21296 = ~new_n21294 & ~new_n21295 ;
  assign new_n21297 = lo0993 & ~new_n21201 ;
  assign new_n21298 = ~new_n15973 & new_n21201 ;
  assign new_n21299 = ~new_n21297 & ~new_n21298 ;
  assign new_n21300 = lo0994 & ~new_n20956 ;
  assign new_n21301 = lo1277 & new_n20956 ;
  assign new_n21302 = ~new_n21300 & ~new_n21301 ;
  assign new_n21303 = lo0995 & ~new_n20979 ;
  assign new_n21304 = lo1095 & new_n20979 ;
  assign new_n21305 = ~new_n21303 & ~new_n21304 ;
  assign new_n21306 = lo0996 & ~new_n20974 ;
  assign new_n21307 = lo1095 & new_n20974 ;
  assign new_n21308 = ~new_n21306 & ~new_n21307 ;
  assign new_n21309 = lo0997 & ~new_n20983 ;
  assign new_n21310 = lo1095 & new_n20983 ;
  assign new_n21311 = ~new_n21309 & ~new_n21310 ;
  assign new_n21312 = lo0998 & ~new_n20987 ;
  assign new_n21313 = lo1095 & new_n20987 ;
  assign new_n21314 = ~new_n21312 & ~new_n21313 ;
  assign new_n21315 = lo0999 & ~new_n20934 ;
  assign new_n21316 = lo1446 & new_n20934 ;
  assign new_n21317 = ~new_n21315 & ~new_n21316 ;
  assign new_n21318 = lo1000 & ~new_n20956 ;
  assign new_n21319 = lo1446 & new_n20956 ;
  assign new_n21320 = ~new_n21318 & ~new_n21319 ;
  assign new_n21321 = lo1001 & ~new_n21201 ;
  assign new_n21322 = ~new_n15288 & new_n21201 ;
  assign new_n21323 = ~new_n21321 & ~new_n21322 ;
  assign new_n21324 = lo1002 & ~new_n21201 ;
  assign new_n21325 = ~new_n16052 & new_n21201 ;
  assign new_n21326 = ~new_n21324 & ~new_n21325 ;
  assign new_n21327 = lo1003 & ~new_n20956 ;
  assign new_n21328 = lo1274 & new_n20956 ;
  assign new_n21329 = ~new_n21327 & ~new_n21328 ;
  assign new_n21330 = lo1004 & ~new_n20974 ;
  assign new_n21331 = lo1096 & new_n20974 ;
  assign new_n21332 = ~new_n21330 & ~new_n21331 ;
  assign new_n21333 = lo1005 & ~new_n20979 ;
  assign new_n21334 = lo1096 & new_n20979 ;
  assign new_n21335 = ~new_n21333 & ~new_n21334 ;
  assign new_n21336 = lo1006 & ~new_n20983 ;
  assign new_n21337 = lo1096 & new_n20983 ;
  assign new_n21338 = ~new_n21336 & ~new_n21337 ;
  assign new_n21339 = lo1007 & ~new_n20987 ;
  assign new_n21340 = lo1096 & new_n20987 ;
  assign new_n21341 = ~new_n21339 & ~new_n21340 ;
  assign new_n21342 = lo1008 & ~new_n20956 ;
  assign new_n21343 = lo1282 & new_n20956 ;
  assign new_n21344 = ~new_n21342 & ~new_n21343 ;
  assign new_n21345 = lo1009 & ~new_n20934 ;
  assign new_n21346 = lo1282 & new_n20934 ;
  assign new_n21347 = ~new_n21345 & ~new_n21346 ;
  assign new_n21348 = lo1010 & ~new_n21201 ;
  assign new_n21349 = ~new_n16105 & new_n21201 ;
  assign new_n21350 = ~new_n21348 & ~new_n21349 ;
  assign new_n21351 = lo1011 & ~new_n20956 ;
  assign new_n21352 = lo1422 & new_n20956 ;
  assign new_n21353 = ~new_n21351 & ~new_n21352 ;
  assign new_n21354 = lo1012 & ~new_n20963 ;
  assign new_n21355 = lo1052 & new_n20963 ;
  assign new_n21356 = ~new_n21354 & ~new_n21355 ;
  assign new_n21357 = lo1013 & ~new_n20956 ;
  assign new_n21358 = lo1052 & new_n20956 ;
  assign new_n21359 = ~new_n21357 & ~new_n21358 ;
  assign new_n21360 = lo1014 & ~new_n21201 ;
  assign new_n21361 = ~new_n16153 & new_n21201 ;
  assign new_n21362 = ~new_n21360 & ~new_n21361 ;
  assign new_n21363 = lo1015 & ~new_n20956 ;
  assign new_n21364 = lo1421 & new_n20956 ;
  assign new_n21365 = ~new_n21363 & ~new_n21364 ;
  assign new_n21366 = lo1016 & ~new_n20963 ;
  assign new_n21367 = lo1054 & new_n20963 ;
  assign new_n21368 = ~new_n21366 & ~new_n21367 ;
  assign new_n21369 = lo1017 & ~new_n20956 ;
  assign new_n21370 = lo1054 & new_n20956 ;
  assign new_n21371 = ~new_n21369 & ~new_n21370 ;
  assign new_n21372 = lo1018 & ~new_n21201 ;
  assign new_n21373 = ~new_n15262 & new_n21201 ;
  assign new_n21374 = ~new_n21372 & ~new_n21373 ;
  assign new_n21375 = lo1019 & ~new_n21201 ;
  assign new_n21376 = ~new_n16229 & new_n21201 ;
  assign new_n21377 = ~new_n21375 & ~new_n21376 ;
  assign new_n21378 = lo1020 & ~new_n20956 ;
  assign new_n21379 = lo1278 & new_n20956 ;
  assign new_n21380 = ~new_n21378 & ~new_n21379 ;
  assign new_n21381 = lo1021 & ~new_n20979 ;
  assign new_n21382 = lo1097 & new_n20979 ;
  assign new_n21383 = ~new_n21381 & ~new_n21382 ;
  assign new_n21384 = lo1022 & ~new_n20974 ;
  assign new_n21385 = lo1097 & new_n20974 ;
  assign new_n21386 = ~new_n21384 & ~new_n21385 ;
  assign new_n21387 = lo1023 & ~new_n20983 ;
  assign new_n21388 = lo1097 & new_n20983 ;
  assign new_n21389 = ~new_n21387 & ~new_n21388 ;
  assign new_n21390 = lo1024 & ~new_n20987 ;
  assign new_n21391 = lo1097 & new_n20987 ;
  assign new_n21392 = ~new_n21390 & ~new_n21391 ;
  assign new_n21393 = lo1025 & ~new_n20934 ;
  assign new_n21394 = lo1445 & new_n20934 ;
  assign new_n21395 = ~new_n21393 & ~new_n21394 ;
  assign new_n21396 = lo1026 & ~new_n20956 ;
  assign new_n21397 = lo1445 & new_n20956 ;
  assign new_n21398 = ~new_n21396 & ~new_n21397 ;
  assign new_n21399 = lo1027 & ~new_n21201 ;
  assign new_n21400 = ~new_n16299 & new_n21201 ;
  assign new_n21401 = ~new_n21399 & ~new_n21400 ;
  assign new_n21402 = lo1028 & ~new_n20956 ;
  assign new_n21403 = lo1273 & new_n20956 ;
  assign new_n21404 = ~new_n21402 & ~new_n21403 ;
  assign new_n21405 = lo1029 & ~new_n20979 ;
  assign new_n21406 = lo1098 & new_n20979 ;
  assign new_n21407 = ~new_n21405 & ~new_n21406 ;
  assign new_n21408 = lo1030 & ~new_n20974 ;
  assign new_n21409 = lo1098 & new_n20974 ;
  assign new_n21410 = ~new_n21408 & ~new_n21409 ;
  assign new_n21411 = lo1031 & ~new_n20983 ;
  assign new_n21412 = lo1098 & new_n20983 ;
  assign new_n21413 = ~new_n21411 & ~new_n21412 ;
  assign new_n21414 = lo1032 & ~new_n20987 ;
  assign new_n21415 = lo1098 & new_n20987 ;
  assign new_n21416 = ~new_n21414 & ~new_n21415 ;
  assign new_n21417 = lo1033 & ~new_n20956 ;
  assign new_n21418 = lo1281 & new_n20956 ;
  assign new_n21419 = ~new_n21417 & ~new_n21418 ;
  assign new_n21420 = lo1034 & ~new_n20934 ;
  assign new_n21421 = lo1281 & new_n20934 ;
  assign new_n21422 = ~new_n21420 & ~new_n21421 ;
  assign new_n21423 = lo1035 & ~new_n21201 ;
  assign new_n21424 = ~new_n16371 & new_n21201 ;
  assign new_n21425 = ~new_n21423 & ~new_n21424 ;
  assign new_n21426 = lo1036 & ~new_n20956 ;
  assign new_n21427 = lo1276 & new_n20956 ;
  assign new_n21428 = ~new_n21426 & ~new_n21427 ;
  assign new_n21429 = lo1037 & ~new_n20979 ;
  assign new_n21430 = lo1099 & new_n20979 ;
  assign new_n21431 = ~new_n21429 & ~new_n21430 ;
  assign new_n21432 = lo1038 & ~new_n20974 ;
  assign new_n21433 = lo1099 & new_n20974 ;
  assign new_n21434 = ~new_n21432 & ~new_n21433 ;
  assign new_n21435 = lo1039 & ~new_n20983 ;
  assign new_n21436 = lo1099 & new_n20983 ;
  assign new_n21437 = ~new_n21435 & ~new_n21436 ;
  assign new_n21438 = lo1040 & ~new_n20987 ;
  assign new_n21439 = lo1099 & new_n20987 ;
  assign new_n21440 = ~new_n21438 & ~new_n21439 ;
  assign new_n21441 = lo1041 & ~new_n20956 ;
  assign new_n21442 = lo1284 & new_n20956 ;
  assign new_n21443 = ~new_n21441 & ~new_n21442 ;
  assign new_n21444 = lo1042 & ~new_n20934 ;
  assign new_n21445 = lo1284 & new_n20934 ;
  assign new_n21446 = ~new_n21444 & ~new_n21445 ;
  assign new_n21447 = lo1043 & ~new_n21201 ;
  assign new_n21448 = ~new_n16443 & new_n21201 ;
  assign new_n21449 = ~new_n21447 & ~new_n21448 ;
  assign new_n21450 = lo1044 & ~new_n20956 ;
  assign new_n21451 = lo1272 & new_n20956 ;
  assign new_n21452 = ~new_n21450 & ~new_n21451 ;
  assign new_n21453 = lo1045 & ~new_n20974 ;
  assign new_n21454 = lo1100 & new_n20974 ;
  assign new_n21455 = ~new_n21453 & ~new_n21454 ;
  assign new_n21456 = lo1046 & ~new_n20979 ;
  assign new_n21457 = lo1100 & new_n20979 ;
  assign new_n21458 = ~new_n21456 & ~new_n21457 ;
  assign new_n21459 = lo1047 & ~new_n20983 ;
  assign new_n21460 = lo1100 & new_n20983 ;
  assign new_n21461 = ~new_n21459 & ~new_n21460 ;
  assign new_n21462 = lo1048 & ~new_n20987 ;
  assign new_n21463 = lo1100 & new_n20987 ;
  assign new_n21464 = ~new_n21462 & ~new_n21463 ;
  assign new_n21465 = lo1049 & ~new_n20956 ;
  assign new_n21466 = lo1280 & new_n20956 ;
  assign new_n21467 = ~new_n21465 & ~new_n21466 ;
  assign new_n21468 = lo1050 & ~new_n20934 ;
  assign new_n21469 = lo1280 & new_n20934 ;
  assign new_n21470 = ~new_n21468 & ~new_n21469 ;
  assign new_n21471 = lo1051 & ~new_n13928 ;
  assign new_n21472 = ~new_n14609 & ~new_n14619 ;
  assign new_n21473 = new_n14607 & ~new_n21472 ;
  assign new_n21474 = ~new_n14610 & ~new_n21473 ;
  assign new_n21475 = ~new_n2261 & ~new_n21474 ;
  assign new_n21476 = ~new_n14643 & ~new_n21475 ;
  assign new_n21477 = new_n13928 & ~new_n21476 ;
  assign new_n21478 = ~new_n21471 & ~new_n21477 ;
  assign new_n21479 = lo1290 & new_n13928 ;
  assign new_n21480 = lo1052 & ~new_n21479 ;
  assign new_n21481 = lo0112 & lo0113 ;
  assign new_n21482 = ~new_n14609 & ~new_n21481 ;
  assign new_n21483 = lo0113 & new_n21482 ;
  assign new_n21484 = ~new_n14128 & new_n21483 ;
  assign new_n21485 = lo0113 & ~new_n21482 ;
  assign new_n21486 = lo0112 & new_n16716 ;
  assign new_n21487 = new_n16716 & ~new_n21486 ;
  assign new_n21488 = ~new_n8780 & ~new_n21487 ;
  assign new_n21489 = ~lo0112 & new_n8780 ;
  assign new_n21490 = ~new_n16716 & new_n21489 ;
  assign new_n21491 = ~new_n21488 & ~new_n21490 ;
  assign new_n21492 = ~lo0113 & ~new_n21491 ;
  assign new_n21493 = new_n21482 & new_n21492 ;
  assign new_n21494 = ~new_n21485 & ~new_n21493 ;
  assign new_n21495 = ~new_n21484 & new_n21494 ;
  assign new_n21496 = new_n21482 & ~new_n21495 ;
  assign new_n21497 = ~new_n21482 & new_n21495 ;
  assign new_n21498 = ~new_n21496 & ~new_n21497 ;
  assign new_n21499 = lo1469 & ~new_n21498 ;
  assign new_n21500 = ~lo1469 & new_n21496 ;
  assign new_n21501 = ~new_n4003 & ~new_n21482 ;
  assign new_n21502 = ~new_n21495 & new_n21501 ;
  assign new_n21503 = ~new_n21500 & ~new_n21502 ;
  assign new_n21504 = ~new_n21499 & new_n21503 ;
  assign new_n21505 = new_n21479 & ~new_n21504 ;
  assign new_n21506 = ~new_n21480 & ~new_n21505 ;
  assign new_n21507 = lo1053 & ~new_n21479 ;
  assign new_n21508 = ~new_n14181 & new_n21483 ;
  assign new_n21509 = lo0112 & new_n18863 ;
  assign new_n21510 = new_n18863 & ~new_n21509 ;
  assign new_n21511 = ~new_n9021 & ~new_n21510 ;
  assign new_n21512 = ~lo0112 & new_n9021 ;
  assign new_n21513 = ~new_n18863 & new_n21512 ;
  assign new_n21514 = ~new_n21511 & ~new_n21513 ;
  assign new_n21515 = ~lo0113 & ~new_n21514 ;
  assign new_n21516 = new_n21482 & new_n21515 ;
  assign new_n21517 = ~new_n21485 & ~new_n21516 ;
  assign new_n21518 = ~new_n21508 & new_n21517 ;
  assign new_n21519 = new_n21482 & ~new_n21518 ;
  assign new_n21520 = ~new_n21482 & new_n21518 ;
  assign new_n21521 = ~new_n21519 & ~new_n21520 ;
  assign new_n21522 = lo1470 & ~new_n21521 ;
  assign new_n21523 = ~lo1470 & new_n21519 ;
  assign new_n21524 = ~new_n4724 & ~new_n21482 ;
  assign new_n21525 = ~new_n21518 & new_n21524 ;
  assign new_n21526 = ~new_n21523 & ~new_n21525 ;
  assign new_n21527 = ~new_n21522 & new_n21526 ;
  assign new_n21528 = new_n21479 & ~new_n21527 ;
  assign new_n21529 = ~new_n21507 & ~new_n21528 ;
  assign new_n21530 = lo1054 & ~new_n21479 ;
  assign new_n21531 = ~new_n14154 & new_n21483 ;
  assign new_n21532 = lo0112 & new_n16735 ;
  assign new_n21533 = new_n16735 & ~new_n21532 ;
  assign new_n21534 = ~new_n8902 & ~new_n21533 ;
  assign new_n21535 = ~lo0112 & new_n8902 ;
  assign new_n21536 = ~new_n16735 & new_n21535 ;
  assign new_n21537 = ~new_n21534 & ~new_n21536 ;
  assign new_n21538 = ~lo0113 & ~new_n21537 ;
  assign new_n21539 = new_n21482 & new_n21538 ;
  assign new_n21540 = ~new_n21485 & ~new_n21539 ;
  assign new_n21541 = ~new_n21531 & new_n21540 ;
  assign new_n21542 = new_n21482 & ~new_n21541 ;
  assign new_n21543 = ~new_n21482 & new_n21541 ;
  assign new_n21544 = ~new_n21542 & ~new_n21543 ;
  assign new_n21545 = lo1471 & ~new_n21544 ;
  assign new_n21546 = ~lo1471 & new_n21542 ;
  assign new_n21547 = ~new_n4362 & ~new_n21482 ;
  assign new_n21548 = ~new_n21541 & new_n21547 ;
  assign new_n21549 = ~new_n21546 & ~new_n21548 ;
  assign new_n21550 = ~new_n21545 & new_n21549 ;
  assign new_n21551 = new_n21479 & ~new_n21550 ;
  assign new_n21552 = ~new_n21530 & ~new_n21551 ;
  assign new_n21553 = lo1055 & ~new_n21479 ;
  assign new_n21554 = ~new_n14101 & new_n21483 ;
  assign new_n21555 = lo0112 & new_n16697 ;
  assign new_n21556 = new_n16697 & ~new_n21555 ;
  assign new_n21557 = ~new_n8659 & ~new_n21556 ;
  assign new_n21558 = ~lo0112 & new_n8659 ;
  assign new_n21559 = ~new_n16697 & new_n21558 ;
  assign new_n21560 = ~new_n21557 & ~new_n21559 ;
  assign new_n21561 = ~lo0113 & ~new_n21560 ;
  assign new_n21562 = new_n21482 & new_n21561 ;
  assign new_n21563 = ~new_n21485 & ~new_n21562 ;
  assign new_n21564 = ~new_n21554 & new_n21563 ;
  assign new_n21565 = new_n21482 & ~new_n21564 ;
  assign new_n21566 = ~new_n21482 & new_n21564 ;
  assign new_n21567 = ~new_n21565 & ~new_n21566 ;
  assign new_n21568 = lo1472 & ~new_n21567 ;
  assign new_n21569 = ~lo1472 & new_n21565 ;
  assign new_n21570 = ~new_n3639 & ~new_n21482 ;
  assign new_n21571 = ~new_n21564 & new_n21570 ;
  assign new_n21572 = ~new_n21569 & ~new_n21571 ;
  assign new_n21573 = ~new_n21568 & new_n21572 ;
  assign new_n21574 = new_n21479 & ~new_n21573 ;
  assign new_n21575 = ~new_n21553 & ~new_n21574 ;
  assign new_n21576 = lo1056 & ~new_n13928 ;
  assign new_n21577 = new_n13978 & ~new_n16735 ;
  assign new_n21578 = ~new_n13937 & ~new_n16920 ;
  assign new_n21579 = new_n13943 & new_n21578 ;
  assign new_n21580 = ~new_n13955 & ~new_n21579 ;
  assign new_n21581 = ~new_n21577 & new_n21580 ;
  assign new_n21582 = ~new_n13937 & ~new_n21581 ;
  assign new_n21583 = new_n13937 & new_n21581 ;
  assign new_n21584 = ~new_n21582 & ~new_n21583 ;
  assign new_n21585 = ~new_n6461 & ~new_n21584 ;
  assign new_n21586 = new_n6461 & new_n21582 ;
  assign new_n21587 = lo0321 & new_n13937 ;
  assign new_n21588 = ~new_n21581 & new_n21587 ;
  assign new_n21589 = ~new_n21586 & ~new_n21588 ;
  assign new_n21590 = ~new_n21585 & new_n21589 ;
  assign new_n21591 = new_n13928 & ~new_n21590 ;
  assign new_n21592 = ~new_n21576 & ~new_n21591 ;
  assign new_n21593 = lo1057 & ~new_n13928 ;
  assign new_n21594 = ~new_n13937 & ~new_n19091 ;
  assign new_n21595 = new_n13943 & new_n21594 ;
  assign new_n21596 = ~new_n6225 & new_n13937 ;
  assign new_n21597 = new_n13943 & new_n21596 ;
  assign new_n21598 = ~new_n13955 & ~new_n21597 ;
  assign new_n21599 = ~new_n21595 & new_n21598 ;
  assign new_n21600 = new_n13943 & ~new_n21599 ;
  assign new_n21601 = new_n16716 & new_n21600 ;
  assign new_n21602 = ~new_n13943 & new_n21599 ;
  assign new_n21603 = ~new_n21600 & ~new_n21602 ;
  assign new_n21604 = ~new_n16716 & ~new_n21603 ;
  assign new_n21605 = lo0601 & ~new_n13943 ;
  assign new_n21606 = ~new_n21599 & new_n21605 ;
  assign new_n21607 = ~new_n21604 & ~new_n21606 ;
  assign new_n21608 = ~new_n21601 & new_n21607 ;
  assign new_n21609 = new_n13928 & ~new_n21608 ;
  assign new_n21610 = ~new_n21593 & ~new_n21609 ;
  assign new_n21611 = lo1058 & ~new_n13928 ;
  assign new_n21612 = ~new_n13937 & ~new_n17933 ;
  assign new_n21613 = new_n13943 & new_n21612 ;
  assign new_n21614 = ~new_n5766 & new_n13937 ;
  assign new_n21615 = new_n13943 & new_n21614 ;
  assign new_n21616 = ~new_n13955 & ~new_n21615 ;
  assign new_n21617 = ~new_n21613 & new_n21616 ;
  assign new_n21618 = new_n13943 & ~new_n21617 ;
  assign new_n21619 = new_n16677 & new_n21618 ;
  assign new_n21620 = ~new_n13943 & new_n21617 ;
  assign new_n21621 = ~new_n21618 & ~new_n21620 ;
  assign new_n21622 = ~new_n16677 & ~new_n21621 ;
  assign new_n21623 = lo0559 & ~new_n13943 ;
  assign new_n21624 = ~new_n21617 & new_n21623 ;
  assign new_n21625 = ~new_n21622 & ~new_n21624 ;
  assign new_n21626 = ~new_n21619 & new_n21625 ;
  assign new_n21627 = new_n13928 & ~new_n21626 ;
  assign new_n21628 = ~new_n21611 & ~new_n21627 ;
  assign new_n21629 = lo1059 & ~new_n13928 ;
  assign new_n21630 = new_n13978 & ~new_n16697 ;
  assign new_n21631 = ~new_n13937 & ~new_n18614 ;
  assign new_n21632 = new_n13943 & new_n21631 ;
  assign new_n21633 = ~new_n13955 & ~new_n21632 ;
  assign new_n21634 = ~new_n21630 & new_n21633 ;
  assign new_n21635 = ~new_n13937 & ~new_n21634 ;
  assign new_n21636 = new_n13937 & new_n21634 ;
  assign new_n21637 = ~new_n21635 & ~new_n21636 ;
  assign new_n21638 = ~new_n5996 & ~new_n21637 ;
  assign new_n21639 = new_n5996 & new_n21635 ;
  assign new_n21640 = lo0517 & new_n13937 ;
  assign new_n21641 = ~new_n21634 & new_n21640 ;
  assign new_n21642 = ~new_n21639 & ~new_n21641 ;
  assign new_n21643 = ~new_n21638 & new_n21642 ;
  assign new_n21644 = new_n13928 & ~new_n21643 ;
  assign new_n21645 = ~new_n21629 & ~new_n21644 ;
  assign new_n21646 = lo1060 & ~new_n13928 ;
  assign new_n21647 = ~new_n13937 & ~new_n18974 ;
  assign new_n21648 = new_n13943 & new_n21647 ;
  assign new_n21649 = ~new_n6690 & new_n13937 ;
  assign new_n21650 = new_n13943 & new_n21649 ;
  assign new_n21651 = ~new_n13955 & ~new_n21650 ;
  assign new_n21652 = ~new_n21648 & new_n21651 ;
  assign new_n21653 = new_n13943 & ~new_n21652 ;
  assign new_n21654 = new_n18863 & new_n21653 ;
  assign new_n21655 = ~new_n13943 & new_n21652 ;
  assign new_n21656 = ~new_n21653 & ~new_n21655 ;
  assign new_n21657 = ~new_n18863 & ~new_n21656 ;
  assign new_n21658 = lo0581 & ~new_n13943 ;
  assign new_n21659 = ~new_n21652 & new_n21658 ;
  assign new_n21660 = ~new_n21657 & ~new_n21659 ;
  assign new_n21661 = ~new_n21654 & new_n21660 ;
  assign new_n21662 = new_n13928 & ~new_n21661 ;
  assign new_n21663 = ~new_n21646 & ~new_n21662 ;
  assign new_n21664 = lo1061 & ~new_n21479 ;
  assign new_n21665 = ~new_n14060 & new_n21483 ;
  assign new_n21666 = lo0112 & new_n16677 ;
  assign new_n21667 = new_n16677 & ~new_n21666 ;
  assign new_n21668 = ~new_n8533 & ~new_n21667 ;
  assign new_n21669 = ~lo0112 & new_n8533 ;
  assign new_n21670 = ~new_n16677 & new_n21669 ;
  assign new_n21671 = ~new_n21668 & ~new_n21670 ;
  assign new_n21672 = ~lo0113 & ~new_n21671 ;
  assign new_n21673 = new_n21482 & new_n21672 ;
  assign new_n21674 = ~new_n21485 & ~new_n21673 ;
  assign new_n21675 = ~new_n21665 & new_n21674 ;
  assign new_n21676 = new_n21482 & ~new_n21675 ;
  assign new_n21677 = ~new_n21482 & new_n21675 ;
  assign new_n21678 = ~new_n21676 & ~new_n21677 ;
  assign new_n21679 = lo1473 & ~new_n21678 ;
  assign new_n21680 = ~lo1473 & new_n21676 ;
  assign new_n21681 = ~new_n3281 & ~new_n21482 ;
  assign new_n21682 = ~new_n21675 & new_n21681 ;
  assign new_n21683 = ~new_n21680 & ~new_n21682 ;
  assign new_n21684 = ~new_n21679 & new_n21683 ;
  assign new_n21685 = new_n21479 & ~new_n21684 ;
  assign new_n21686 = ~new_n21664 & ~new_n21685 ;
  assign new_n21687 = new_n15611 & new_n16664 ;
  assign new_n21688 = lo1062 & ~new_n21687 ;
  assign new_n21689 = ~new_n2415 & new_n21687 ;
  assign new_n21690 = ~new_n21688 & ~new_n21689 ;
  assign new_n21691 = lo1063 & ~new_n21687 ;
  assign new_n21692 = ~new_n2417 & new_n21687 ;
  assign new_n21693 = ~new_n21691 & ~new_n21692 ;
  assign new_n21694 = lo1064 & ~new_n21687 ;
  assign new_n21695 = ~new_n2419 & new_n21687 ;
  assign new_n21696 = ~new_n21694 & ~new_n21695 ;
  assign new_n21697 = lo1065 & ~new_n21687 ;
  assign new_n21698 = ~new_n2422 & new_n21687 ;
  assign new_n21699 = ~new_n21697 & ~new_n21698 ;
  assign new_n21700 = lo1066 & new_n2252 ;
  assign new_n21701 = new_n12523 & new_n13807 ;
  assign new_n21702 = new_n21010 & new_n21701 ;
  assign new_n21703 = new_n2450 & new_n17075 ;
  assign new_n21704 = new_n12325 & new_n15526 ;
  assign new_n21705 = ~new_n12377 & ~new_n21704 ;
  assign new_n21706 = ~new_n2450 & ~new_n21705 ;
  assign new_n21707 = new_n12386 & new_n21706 ;
  assign new_n21708 = ~new_n21703 & ~new_n21707 ;
  assign new_n21709 = new_n14790 & ~new_n21708 ;
  assign new_n21710 = ~new_n21702 & ~new_n21709 ;
  assign new_n21711 = ~new_n2252 & ~new_n21710 ;
  assign new_n21712 = new_n17045 & new_n21711 ;
  assign new_n21713 = ~new_n21700 & ~new_n21712 ;
  assign new_n21714 = lo1067 & new_n2252 ;
  assign new_n21715 = lo1101 & ~new_n2252 ;
  assign new_n21716 = ~new_n21714 & ~new_n21715 ;
  assign new_n21717 = ~new_n12329 & new_n12720 ;
  assign new_n21718 = new_n12442 & new_n21717 ;
  assign new_n21719 = ~new_n20787 & ~new_n21718 ;
  assign new_n21720 = new_n12383 & new_n13807 ;
  assign new_n21721 = ~new_n21719 & new_n21720 ;
  assign new_n21722 = lo1384 & new_n21721 ;
  assign new_n21723 = lo1068 & ~new_n21721 ;
  assign new_n21724 = ~new_n21722 & ~new_n21723 ;
  assign new_n21725 = lo1069 & ~new_n20863 ;
  assign new_n21726 = lo1102 & ~new_n14656 ;
  assign new_n21727 = ~lo0980 & lo1105 ;
  assign new_n21728 = ~lo0977 & new_n21727 ;
  assign new_n21729 = ~lo0980 & lo1104 ;
  assign new_n21730 = lo0977 & new_n21729 ;
  assign new_n21731 = ~new_n20868 & ~new_n21730 ;
  assign new_n21732 = ~new_n21728 & new_n21731 ;
  assign new_n21733 = ~lo0980 & ~new_n21732 ;
  assign new_n21734 = lo0980 & new_n21732 ;
  assign new_n21735 = ~new_n21733 & ~new_n21734 ;
  assign new_n21736 = lo1103 & ~new_n21735 ;
  assign new_n21737 = ~lo1103 & new_n21733 ;
  assign new_n21738 = lo0980 & lo1106 ;
  assign new_n21739 = ~new_n21732 & new_n21738 ;
  assign new_n21740 = ~new_n21737 & ~new_n21739 ;
  assign new_n21741 = ~new_n21736 & new_n21740 ;
  assign new_n21742 = new_n14656 & ~new_n21741 ;
  assign new_n21743 = ~new_n21726 & ~new_n21742 ;
  assign new_n21744 = new_n20863 & ~new_n21743 ;
  assign new_n21745 = ~new_n21725 & ~new_n21744 ;
  assign new_n21746 = lo0978 & new_n21257 ;
  assign new_n21747 = lo1070 & ~new_n21746 ;
  assign new_n21748 = lo1107 & new_n21746 ;
  assign new_n21749 = ~new_n21747 & ~new_n21748 ;
  assign new_n21750 = lo0979 & new_n21249 ;
  assign new_n21751 = ~lo0978 & new_n21750 ;
  assign new_n21752 = lo1071 & ~new_n21751 ;
  assign new_n21753 = lo1107 & new_n21751 ;
  assign new_n21754 = ~new_n21752 & ~new_n21753 ;
  assign new_n21755 = ~lo0978 & new_n21257 ;
  assign new_n21756 = lo1072 & ~new_n21755 ;
  assign new_n21757 = lo1107 & new_n21755 ;
  assign new_n21758 = ~new_n21756 & ~new_n21757 ;
  assign new_n21759 = lo0978 & new_n21750 ;
  assign new_n21760 = lo1073 & ~new_n21759 ;
  assign new_n21761 = lo1107 & new_n21759 ;
  assign new_n21762 = ~new_n21760 & ~new_n21761 ;
  assign new_n21763 = lo1042 & ~lo1457 ;
  assign new_n21764 = ~lo1042 & lo1457 ;
  assign new_n21765 = ~new_n21763 & ~new_n21764 ;
  assign new_n21766 = lo1034 & ~lo1452 ;
  assign new_n21767 = ~lo0971 & lo1456 ;
  assign new_n21768 = ~new_n21766 & ~new_n21767 ;
  assign new_n21769 = new_n21765 & new_n21768 ;
  assign new_n21770 = lo1009 & ~lo1459 ;
  assign new_n21771 = ~lo1009 & lo1459 ;
  assign new_n21772 = ~new_n21770 & ~new_n21771 ;
  assign new_n21773 = lo1025 & ~lo1458 ;
  assign new_n21774 = ~lo1025 & lo1458 ;
  assign new_n21775 = ~new_n21773 & ~new_n21774 ;
  assign new_n21776 = new_n21772 & new_n21775 ;
  assign new_n21777 = new_n21769 & new_n21776 ;
  assign new_n21778 = lo0916 & ~lo1453 ;
  assign new_n21779 = ~lo0916 & lo1453 ;
  assign new_n21780 = ~new_n21778 & ~new_n21779 ;
  assign new_n21781 = ~lo1034 & lo1452 ;
  assign new_n21782 = lo0971 & ~lo1456 ;
  assign new_n21783 = ~new_n21781 & ~new_n21782 ;
  assign new_n21784 = new_n21780 & new_n21783 ;
  assign new_n21785 = lo0999 & ~lo1455 ;
  assign new_n21786 = ~lo0999 & lo1455 ;
  assign new_n21787 = ~new_n21785 & ~new_n21786 ;
  assign new_n21788 = lo1050 & ~lo1454 ;
  assign new_n21789 = ~lo1050 & lo1454 ;
  assign new_n21790 = ~new_n21788 & ~new_n21789 ;
  assign new_n21791 = new_n21787 & new_n21790 ;
  assign new_n21792 = new_n21784 & new_n21791 ;
  assign new_n21793 = new_n21777 & new_n21792 ;
  assign new_n21794 = lo1076 & new_n2252 ;
  assign new_n21795 = ~new_n2456 & new_n12442 ;
  assign new_n21796 = ~new_n12420 & ~new_n21795 ;
  assign new_n21797 = new_n12477 & new_n12594 ;
  assign new_n21798 = new_n12486 & new_n20845 ;
  assign new_n21799 = ~new_n12479 & ~new_n21798 ;
  assign new_n21800 = ~new_n21797 & new_n21799 ;
  assign new_n21801 = new_n12452 & ~new_n21800 ;
  assign new_n21802 = ~new_n12452 & new_n21800 ;
  assign new_n21803 = ~new_n21801 & ~new_n21802 ;
  assign new_n21804 = new_n21796 & ~new_n21803 ;
  assign new_n21805 = ~new_n21796 & new_n21801 ;
  assign new_n21806 = ~new_n12452 & ~new_n13278 ;
  assign new_n21807 = ~new_n21800 & new_n21806 ;
  assign new_n21808 = ~new_n21805 & ~new_n21807 ;
  assign new_n21809 = ~new_n21804 & new_n21808 ;
  assign new_n21810 = new_n2446 & ~new_n21809 ;
  assign new_n21811 = new_n13558 & new_n13781 ;
  assign new_n21812 = new_n12369 & new_n12376 ;
  assign new_n21813 = ~new_n20838 & ~new_n21812 ;
  assign new_n21814 = ~new_n12329 & ~new_n21813 ;
  assign new_n21815 = ~new_n21811 & ~new_n21814 ;
  assign new_n21816 = ~new_n2446 & ~new_n21815 ;
  assign new_n21817 = ~new_n21810 & ~new_n21816 ;
  assign new_n21818 = new_n2455 & ~new_n21817 ;
  assign new_n21819 = new_n20654 & ~new_n21818 ;
  assign new_n21820 = new_n2454 & ~new_n21819 ;
  assign new_n21821 = ~new_n2454 & new_n21819 ;
  assign new_n21822 = ~new_n21820 & ~new_n21821 ;
  assign new_n21823 = ~new_n12508 & ~new_n21822 ;
  assign new_n21824 = new_n12508 & new_n21820 ;
  assign new_n21825 = ~new_n12325 & new_n12471 ;
  assign new_n21826 = ~new_n14759 & ~new_n21825 ;
  assign new_n21827 = new_n12386 & ~new_n21826 ;
  assign new_n21828 = ~new_n12580 & ~new_n21827 ;
  assign new_n21829 = ~new_n2454 & new_n12522 ;
  assign new_n21830 = ~new_n21828 & new_n21829 ;
  assign new_n21831 = ~new_n21819 & new_n21830 ;
  assign new_n21832 = ~new_n21824 & ~new_n21831 ;
  assign new_n21833 = ~new_n21823 & new_n21832 ;
  assign new_n21834 = ~new_n2252 & ~new_n21833 ;
  assign new_n21835 = ~new_n21794 & ~new_n21834 ;
  assign new_n21836 = lo1108 & lo1109 ;
  assign new_n21837 = lo1077 & ~new_n21836 ;
  assign new_n21838 = lo1110 & new_n21836 ;
  assign new_n21839 = ~new_n21837 & ~new_n21838 ;
  assign new_n21840 = lo1078 & ~new_n21479 ;
  assign new_n21841 = ~new_n14260 & new_n21483 ;
  assign new_n21842 = lo0112 & new_n10308 ;
  assign new_n21843 = new_n10308 & ~new_n21842 ;
  assign new_n21844 = ~new_n9389 & ~new_n21843 ;
  assign new_n21845 = ~lo0112 & new_n9389 ;
  assign new_n21846 = ~new_n10308 & new_n21845 ;
  assign new_n21847 = ~new_n21844 & ~new_n21846 ;
  assign new_n21848 = ~lo0113 & ~new_n21847 ;
  assign new_n21849 = new_n21482 & new_n21848 ;
  assign new_n21850 = ~new_n21485 & ~new_n21849 ;
  assign new_n21851 = ~new_n21841 & new_n21850 ;
  assign new_n21852 = new_n21482 & ~new_n21851 ;
  assign new_n21853 = ~new_n21482 & new_n21851 ;
  assign new_n21854 = ~new_n21852 & ~new_n21853 ;
  assign new_n21855 = lo1474 & ~new_n21854 ;
  assign new_n21856 = ~lo1474 & new_n21852 ;
  assign new_n21857 = ~new_n5654 & ~new_n21482 ;
  assign new_n21858 = ~new_n21851 & new_n21857 ;
  assign new_n21859 = ~new_n21856 & ~new_n21858 ;
  assign new_n21860 = ~new_n21855 & new_n21859 ;
  assign new_n21861 = new_n21479 & ~new_n21860 ;
  assign new_n21862 = ~new_n21840 & ~new_n21861 ;
  assign new_n21863 = lo1079 & new_n2252 ;
  assign new_n21864 = lo1115 & ~new_n2252 ;
  assign new_n21865 = ~new_n21863 & ~new_n21864 ;
  assign new_n21866 = lo1080 & new_n2252 ;
  assign new_n21867 = lo1116 & ~new_n2252 ;
  assign new_n21868 = ~new_n21866 & ~new_n21867 ;
  assign new_n21869 = lo1081 & new_n2252 ;
  assign new_n21870 = lo1117 & ~new_n2252 ;
  assign new_n21871 = ~new_n21869 & ~new_n21870 ;
  assign new_n21872 = lo1082 & new_n2252 ;
  assign new_n21873 = lo1118 & ~new_n2252 ;
  assign new_n21874 = ~new_n21872 & ~new_n21873 ;
  assign new_n21875 = lo1083 & new_n2252 ;
  assign new_n21876 = lo1119 & ~new_n2252 ;
  assign new_n21877 = ~new_n21875 & ~new_n21876 ;
  assign new_n21878 = lo1084 & new_n2252 ;
  assign new_n21879 = lo1129 & ~new_n2252 ;
  assign new_n21880 = ~new_n21878 & ~new_n21879 ;
  assign new_n21881 = lo1085 & new_n2252 ;
  assign new_n21882 = lo1130 & ~new_n2252 ;
  assign new_n21883 = ~new_n21881 & ~new_n21882 ;
  assign new_n21884 = lo1086 & new_n2252 ;
  assign new_n21885 = lo1131 & ~new_n2252 ;
  assign new_n21886 = ~new_n21884 & ~new_n21885 ;
  assign new_n21887 = lo1087 & new_n2252 ;
  assign new_n21888 = lo1132 & ~new_n2252 ;
  assign new_n21889 = ~new_n21887 & ~new_n21888 ;
  assign new_n21890 = lo1088 & new_n2252 ;
  assign new_n21891 = lo1133 & ~new_n2252 ;
  assign new_n21892 = ~new_n21890 & ~new_n21891 ;
  assign new_n21893 = lo1089 & new_n2252 ;
  assign new_n21894 = lo1134 & ~new_n2252 ;
  assign new_n21895 = ~new_n21893 & ~new_n21894 ;
  assign new_n21896 = lo1090 & new_n2252 ;
  assign new_n21897 = lo1135 & ~new_n2252 ;
  assign new_n21898 = ~new_n21896 & ~new_n21897 ;
  assign new_n21899 = lo1091 & ~new_n21836 ;
  assign new_n21900 = lo1099 & new_n21836 ;
  assign new_n21901 = ~new_n21899 & ~new_n21900 ;
  assign new_n21902 = lo1093 & ~new_n21479 ;
  assign new_n21903 = ~new_n14234 & new_n21483 ;
  assign new_n21904 = lo0112 & new_n13907 ;
  assign new_n21905 = new_n13907 & ~new_n21904 ;
  assign new_n21906 = ~new_n9266 & ~new_n21905 ;
  assign new_n21907 = ~lo0112 & new_n9266 ;
  assign new_n21908 = ~new_n13907 & new_n21907 ;
  assign new_n21909 = ~new_n21906 & ~new_n21908 ;
  assign new_n21910 = ~lo0113 & ~new_n21909 ;
  assign new_n21911 = new_n21482 & new_n21910 ;
  assign new_n21912 = ~new_n21485 & ~new_n21911 ;
  assign new_n21913 = ~new_n21903 & new_n21912 ;
  assign new_n21914 = new_n21482 & ~new_n21913 ;
  assign new_n21915 = ~new_n21482 & new_n21913 ;
  assign new_n21916 = ~new_n21914 & ~new_n21915 ;
  assign new_n21917 = lo1475 & ~new_n21916 ;
  assign new_n21918 = ~lo1475 & new_n21914 ;
  assign new_n21919 = ~new_n5370 & ~new_n21482 ;
  assign new_n21920 = ~new_n21913 & new_n21919 ;
  assign new_n21921 = ~new_n21918 & ~new_n21920 ;
  assign new_n21922 = ~new_n21917 & new_n21921 ;
  assign new_n21923 = new_n21479 & ~new_n21922 ;
  assign new_n21924 = ~new_n21902 & ~new_n21923 ;
  assign new_n21925 = lo1094 & ~new_n21479 ;
  assign new_n21926 = ~new_n14207 & new_n21483 ;
  assign new_n21927 = lo0112 & new_n19223 ;
  assign new_n21928 = new_n19223 & ~new_n21927 ;
  assign new_n21929 = ~new_n9141 & ~new_n21928 ;
  assign new_n21930 = ~lo0112 & new_n9141 ;
  assign new_n21931 = ~new_n19223 & new_n21930 ;
  assign new_n21932 = ~new_n21929 & ~new_n21931 ;
  assign new_n21933 = ~lo0113 & ~new_n21932 ;
  assign new_n21934 = new_n21482 & new_n21933 ;
  assign new_n21935 = ~new_n21485 & ~new_n21934 ;
  assign new_n21936 = ~new_n21926 & new_n21935 ;
  assign new_n21937 = new_n21482 & ~new_n21936 ;
  assign new_n21938 = ~new_n21482 & new_n21936 ;
  assign new_n21939 = ~new_n21937 & ~new_n21938 ;
  assign new_n21940 = lo1476 & ~new_n21939 ;
  assign new_n21941 = ~lo1476 & new_n21937 ;
  assign new_n21942 = ~new_n5086 & ~new_n21482 ;
  assign new_n21943 = ~new_n21936 & new_n21942 ;
  assign new_n21944 = ~new_n21941 & ~new_n21943 ;
  assign new_n21945 = ~new_n21940 & new_n21944 ;
  assign new_n21946 = new_n21479 & ~new_n21945 ;
  assign new_n21947 = ~new_n21925 & ~new_n21946 ;
  assign new_n21948 = lo1095 & ~new_n21836 ;
  assign new_n21949 = lo1097 & new_n21836 ;
  assign new_n21950 = ~new_n21948 & ~new_n21949 ;
  assign new_n21951 = lo1096 & ~new_n21836 ;
  assign new_n21952 = lo1091 & new_n21836 ;
  assign new_n21953 = ~new_n21951 & ~new_n21952 ;
  assign new_n21954 = lo1097 & ~new_n21836 ;
  assign new_n21955 = lo1077 & new_n21836 ;
  assign new_n21956 = ~new_n21954 & ~new_n21955 ;
  assign new_n21957 = lo1098 & ~new_n21836 ;
  assign new_n21958 = lo1096 & new_n21836 ;
  assign new_n21959 = ~new_n21957 & ~new_n21958 ;
  assign new_n21960 = lo1099 & ~new_n21836 ;
  assign new_n21961 = lo1095 & new_n21836 ;
  assign new_n21962 = ~new_n21960 & ~new_n21961 ;
  assign new_n21963 = lo1100 & ~new_n21836 ;
  assign new_n21964 = lo1098 & new_n21836 ;
  assign new_n21965 = ~new_n21963 & ~new_n21964 ;
  assign new_n21966 = lo1101 & new_n2252 ;
  assign new_n21967 = new_n12383 & new_n12592 ;
  assign new_n21968 = new_n13046 & new_n21967 ;
  assign new_n21969 = new_n2264 & new_n12553 ;
  assign new_n21970 = new_n21195 & new_n21969 ;
  assign new_n21971 = ~new_n21968 & ~new_n21970 ;
  assign new_n21972 = ~new_n2252 & new_n12442 ;
  assign new_n21973 = ~new_n21971 & new_n21972 ;
  assign new_n21974 = new_n20585 & new_n21973 ;
  assign new_n21975 = ~new_n21966 & ~new_n21974 ;
  assign new_n21976 = lo1102 & ~new_n20863 ;
  assign new_n21977 = lo1136 & ~new_n14656 ;
  assign new_n21978 = ~lo0977 & lo1139 ;
  assign new_n21979 = ~lo0980 & new_n21978 ;
  assign new_n21980 = ~lo0977 & lo1138 ;
  assign new_n21981 = lo0980 & new_n21980 ;
  assign new_n21982 = ~new_n20868 & ~new_n21981 ;
  assign new_n21983 = ~new_n21979 & new_n21982 ;
  assign new_n21984 = ~lo0977 & ~new_n21983 ;
  assign new_n21985 = lo0977 & new_n21983 ;
  assign new_n21986 = ~new_n21984 & ~new_n21985 ;
  assign new_n21987 = lo1137 & ~new_n21986 ;
  assign new_n21988 = ~lo1137 & new_n21984 ;
  assign new_n21989 = lo0977 & lo1140 ;
  assign new_n21990 = ~new_n21983 & new_n21989 ;
  assign new_n21991 = ~new_n21988 & ~new_n21990 ;
  assign new_n21992 = ~new_n21987 & new_n21991 ;
  assign new_n21993 = new_n14656 & ~new_n21992 ;
  assign new_n21994 = ~new_n21977 & ~new_n21993 ;
  assign new_n21995 = new_n20863 & ~new_n21994 ;
  assign new_n21996 = ~new_n21976 & ~new_n21995 ;
  assign new_n21997 = lo1103 & ~new_n21751 ;
  assign new_n21998 = lo1141 & new_n21751 ;
  assign new_n21999 = ~new_n21997 & ~new_n21998 ;
  assign new_n22000 = lo1104 & ~new_n21746 ;
  assign new_n22001 = lo1141 & new_n21746 ;
  assign new_n22002 = ~new_n22000 & ~new_n22001 ;
  assign new_n22003 = lo1105 & ~new_n21755 ;
  assign new_n22004 = lo1141 & new_n21755 ;
  assign new_n22005 = ~new_n22003 & ~new_n22004 ;
  assign new_n22006 = lo1106 & ~new_n21759 ;
  assign new_n22007 = lo1141 & new_n21759 ;
  assign new_n22008 = ~new_n22006 & ~new_n22007 ;
  assign new_n22009 = lo1107 & ~new_n21248 ;
  assign new_n22010 = lo1272 & new_n21248 ;
  assign new_n22011 = ~new_n22009 & ~new_n22010 ;
  assign new_n22012 = ~lo1448 & lo1449 ;
  assign new_n22013 = new_n20888 & new_n22012 ;
  assign new_n22014 = lo1143 & ~lo1144 ;
  assign new_n22015 = lo1112 & ~new_n20794 ;
  assign new_n22016 = lo0950 & ~new_n14060 ;
  assign new_n22017 = ~lo0950 & ~new_n3281 ;
  assign new_n22018 = ~new_n22016 & ~new_n22017 ;
  assign new_n22019 = lo0949 & new_n22018 ;
  assign new_n22020 = new_n22018 & ~new_n22019 ;
  assign new_n22021 = new_n2718 & ~new_n22020 ;
  assign new_n22022 = ~lo0949 & ~new_n2718 ;
  assign new_n22023 = ~new_n22018 & new_n22022 ;
  assign new_n22024 = ~new_n22021 & ~new_n22023 ;
  assign new_n22025 = new_n20794 & ~new_n22024 ;
  assign new_n22026 = ~new_n22015 & ~new_n22025 ;
  assign new_n22027 = lo0943 & new_n20799 ;
  assign new_n22028 = new_n21039 & new_n22027 ;
  assign new_n22029 = new_n20794 & new_n22028 ;
  assign new_n22030 = lo1113 & ~new_n22029 ;
  assign new_n22031 = lo1114 & new_n22029 ;
  assign new_n22032 = ~new_n22030 & ~new_n22031 ;
  assign new_n22033 = lo1145 & ~new_n2252 ;
  assign new_n22034 = lo1114 & ~new_n22033 ;
  assign new_n22035 = lo0961 & ~new_n14060 ;
  assign new_n22036 = ~lo0961 & ~new_n2739 ;
  assign new_n22037 = ~new_n22035 & ~new_n22036 ;
  assign new_n22038 = lo0960 & new_n22037 ;
  assign new_n22039 = new_n22037 & ~new_n22038 ;
  assign new_n22040 = new_n2718 & ~new_n22039 ;
  assign new_n22041 = ~lo0960 & ~new_n2718 ;
  assign new_n22042 = ~new_n22037 & new_n22041 ;
  assign new_n22043 = ~new_n22040 & ~new_n22042 ;
  assign new_n22044 = new_n22033 & ~new_n22043 ;
  assign new_n22045 = ~new_n22034 & ~new_n22044 ;
  assign new_n22046 = lo1115 & new_n2252 ;
  assign new_n22047 = ~new_n2252 & new_n21721 ;
  assign new_n22048 = new_n15451 & new_n22047 ;
  assign new_n22049 = ~new_n22046 & ~new_n22048 ;
  assign new_n22050 = lo1116 & new_n2252 ;
  assign new_n22051 = new_n20585 & ~new_n21719 ;
  assign new_n22052 = new_n12383 & new_n22051 ;
  assign new_n22053 = new_n16510 & new_n22052 ;
  assign new_n22054 = ~new_n22050 & ~new_n22053 ;
  assign new_n22055 = lo1117 & new_n2252 ;
  assign new_n22056 = new_n16893 & new_n22052 ;
  assign new_n22057 = ~new_n22055 & ~new_n22056 ;
  assign new_n22058 = lo1118 & new_n2252 ;
  assign new_n22059 = new_n18968 & new_n22052 ;
  assign new_n22060 = ~new_n22058 & ~new_n22059 ;
  assign new_n22061 = lo1119 & new_n2252 ;
  assign new_n22062 = new_n19328 & new_n22052 ;
  assign new_n22063 = ~new_n22061 & ~new_n22062 ;
  assign new_n22064 = lo1120 & ~new_n22029 ;
  assign new_n22065 = lo1121 & new_n22029 ;
  assign new_n22066 = ~new_n22064 & ~new_n22065 ;
  assign new_n22067 = lo1121 & ~new_n22033 ;
  assign new_n22068 = lo0960 & new_n5549 ;
  assign new_n22069 = lo0961 & ~new_n14036 ;
  assign new_n22070 = ~lo0961 & ~new_n5560 ;
  assign new_n22071 = ~new_n22069 & ~new_n22070 ;
  assign new_n22072 = ~lo0960 & ~new_n22071 ;
  assign new_n22073 = ~new_n22068 & ~new_n22072 ;
  assign new_n22074 = new_n22033 & ~new_n22073 ;
  assign new_n22075 = ~new_n22067 & ~new_n22074 ;
  assign new_n22076 = lo1122 & ~new_n20794 ;
  assign new_n22077 = lo0949 & new_n5549 ;
  assign new_n22078 = lo0950 & ~new_n14036 ;
  assign new_n22079 = ~lo0950 & ~new_n7374 ;
  assign new_n22080 = ~new_n22078 & ~new_n22079 ;
  assign new_n22081 = ~lo0949 & ~new_n22080 ;
  assign new_n22082 = ~new_n22077 & ~new_n22081 ;
  assign new_n22083 = new_n20794 & ~new_n22082 ;
  assign new_n22084 = ~new_n22076 & ~new_n22083 ;
  assign new_n22085 = lo1123 & ~new_n20794 ;
  assign new_n22086 = lo0949 & new_n2899 ;
  assign new_n22087 = lo0950 & ~new_n14472 ;
  assign new_n22088 = ~lo0950 & ~new_n7512 ;
  assign new_n22089 = ~new_n22087 & ~new_n22088 ;
  assign new_n22090 = ~lo0949 & ~new_n22089 ;
  assign new_n22091 = ~new_n22086 & ~new_n22090 ;
  assign new_n22092 = new_n20794 & ~new_n22091 ;
  assign new_n22093 = ~new_n22085 & ~new_n22092 ;
  assign new_n22094 = lo1124 & ~new_n22029 ;
  assign new_n22095 = lo1125 & new_n22029 ;
  assign new_n22096 = ~new_n22094 & ~new_n22095 ;
  assign new_n22097 = lo1125 & ~new_n22033 ;
  assign new_n22098 = lo0960 & new_n2899 ;
  assign new_n22099 = lo0961 & ~new_n14472 ;
  assign new_n22100 = ~lo0961 & ~new_n2910 ;
  assign new_n22101 = ~new_n22099 & ~new_n22100 ;
  assign new_n22102 = ~lo0960 & ~new_n22101 ;
  assign new_n22103 = ~new_n22098 & ~new_n22102 ;
  assign new_n22104 = new_n22033 & ~new_n22103 ;
  assign new_n22105 = ~new_n22097 & ~new_n22104 ;
  assign new_n22106 = lo1126 & ~new_n20794 ;
  assign new_n22107 = lo0949 & new_n2586 ;
  assign new_n22108 = lo0950 & ~new_n10308 ;
  assign new_n22109 = ~lo0950 & ~new_n9389 ;
  assign new_n22110 = ~new_n22108 & ~new_n22109 ;
  assign new_n22111 = ~lo0949 & ~new_n22110 ;
  assign new_n22112 = ~new_n22107 & ~new_n22111 ;
  assign new_n22113 = new_n20794 & ~new_n22112 ;
  assign new_n22114 = ~new_n22106 & ~new_n22113 ;
  assign new_n22115 = lo1127 & ~new_n22029 ;
  assign new_n22116 = lo1128 & new_n22029 ;
  assign new_n22117 = ~new_n22115 & ~new_n22116 ;
  assign new_n22118 = lo1128 & ~new_n22033 ;
  assign new_n22119 = lo0961 & ~new_n10308 ;
  assign new_n22120 = ~lo0961 & ~new_n2619 ;
  assign new_n22121 = ~new_n22119 & ~new_n22120 ;
  assign new_n22122 = lo0960 & new_n22121 ;
  assign new_n22123 = new_n22121 & ~new_n22122 ;
  assign new_n22124 = new_n2586 & ~new_n22123 ;
  assign new_n22125 = ~lo0960 & ~new_n2586 ;
  assign new_n22126 = ~new_n22121 & new_n22125 ;
  assign new_n22127 = ~new_n22124 & ~new_n22126 ;
  assign new_n22128 = new_n22033 & ~new_n22127 ;
  assign new_n22129 = ~new_n22118 & ~new_n22128 ;
  assign new_n22130 = lo1129 & new_n2252 ;
  assign new_n22131 = ~new_n12441 & ~new_n15547 ;
  assign new_n22132 = ~new_n12887 & new_n22131 ;
  assign new_n22133 = new_n12523 & new_n20535 ;
  assign new_n22134 = ~new_n12496 & ~new_n22133 ;
  assign new_n22135 = new_n22132 & ~new_n22134 ;
  assign new_n22136 = ~new_n12384 & ~new_n22135 ;
  assign new_n22137 = new_n20790 & ~new_n22136 ;
  assign new_n22138 = new_n15451 & new_n22137 ;
  assign new_n22139 = ~new_n22130 & ~new_n22138 ;
  assign new_n22140 = lo1130 & new_n2252 ;
  assign new_n22141 = new_n14732 & new_n20764 ;
  assign new_n22142 = ~new_n22140 & ~new_n22141 ;
  assign new_n22143 = lo1131 & new_n2252 ;
  assign new_n22144 = new_n12761 & new_n20763 ;
  assign new_n22145 = new_n14732 & new_n22144 ;
  assign new_n22146 = ~new_n22143 & ~new_n22145 ;
  assign new_n22147 = lo1132 & new_n2252 ;
  assign new_n22148 = new_n17927 & new_n22144 ;
  assign new_n22149 = ~new_n22147 & ~new_n22148 ;
  assign new_n22150 = lo1133 & new_n2252 ;
  assign new_n22151 = ~new_n2252 & ~new_n12329 ;
  assign new_n22152 = new_n22052 & new_n22151 ;
  assign new_n22153 = ~new_n22150 & ~new_n22152 ;
  assign new_n22154 = lo1134 & new_n2252 ;
  assign new_n22155 = new_n2264 & ~new_n12420 ;
  assign new_n22156 = new_n12420 & new_n12468 ;
  assign new_n22157 = ~new_n22155 & ~new_n22156 ;
  assign new_n22158 = ~new_n12329 & new_n22132 ;
  assign new_n22159 = ~new_n22157 & new_n22158 ;
  assign new_n22160 = ~new_n12547 & ~new_n22159 ;
  assign new_n22161 = ~new_n2252 & ~new_n20788 ;
  assign new_n22162 = ~new_n22160 & new_n22161 ;
  assign new_n22163 = new_n20585 & new_n22162 ;
  assign new_n22164 = ~new_n22154 & ~new_n22163 ;
  assign new_n22165 = lo1135 & new_n2252 ;
  assign new_n22166 = new_n14806 & new_n20764 ;
  assign new_n22167 = ~new_n22165 & ~new_n22166 ;
  assign new_n22168 = lo1136 & ~new_n20863 ;
  assign new_n22169 = lo1230 & ~new_n14656 ;
  assign new_n22170 = ~lo0980 & lo1233 ;
  assign new_n22171 = ~lo0977 & new_n22170 ;
  assign new_n22172 = ~lo0980 & lo1232 ;
  assign new_n22173 = lo0977 & new_n22172 ;
  assign new_n22174 = ~new_n20868 & ~new_n22173 ;
  assign new_n22175 = ~new_n22171 & new_n22174 ;
  assign new_n22176 = ~lo0980 & ~new_n22175 ;
  assign new_n22177 = lo0980 & new_n22175 ;
  assign new_n22178 = ~new_n22176 & ~new_n22177 ;
  assign new_n22179 = lo1231 & ~new_n22178 ;
  assign new_n22180 = ~lo1231 & new_n22176 ;
  assign new_n22181 = lo0980 & lo1234 ;
  assign new_n22182 = ~new_n22175 & new_n22181 ;
  assign new_n22183 = ~new_n22180 & ~new_n22182 ;
  assign new_n22184 = ~new_n22179 & new_n22183 ;
  assign new_n22185 = new_n14656 & ~new_n22184 ;
  assign new_n22186 = ~new_n22169 & ~new_n22185 ;
  assign new_n22187 = new_n20863 & ~new_n22186 ;
  assign new_n22188 = ~new_n22168 & ~new_n22187 ;
  assign new_n22189 = lo1137 & ~new_n21746 ;
  assign new_n22190 = lo1235 & new_n21746 ;
  assign new_n22191 = ~new_n22189 & ~new_n22190 ;
  assign new_n22192 = lo1138 & ~new_n21751 ;
  assign new_n22193 = lo1235 & new_n21751 ;
  assign new_n22194 = ~new_n22192 & ~new_n22193 ;
  assign new_n22195 = lo1139 & ~new_n21755 ;
  assign new_n22196 = lo1235 & new_n21755 ;
  assign new_n22197 = ~new_n22195 & ~new_n22196 ;
  assign new_n22198 = lo1140 & ~new_n21759 ;
  assign new_n22199 = lo1235 & new_n21759 ;
  assign new_n22200 = ~new_n22198 & ~new_n22199 ;
  assign new_n22201 = lo1141 & ~new_n21248 ;
  assign new_n22202 = lo1273 & new_n21248 ;
  assign new_n22203 = ~new_n22201 & ~new_n22202 ;
  assign new_n22204 = lo1016 & ~lo1465 ;
  assign new_n22205 = ~lo1016 & lo1465 ;
  assign new_n22206 = ~new_n22204 & ~new_n22205 ;
  assign new_n22207 = lo0982 & ~lo1460 ;
  assign new_n22208 = ~lo0987 & lo1464 ;
  assign new_n22209 = ~new_n22207 & ~new_n22208 ;
  assign new_n22210 = new_n22206 & new_n22209 ;
  assign new_n22211 = lo0991 & ~lo1467 ;
  assign new_n22212 = ~lo0991 & lo1467 ;
  assign new_n22213 = ~new_n22211 & ~new_n22212 ;
  assign new_n22214 = lo0974 & ~lo1466 ;
  assign new_n22215 = ~lo0974 & lo1466 ;
  assign new_n22216 = ~new_n22214 & ~new_n22215 ;
  assign new_n22217 = new_n22213 & new_n22216 ;
  assign new_n22218 = new_n22210 & new_n22217 ;
  assign new_n22219 = lo0920 & ~lo1461 ;
  assign new_n22220 = ~lo0920 & lo1461 ;
  assign new_n22221 = ~new_n22219 & ~new_n22220 ;
  assign new_n22222 = ~lo0982 & lo1460 ;
  assign new_n22223 = lo0987 & ~lo1464 ;
  assign new_n22224 = ~new_n22222 & ~new_n22223 ;
  assign new_n22225 = new_n22221 & new_n22224 ;
  assign new_n22226 = lo1012 & ~lo1463 ;
  assign new_n22227 = ~lo1012 & lo1463 ;
  assign new_n22228 = ~new_n22226 & ~new_n22227 ;
  assign new_n22229 = lo0928 & ~lo1462 ;
  assign new_n22230 = ~lo0928 & lo1462 ;
  assign new_n22231 = ~new_n22229 & ~new_n22230 ;
  assign new_n22232 = new_n22228 & new_n22231 ;
  assign new_n22233 = new_n22225 & new_n22232 ;
  assign new_n22234 = new_n22218 & new_n22233 ;
  assign new_n22235 = lo1145 & new_n2252 ;
  assign new_n22236 = ~lo1237 & ~new_n21055 ;
  assign new_n22237 = ~new_n2252 & ~new_n22236 ;
  assign new_n22238 = ~new_n22235 & ~new_n22237 ;
  assign new_n22239 = lo1146 & ~new_n22029 ;
  assign new_n22240 = lo1147 & new_n22029 ;
  assign new_n22241 = ~new_n22239 & ~new_n22240 ;
  assign new_n22242 = lo1147 & ~new_n22033 ;
  assign new_n22243 = lo0960 & new_n7122 ;
  assign new_n22244 = lo0961 & ~new_n13907 ;
  assign new_n22245 = ~lo0961 & ~new_n7138 ;
  assign new_n22246 = ~new_n22244 & ~new_n22245 ;
  assign new_n22247 = ~lo0960 & ~new_n22246 ;
  assign new_n22248 = ~new_n22243 & ~new_n22247 ;
  assign new_n22249 = new_n22033 & ~new_n22248 ;
  assign new_n22250 = ~new_n22242 & ~new_n22249 ;
  assign new_n22251 = lo1148 & ~new_n22029 ;
  assign new_n22252 = lo1149 & new_n22029 ;
  assign new_n22253 = ~new_n22251 & ~new_n22252 ;
  assign new_n22254 = lo1149 & ~new_n22033 ;
  assign new_n22255 = lo0960 & new_n6899 ;
  assign new_n22256 = lo0961 & ~new_n19223 ;
  assign new_n22257 = ~lo0961 & ~new_n6917 ;
  assign new_n22258 = ~new_n22256 & ~new_n22257 ;
  assign new_n22259 = ~lo0960 & ~new_n22258 ;
  assign new_n22260 = ~new_n22255 & ~new_n22259 ;
  assign new_n22261 = new_n22033 & ~new_n22260 ;
  assign new_n22262 = ~new_n22254 & ~new_n22261 ;
  assign new_n22263 = lo1150 & ~new_n22029 ;
  assign new_n22264 = lo1151 & new_n22029 ;
  assign new_n22265 = ~new_n22263 & ~new_n22264 ;
  assign new_n22266 = lo1151 & ~new_n22033 ;
  assign new_n22267 = lo0960 & new_n6667 ;
  assign new_n22268 = lo0961 & ~new_n18863 ;
  assign new_n22269 = ~lo0961 & ~new_n6690 ;
  assign new_n22270 = ~new_n22268 & ~new_n22269 ;
  assign new_n22271 = ~lo0960 & ~new_n22270 ;
  assign new_n22272 = ~new_n22267 & ~new_n22271 ;
  assign new_n22273 = new_n22033 & ~new_n22272 ;
  assign new_n22274 = ~new_n22266 & ~new_n22273 ;
  assign new_n22275 = lo1152 & ~new_n22029 ;
  assign new_n22276 = lo1153 & new_n22029 ;
  assign new_n22277 = ~new_n22275 & ~new_n22276 ;
  assign new_n22278 = lo1153 & ~new_n22033 ;
  assign new_n22279 = lo0960 & new_n6433 ;
  assign new_n22280 = lo0961 & ~new_n16735 ;
  assign new_n22281 = ~lo0961 & ~new_n6461 ;
  assign new_n22282 = ~new_n22280 & ~new_n22281 ;
  assign new_n22283 = ~lo0960 & ~new_n22282 ;
  assign new_n22284 = ~new_n22279 & ~new_n22283 ;
  assign new_n22285 = new_n22033 & ~new_n22284 ;
  assign new_n22286 = ~new_n22278 & ~new_n22285 ;
  assign new_n22287 = lo1154 & ~new_n22029 ;
  assign new_n22288 = lo1155 & new_n22029 ;
  assign new_n22289 = ~new_n22287 & ~new_n22288 ;
  assign new_n22290 = lo1155 & ~new_n22033 ;
  assign new_n22291 = lo0960 & new_n6202 ;
  assign new_n22292 = lo0961 & ~new_n16716 ;
  assign new_n22293 = ~lo0961 & ~new_n6225 ;
  assign new_n22294 = ~new_n22292 & ~new_n22293 ;
  assign new_n22295 = ~lo0960 & ~new_n22294 ;
  assign new_n22296 = ~new_n22291 & ~new_n22295 ;
  assign new_n22297 = new_n22033 & ~new_n22296 ;
  assign new_n22298 = ~new_n22290 & ~new_n22297 ;
  assign new_n22299 = lo1156 & ~new_n22029 ;
  assign new_n22300 = lo1157 & new_n22029 ;
  assign new_n22301 = ~new_n22299 & ~new_n22300 ;
  assign new_n22302 = lo1157 & ~new_n22033 ;
  assign new_n22303 = lo0960 & new_n5977 ;
  assign new_n22304 = lo0961 & ~new_n16697 ;
  assign new_n22305 = ~lo0961 & ~new_n5996 ;
  assign new_n22306 = ~new_n22304 & ~new_n22305 ;
  assign new_n22307 = ~lo0960 & ~new_n22306 ;
  assign new_n22308 = ~new_n22303 & ~new_n22307 ;
  assign new_n22309 = new_n22033 & ~new_n22308 ;
  assign new_n22310 = ~new_n22302 & ~new_n22309 ;
  assign new_n22311 = lo1158 & ~new_n22029 ;
  assign new_n22312 = lo1159 & new_n22029 ;
  assign new_n22313 = ~new_n22311 & ~new_n22312 ;
  assign new_n22314 = lo1159 & ~new_n22033 ;
  assign new_n22315 = lo0960 & ~new_n5743 ;
  assign new_n22316 = lo0961 & ~new_n16677 ;
  assign new_n22317 = ~lo0961 & ~new_n5766 ;
  assign new_n22318 = ~new_n22316 & ~new_n22317 ;
  assign new_n22319 = ~lo0960 & ~new_n22318 ;
  assign new_n22320 = ~new_n22315 & ~new_n22319 ;
  assign new_n22321 = new_n22033 & ~new_n22320 ;
  assign new_n22322 = ~new_n22314 & ~new_n22321 ;
  assign new_n22323 = lo1160 & ~new_n22029 ;
  assign new_n22324 = lo1161 & new_n22029 ;
  assign new_n22325 = ~new_n22323 & ~new_n22324 ;
  assign new_n22326 = lo1161 & ~new_n22033 ;
  assign new_n22327 = lo0960 & ~new_n5455 ;
  assign new_n22328 = lo0961 & ~new_n13936 ;
  assign new_n22329 = ~lo0961 & ~new_n5472 ;
  assign new_n22330 = ~new_n22328 & ~new_n22329 ;
  assign new_n22331 = ~lo0960 & ~new_n22330 ;
  assign new_n22332 = ~new_n22327 & ~new_n22331 ;
  assign new_n22333 = new_n22033 & ~new_n22332 ;
  assign new_n22334 = ~new_n22326 & ~new_n22333 ;
  assign new_n22335 = lo1162 & ~new_n22029 ;
  assign new_n22336 = lo1163 & new_n22029 ;
  assign new_n22337 = ~new_n22335 & ~new_n22336 ;
  assign new_n22338 = lo1163 & ~new_n22033 ;
  assign new_n22339 = lo0960 & ~new_n5170 ;
  assign new_n22340 = lo0961 & ~new_n13977 ;
  assign new_n22341 = ~lo0961 & ~new_n5187 ;
  assign new_n22342 = ~new_n22340 & ~new_n22341 ;
  assign new_n22343 = ~lo0960 & ~new_n22342 ;
  assign new_n22344 = ~new_n22339 & ~new_n22343 ;
  assign new_n22345 = new_n22033 & ~new_n22344 ;
  assign new_n22346 = ~new_n22338 & ~new_n22345 ;
  assign new_n22347 = lo1164 & ~new_n22029 ;
  assign new_n22348 = lo1165 & new_n22029 ;
  assign new_n22349 = ~new_n22347 & ~new_n22348 ;
  assign new_n22350 = lo1165 & ~new_n22033 ;
  assign new_n22351 = lo0960 & ~new_n4889 ;
  assign new_n22352 = lo0961 & ~new_n14525 ;
  assign new_n22353 = ~lo0961 & ~new_n4904 ;
  assign new_n22354 = ~new_n22352 & ~new_n22353 ;
  assign new_n22355 = ~lo0960 & ~new_n22354 ;
  assign new_n22356 = ~new_n22351 & ~new_n22355 ;
  assign new_n22357 = new_n22033 & ~new_n22356 ;
  assign new_n22358 = ~new_n22350 & ~new_n22357 ;
  assign new_n22359 = lo1166 & ~new_n22029 ;
  assign new_n22360 = lo1167 & new_n22029 ;
  assign new_n22361 = ~new_n22359 & ~new_n22360 ;
  assign new_n22362 = lo1167 & ~new_n22033 ;
  assign new_n22363 = lo0960 & ~new_n4446 ;
  assign new_n22364 = lo0961 & ~new_n14578 ;
  assign new_n22365 = ~lo0961 & ~new_n4461 ;
  assign new_n22366 = ~new_n22364 & ~new_n22365 ;
  assign new_n22367 = ~lo0960 & ~new_n22366 ;
  assign new_n22368 = ~new_n22363 & ~new_n22367 ;
  assign new_n22369 = new_n22033 & ~new_n22368 ;
  assign new_n22370 = ~new_n22362 & ~new_n22369 ;
  assign new_n22371 = lo1168 & ~new_n22029 ;
  assign new_n22372 = lo1169 & new_n22029 ;
  assign new_n22373 = ~new_n22371 & ~new_n22372 ;
  assign new_n22374 = lo1169 & ~new_n22033 ;
  assign new_n22375 = lo0960 & ~new_n4168 ;
  assign new_n22376 = lo0961 & ~new_n14552 ;
  assign new_n22377 = ~lo0961 & ~new_n4179 ;
  assign new_n22378 = ~new_n22376 & ~new_n22377 ;
  assign new_n22379 = ~lo0960 & ~new_n22378 ;
  assign new_n22380 = ~new_n22375 & ~new_n22379 ;
  assign new_n22381 = new_n22033 & ~new_n22380 ;
  assign new_n22382 = ~new_n22374 & ~new_n22381 ;
  assign new_n22383 = lo1170 & ~new_n22029 ;
  assign new_n22384 = lo1171 & new_n22029 ;
  assign new_n22385 = ~new_n22383 & ~new_n22384 ;
  assign new_n22386 = lo1171 & ~new_n22033 ;
  assign new_n22387 = lo0960 & ~new_n3723 ;
  assign new_n22388 = lo0961 & ~new_n14005 ;
  assign new_n22389 = ~lo0961 & ~new_n3734 ;
  assign new_n22390 = ~new_n22388 & ~new_n22389 ;
  assign new_n22391 = ~lo0960 & ~new_n22390 ;
  assign new_n22392 = ~new_n22387 & ~new_n22391 ;
  assign new_n22393 = new_n22033 & ~new_n22392 ;
  assign new_n22394 = ~new_n22386 & ~new_n22393 ;
  assign new_n22395 = lo1172 & ~new_n22029 ;
  assign new_n22396 = lo1173 & new_n22029 ;
  assign new_n22397 = ~new_n22395 & ~new_n22396 ;
  assign new_n22398 = lo1173 & ~new_n22033 ;
  assign new_n22399 = lo0960 & ~new_n3372 ;
  assign new_n22400 = lo0961 & ~new_n14499 ;
  assign new_n22401 = ~lo0961 & ~new_n3383 ;
  assign new_n22402 = ~new_n22400 & ~new_n22401 ;
  assign new_n22403 = ~lo0960 & ~new_n22402 ;
  assign new_n22404 = ~new_n22399 & ~new_n22403 ;
  assign new_n22405 = new_n22033 & ~new_n22404 ;
  assign new_n22406 = ~new_n22398 & ~new_n22405 ;
  assign new_n22407 = lo1174 & ~new_n22029 ;
  assign new_n22408 = lo1175 & new_n22029 ;
  assign new_n22409 = ~new_n22407 & ~new_n22408 ;
  assign new_n22410 = lo1175 & ~new_n22033 ;
  assign new_n22411 = lo0960 & new_n5265 ;
  assign new_n22412 = lo0961 & ~new_n14446 ;
  assign new_n22413 = ~lo0961 & ~new_n5276 ;
  assign new_n22414 = ~new_n22412 & ~new_n22413 ;
  assign new_n22415 = ~lo0960 & ~new_n22414 ;
  assign new_n22416 = ~new_n22411 & ~new_n22415 ;
  assign new_n22417 = new_n22033 & ~new_n22416 ;
  assign new_n22418 = ~new_n22410 & ~new_n22417 ;
  assign new_n22419 = lo1176 & ~new_n22029 ;
  assign new_n22420 = lo1177 & new_n22029 ;
  assign new_n22421 = ~new_n22419 & ~new_n22420 ;
  assign new_n22422 = lo1177 & ~new_n22033 ;
  assign new_n22423 = lo0960 & new_n4981 ;
  assign new_n22424 = lo0961 & ~new_n14419 ;
  assign new_n22425 = ~lo0961 & ~new_n4992 ;
  assign new_n22426 = ~new_n22424 & ~new_n22425 ;
  assign new_n22427 = ~lo0960 & ~new_n22426 ;
  assign new_n22428 = ~new_n22423 & ~new_n22427 ;
  assign new_n22429 = new_n22033 & ~new_n22428 ;
  assign new_n22430 = ~new_n22422 & ~new_n22429 ;
  assign new_n22431 = lo1178 & ~new_n22029 ;
  assign new_n22432 = lo1179 & new_n22029 ;
  assign new_n22433 = ~new_n22431 & ~new_n22432 ;
  assign new_n22434 = lo1179 & ~new_n22033 ;
  assign new_n22435 = lo0960 & new_n4619 ;
  assign new_n22436 = lo0961 & ~new_n14393 ;
  assign new_n22437 = ~lo0961 & ~new_n4630 ;
  assign new_n22438 = ~new_n22436 & ~new_n22437 ;
  assign new_n22439 = ~lo0960 & ~new_n22438 ;
  assign new_n22440 = ~new_n22435 & ~new_n22439 ;
  assign new_n22441 = new_n22033 & ~new_n22440 ;
  assign new_n22442 = ~new_n22434 & ~new_n22441 ;
  assign new_n22443 = lo1180 & ~new_n22029 ;
  assign new_n22444 = lo1181 & new_n22029 ;
  assign new_n22445 = ~new_n22443 & ~new_n22444 ;
  assign new_n22446 = lo1181 & ~new_n22033 ;
  assign new_n22447 = lo0960 & new_n4257 ;
  assign new_n22448 = lo0961 & ~new_n14366 ;
  assign new_n22449 = ~lo0961 & ~new_n4268 ;
  assign new_n22450 = ~new_n22448 & ~new_n22449 ;
  assign new_n22451 = ~lo0960 & ~new_n22450 ;
  assign new_n22452 = ~new_n22447 & ~new_n22451 ;
  assign new_n22453 = new_n22033 & ~new_n22452 ;
  assign new_n22454 = ~new_n22446 & ~new_n22453 ;
  assign new_n22455 = lo1182 & ~new_n22029 ;
  assign new_n22456 = lo1183 & new_n22029 ;
  assign new_n22457 = ~new_n22455 & ~new_n22456 ;
  assign new_n22458 = lo1183 & ~new_n22033 ;
  assign new_n22459 = lo0960 & new_n3897 ;
  assign new_n22460 = lo0961 & ~new_n14340 ;
  assign new_n22461 = ~lo0961 & ~new_n3908 ;
  assign new_n22462 = ~new_n22460 & ~new_n22461 ;
  assign new_n22463 = ~lo0960 & ~new_n22462 ;
  assign new_n22464 = ~new_n22459 & ~new_n22463 ;
  assign new_n22465 = new_n22033 & ~new_n22464 ;
  assign new_n22466 = ~new_n22458 & ~new_n22465 ;
  assign new_n22467 = lo1184 & ~new_n22029 ;
  assign new_n22468 = lo1185 & new_n22029 ;
  assign new_n22469 = ~new_n22467 & ~new_n22468 ;
  assign new_n22470 = lo1185 & ~new_n22033 ;
  assign new_n22471 = lo0960 & new_n3538 ;
  assign new_n22472 = lo0961 & ~new_n14313 ;
  assign new_n22473 = ~lo0961 & ~new_n3549 ;
  assign new_n22474 = ~new_n22472 & ~new_n22473 ;
  assign new_n22475 = ~lo0960 & ~new_n22474 ;
  assign new_n22476 = ~new_n22471 & ~new_n22475 ;
  assign new_n22477 = new_n22033 & ~new_n22476 ;
  assign new_n22478 = ~new_n22470 & ~new_n22477 ;
  assign new_n22479 = lo1186 & ~new_n22029 ;
  assign new_n22480 = lo1187 & new_n22029 ;
  assign new_n22481 = ~new_n22479 & ~new_n22480 ;
  assign new_n22482 = lo1187 & ~new_n22033 ;
  assign new_n22483 = lo0960 & new_n2813 ;
  assign new_n22484 = lo0961 & ~new_n14287 ;
  assign new_n22485 = ~lo0961 & ~new_n2824 ;
  assign new_n22486 = ~new_n22484 & ~new_n22485 ;
  assign new_n22487 = ~lo0960 & ~new_n22486 ;
  assign new_n22488 = ~new_n22483 & ~new_n22487 ;
  assign new_n22489 = new_n22033 & ~new_n22488 ;
  assign new_n22490 = ~new_n22482 & ~new_n22489 ;
  assign new_n22491 = lo1188 & ~new_n22029 ;
  assign new_n22492 = lo1189 & new_n22029 ;
  assign new_n22493 = ~new_n22491 & ~new_n22492 ;
  assign new_n22494 = lo1189 & ~new_n22033 ;
  assign new_n22495 = lo0960 & new_n4807 ;
  assign new_n22496 = lo0961 & ~new_n14260 ;
  assign new_n22497 = ~lo0961 & ~new_n4818 ;
  assign new_n22498 = ~new_n22496 & ~new_n22497 ;
  assign new_n22499 = ~lo0960 & ~new_n22498 ;
  assign new_n22500 = ~new_n22495 & ~new_n22499 ;
  assign new_n22501 = new_n22033 & ~new_n22500 ;
  assign new_n22502 = ~new_n22494 & ~new_n22501 ;
  assign new_n22503 = lo1190 & ~new_n22029 ;
  assign new_n22504 = lo1191 & new_n22029 ;
  assign new_n22505 = ~new_n22503 & ~new_n22504 ;
  assign new_n22506 = lo1191 & ~new_n22033 ;
  assign new_n22507 = lo0960 & new_n4530 ;
  assign new_n22508 = lo0961 & ~new_n14234 ;
  assign new_n22509 = ~lo0961 & ~new_n4541 ;
  assign new_n22510 = ~new_n22508 & ~new_n22509 ;
  assign new_n22511 = ~lo0960 & ~new_n22510 ;
  assign new_n22512 = ~new_n22507 & ~new_n22511 ;
  assign new_n22513 = new_n22033 & ~new_n22512 ;
  assign new_n22514 = ~new_n22506 & ~new_n22513 ;
  assign new_n22515 = lo1192 & ~new_n22029 ;
  assign new_n22516 = lo1193 & new_n22029 ;
  assign new_n22517 = ~new_n22515 & ~new_n22516 ;
  assign new_n22518 = lo1193 & ~new_n22033 ;
  assign new_n22519 = lo0960 & new_n4086 ;
  assign new_n22520 = lo0961 & ~new_n14207 ;
  assign new_n22521 = ~lo0961 & ~new_n4097 ;
  assign new_n22522 = ~new_n22520 & ~new_n22521 ;
  assign new_n22523 = ~lo0960 & ~new_n22522 ;
  assign new_n22524 = ~new_n22519 & ~new_n22523 ;
  assign new_n22525 = new_n22033 & ~new_n22524 ;
  assign new_n22526 = ~new_n22518 & ~new_n22525 ;
  assign new_n22527 = lo1194 & ~new_n22029 ;
  assign new_n22528 = lo1195 & new_n22029 ;
  assign new_n22529 = ~new_n22527 & ~new_n22528 ;
  assign new_n22530 = lo1195 & ~new_n22033 ;
  assign new_n22531 = lo0960 & new_n3806 ;
  assign new_n22532 = lo0961 & ~new_n14181 ;
  assign new_n22533 = ~lo0961 & ~new_n3817 ;
  assign new_n22534 = ~new_n22532 & ~new_n22533 ;
  assign new_n22535 = ~lo0960 & ~new_n22534 ;
  assign new_n22536 = ~new_n22531 & ~new_n22535 ;
  assign new_n22537 = new_n22033 & ~new_n22536 ;
  assign new_n22538 = ~new_n22530 & ~new_n22537 ;
  assign new_n22539 = lo1196 & ~new_n22029 ;
  assign new_n22540 = lo1197 & new_n22029 ;
  assign new_n22541 = ~new_n22539 & ~new_n22540 ;
  assign new_n22542 = lo1197 & ~new_n22033 ;
  assign new_n22543 = lo0960 & new_n3453 ;
  assign new_n22544 = lo0961 & ~new_n14154 ;
  assign new_n22545 = ~lo0961 & ~new_n3464 ;
  assign new_n22546 = ~new_n22544 & ~new_n22545 ;
  assign new_n22547 = ~lo0960 & ~new_n22546 ;
  assign new_n22548 = ~new_n22543 & ~new_n22547 ;
  assign new_n22549 = new_n22033 & ~new_n22548 ;
  assign new_n22550 = ~new_n22542 & ~new_n22549 ;
  assign new_n22551 = lo1198 & ~new_n22029 ;
  assign new_n22552 = lo1199 & new_n22029 ;
  assign new_n22553 = ~new_n22551 & ~new_n22552 ;
  assign new_n22554 = lo1199 & ~new_n22033 ;
  assign new_n22555 = lo0960 & new_n2990 ;
  assign new_n22556 = lo0961 & ~new_n14128 ;
  assign new_n22557 = ~lo0961 & ~new_n3001 ;
  assign new_n22558 = ~new_n22556 & ~new_n22557 ;
  assign new_n22559 = ~lo0960 & ~new_n22558 ;
  assign new_n22560 = ~new_n22555 & ~new_n22559 ;
  assign new_n22561 = new_n22033 & ~new_n22560 ;
  assign new_n22562 = ~new_n22554 & ~new_n22561 ;
  assign new_n22563 = lo1200 & ~new_n22029 ;
  assign new_n22564 = lo1201 & new_n22029 ;
  assign new_n22565 = ~new_n22563 & ~new_n22564 ;
  assign new_n22566 = lo1201 & ~new_n22033 ;
  assign new_n22567 = lo0960 & new_n3081 ;
  assign new_n22568 = lo0961 & ~new_n14101 ;
  assign new_n22569 = ~lo0961 & ~new_n3092 ;
  assign new_n22570 = ~new_n22568 & ~new_n22569 ;
  assign new_n22571 = ~lo0960 & ~new_n22570 ;
  assign new_n22572 = ~new_n22567 & ~new_n22571 ;
  assign new_n22573 = new_n22033 & ~new_n22572 ;
  assign new_n22574 = ~new_n22566 & ~new_n22573 ;
  assign new_n22575 = lo1202 & ~new_n20794 ;
  assign new_n22576 = lo0949 & new_n7122 ;
  assign new_n22577 = lo0950 & ~new_n13907 ;
  assign new_n22578 = ~lo0950 & ~new_n9266 ;
  assign new_n22579 = ~new_n22577 & ~new_n22578 ;
  assign new_n22580 = ~lo0949 & ~new_n22579 ;
  assign new_n22581 = ~new_n22576 & ~new_n22580 ;
  assign new_n22582 = new_n20794 & ~new_n22581 ;
  assign new_n22583 = ~new_n22575 & ~new_n22582 ;
  assign new_n22584 = lo1203 & ~new_n20794 ;
  assign new_n22585 = lo0949 & new_n5265 ;
  assign new_n22586 = lo0950 & ~new_n14446 ;
  assign new_n22587 = ~lo0950 & ~new_n7249 ;
  assign new_n22588 = ~new_n22586 & ~new_n22587 ;
  assign new_n22589 = ~lo0949 & ~new_n22588 ;
  assign new_n22590 = ~new_n22585 & ~new_n22589 ;
  assign new_n22591 = new_n20794 & ~new_n22590 ;
  assign new_n22592 = ~new_n22584 & ~new_n22591 ;
  assign new_n22593 = lo1204 & ~new_n20794 ;
  assign new_n22594 = lo0949 & new_n6899 ;
  assign new_n22595 = lo0950 & ~new_n19223 ;
  assign new_n22596 = ~lo0950 & ~new_n9141 ;
  assign new_n22597 = ~new_n22595 & ~new_n22596 ;
  assign new_n22598 = ~lo0949 & ~new_n22597 ;
  assign new_n22599 = ~new_n22594 & ~new_n22598 ;
  assign new_n22600 = new_n20794 & ~new_n22599 ;
  assign new_n22601 = ~new_n22593 & ~new_n22600 ;
  assign new_n22602 = lo1205 & ~new_n20794 ;
  assign new_n22603 = lo0949 & new_n4981 ;
  assign new_n22604 = lo0950 & ~new_n14419 ;
  assign new_n22605 = ~lo0950 & ~new_n7026 ;
  assign new_n22606 = ~new_n22604 & ~new_n22605 ;
  assign new_n22607 = ~lo0949 & ~new_n22606 ;
  assign new_n22608 = ~new_n22603 & ~new_n22607 ;
  assign new_n22609 = new_n20794 & ~new_n22608 ;
  assign new_n22610 = ~new_n22602 & ~new_n22609 ;
  assign new_n22611 = lo1206 & ~new_n20794 ;
  assign new_n22612 = lo0949 & new_n6667 ;
  assign new_n22613 = lo0950 & ~new_n18863 ;
  assign new_n22614 = ~lo0950 & ~new_n9021 ;
  assign new_n22615 = ~new_n22613 & ~new_n22614 ;
  assign new_n22616 = ~lo0949 & ~new_n22615 ;
  assign new_n22617 = ~new_n22612 & ~new_n22616 ;
  assign new_n22618 = new_n20794 & ~new_n22617 ;
  assign new_n22619 = ~new_n22611 & ~new_n22618 ;
  assign new_n22620 = lo1207 & ~new_n20794 ;
  assign new_n22621 = lo0949 & new_n4619 ;
  assign new_n22622 = lo0950 & ~new_n14393 ;
  assign new_n22623 = ~lo0950 & ~new_n6801 ;
  assign new_n22624 = ~new_n22622 & ~new_n22623 ;
  assign new_n22625 = ~lo0949 & ~new_n22624 ;
  assign new_n22626 = ~new_n22621 & ~new_n22625 ;
  assign new_n22627 = new_n20794 & ~new_n22626 ;
  assign new_n22628 = ~new_n22620 & ~new_n22627 ;
  assign new_n22629 = lo1208 & ~new_n20794 ;
  assign new_n22630 = lo0949 & new_n6433 ;
  assign new_n22631 = lo0950 & ~new_n16735 ;
  assign new_n22632 = ~lo0950 & ~new_n8902 ;
  assign new_n22633 = ~new_n22631 & ~new_n22632 ;
  assign new_n22634 = ~lo0949 & ~new_n22633 ;
  assign new_n22635 = ~new_n22630 & ~new_n22634 ;
  assign new_n22636 = new_n20794 & ~new_n22635 ;
  assign new_n22637 = ~new_n22629 & ~new_n22636 ;
  assign new_n22638 = lo1209 & ~new_n20794 ;
  assign new_n22639 = lo0949 & new_n4257 ;
  assign new_n22640 = lo0950 & ~new_n14366 ;
  assign new_n22641 = ~lo0950 & ~new_n6571 ;
  assign new_n22642 = ~new_n22640 & ~new_n22641 ;
  assign new_n22643 = ~lo0949 & ~new_n22642 ;
  assign new_n22644 = ~new_n22639 & ~new_n22643 ;
  assign new_n22645 = new_n20794 & ~new_n22644 ;
  assign new_n22646 = ~new_n22638 & ~new_n22645 ;
  assign new_n22647 = lo1210 & ~new_n20794 ;
  assign new_n22648 = lo0949 & new_n6202 ;
  assign new_n22649 = lo0950 & ~new_n16716 ;
  assign new_n22650 = ~lo0950 & ~new_n8780 ;
  assign new_n22651 = ~new_n22649 & ~new_n22650 ;
  assign new_n22652 = ~lo0949 & ~new_n22651 ;
  assign new_n22653 = ~new_n22648 & ~new_n22652 ;
  assign new_n22654 = new_n20794 & ~new_n22653 ;
  assign new_n22655 = ~new_n22647 & ~new_n22654 ;
  assign new_n22656 = lo1211 & ~new_n20794 ;
  assign new_n22657 = lo0949 & new_n3897 ;
  assign new_n22658 = lo0950 & ~new_n14340 ;
  assign new_n22659 = ~lo0950 & ~new_n6336 ;
  assign new_n22660 = ~new_n22658 & ~new_n22659 ;
  assign new_n22661 = ~lo0949 & ~new_n22660 ;
  assign new_n22662 = ~new_n22657 & ~new_n22661 ;
  assign new_n22663 = new_n20794 & ~new_n22662 ;
  assign new_n22664 = ~new_n22656 & ~new_n22663 ;
  assign new_n22665 = lo1212 & ~new_n20794 ;
  assign new_n22666 = lo0949 & new_n5977 ;
  assign new_n22667 = lo0950 & ~new_n16697 ;
  assign new_n22668 = ~lo0950 & ~new_n8659 ;
  assign new_n22669 = ~new_n22667 & ~new_n22668 ;
  assign new_n22670 = ~lo0949 & ~new_n22669 ;
  assign new_n22671 = ~new_n22666 & ~new_n22670 ;
  assign new_n22672 = new_n20794 & ~new_n22671 ;
  assign new_n22673 = ~new_n22665 & ~new_n22672 ;
  assign new_n22674 = lo1213 & ~new_n20794 ;
  assign new_n22675 = lo0949 & new_n3538 ;
  assign new_n22676 = lo0950 & ~new_n14313 ;
  assign new_n22677 = ~lo0950 & ~new_n6106 ;
  assign new_n22678 = ~new_n22676 & ~new_n22677 ;
  assign new_n22679 = ~lo0949 & ~new_n22678 ;
  assign new_n22680 = ~new_n22675 & ~new_n22679 ;
  assign new_n22681 = new_n20794 & ~new_n22680 ;
  assign new_n22682 = ~new_n22674 & ~new_n22681 ;
  assign new_n22683 = lo1214 & ~new_n20794 ;
  assign new_n22684 = lo0949 & ~new_n5743 ;
  assign new_n22685 = lo0950 & ~new_n16677 ;
  assign new_n22686 = ~lo0950 & ~new_n8533 ;
  assign new_n22687 = ~new_n22685 & ~new_n22686 ;
  assign new_n22688 = ~lo0949 & ~new_n22687 ;
  assign new_n22689 = ~new_n22684 & ~new_n22688 ;
  assign new_n22690 = new_n20794 & ~new_n22689 ;
  assign new_n22691 = ~new_n22683 & ~new_n22690 ;
  assign new_n22692 = lo1215 & ~new_n20794 ;
  assign new_n22693 = lo0949 & new_n2813 ;
  assign new_n22694 = lo0950 & ~new_n14287 ;
  assign new_n22695 = ~lo0950 & ~new_n5880 ;
  assign new_n22696 = ~new_n22694 & ~new_n22695 ;
  assign new_n22697 = ~lo0949 & ~new_n22696 ;
  assign new_n22698 = ~new_n22693 & ~new_n22697 ;
  assign new_n22699 = new_n20794 & ~new_n22698 ;
  assign new_n22700 = ~new_n22692 & ~new_n22699 ;
  assign new_n22701 = lo1216 & ~new_n20794 ;
  assign new_n22702 = lo0949 & ~new_n5455 ;
  assign new_n22703 = lo0950 & ~new_n13936 ;
  assign new_n22704 = ~lo0950 & ~new_n8411 ;
  assign new_n22705 = ~new_n22703 & ~new_n22704 ;
  assign new_n22706 = ~lo0949 & ~new_n22705 ;
  assign new_n22707 = ~new_n22702 & ~new_n22706 ;
  assign new_n22708 = new_n20794 & ~new_n22707 ;
  assign new_n22709 = ~new_n22701 & ~new_n22708 ;
  assign new_n22710 = lo1217 & ~new_n20794 ;
  assign new_n22711 = lo0949 & new_n4807 ;
  assign new_n22712 = lo0950 & ~new_n14260 ;
  assign new_n22713 = ~lo0950 & ~new_n5654 ;
  assign new_n22714 = ~new_n22712 & ~new_n22713 ;
  assign new_n22715 = ~lo0949 & ~new_n22714 ;
  assign new_n22716 = ~new_n22711 & ~new_n22715 ;
  assign new_n22717 = new_n20794 & ~new_n22716 ;
  assign new_n22718 = ~new_n22710 & ~new_n22717 ;
  assign new_n22719 = lo1218 & ~new_n20794 ;
  assign new_n22720 = lo0949 & ~new_n5170 ;
  assign new_n22721 = lo0950 & ~new_n13977 ;
  assign new_n22722 = ~lo0950 & ~new_n8281 ;
  assign new_n22723 = ~new_n22721 & ~new_n22722 ;
  assign new_n22724 = ~lo0949 & ~new_n22723 ;
  assign new_n22725 = ~new_n22720 & ~new_n22724 ;
  assign new_n22726 = new_n20794 & ~new_n22725 ;
  assign new_n22727 = ~new_n22719 & ~new_n22726 ;
  assign new_n22728 = lo1219 & ~new_n20794 ;
  assign new_n22729 = lo0949 & new_n4530 ;
  assign new_n22730 = lo0950 & ~new_n14234 ;
  assign new_n22731 = ~lo0950 & ~new_n5370 ;
  assign new_n22732 = ~new_n22730 & ~new_n22731 ;
  assign new_n22733 = ~lo0949 & ~new_n22732 ;
  assign new_n22734 = ~new_n22729 & ~new_n22733 ;
  assign new_n22735 = new_n20794 & ~new_n22734 ;
  assign new_n22736 = ~new_n22728 & ~new_n22735 ;
  assign new_n22737 = lo1220 & ~new_n20794 ;
  assign new_n22738 = lo0949 & ~new_n4889 ;
  assign new_n22739 = lo0950 & ~new_n14525 ;
  assign new_n22740 = ~lo0950 & ~new_n8149 ;
  assign new_n22741 = ~new_n22739 & ~new_n22740 ;
  assign new_n22742 = ~lo0949 & ~new_n22741 ;
  assign new_n22743 = ~new_n22738 & ~new_n22742 ;
  assign new_n22744 = new_n20794 & ~new_n22743 ;
  assign new_n22745 = ~new_n22737 & ~new_n22744 ;
  assign new_n22746 = lo1221 & ~new_n20794 ;
  assign new_n22747 = lo0949 & new_n4086 ;
  assign new_n22748 = lo0950 & ~new_n14207 ;
  assign new_n22749 = ~lo0950 & ~new_n5086 ;
  assign new_n22750 = ~new_n22748 & ~new_n22749 ;
  assign new_n22751 = ~lo0949 & ~new_n22750 ;
  assign new_n22752 = ~new_n22747 & ~new_n22751 ;
  assign new_n22753 = new_n20794 & ~new_n22752 ;
  assign new_n22754 = ~new_n22746 & ~new_n22753 ;
  assign new_n22755 = lo1222 & ~new_n20794 ;
  assign new_n22756 = lo0949 & ~new_n4446 ;
  assign new_n22757 = lo0950 & ~new_n14578 ;
  assign new_n22758 = ~lo0950 & ~new_n8008 ;
  assign new_n22759 = ~new_n22757 & ~new_n22758 ;
  assign new_n22760 = ~lo0949 & ~new_n22759 ;
  assign new_n22761 = ~new_n22756 & ~new_n22760 ;
  assign new_n22762 = new_n20794 & ~new_n22761 ;
  assign new_n22763 = ~new_n22755 & ~new_n22762 ;
  assign new_n22764 = lo1223 & ~new_n20794 ;
  assign new_n22765 = lo0949 & new_n3806 ;
  assign new_n22766 = lo0950 & ~new_n14181 ;
  assign new_n22767 = ~lo0950 & ~new_n4724 ;
  assign new_n22768 = ~new_n22766 & ~new_n22767 ;
  assign new_n22769 = ~lo0949 & ~new_n22768 ;
  assign new_n22770 = ~new_n22765 & ~new_n22769 ;
  assign new_n22771 = new_n20794 & ~new_n22770 ;
  assign new_n22772 = ~new_n22764 & ~new_n22771 ;
  assign new_n22773 = lo1224 & ~new_n20794 ;
  assign new_n22774 = lo0949 & ~new_n4168 ;
  assign new_n22775 = lo0950 & ~new_n14552 ;
  assign new_n22776 = ~lo0950 & ~new_n7883 ;
  assign new_n22777 = ~new_n22775 & ~new_n22776 ;
  assign new_n22778 = ~lo0949 & ~new_n22777 ;
  assign new_n22779 = ~new_n22774 & ~new_n22778 ;
  assign new_n22780 = new_n20794 & ~new_n22779 ;
  assign new_n22781 = ~new_n22773 & ~new_n22780 ;
  assign new_n22782 = lo1225 & ~new_n20794 ;
  assign new_n22783 = lo0949 & new_n3453 ;
  assign new_n22784 = lo0950 & ~new_n14154 ;
  assign new_n22785 = ~lo0950 & ~new_n4362 ;
  assign new_n22786 = ~new_n22784 & ~new_n22785 ;
  assign new_n22787 = ~lo0949 & ~new_n22786 ;
  assign new_n22788 = ~new_n22783 & ~new_n22787 ;
  assign new_n22789 = new_n20794 & ~new_n22788 ;
  assign new_n22790 = ~new_n22782 & ~new_n22789 ;
  assign new_n22791 = lo1226 & ~new_n20794 ;
  assign new_n22792 = lo0949 & ~new_n3723 ;
  assign new_n22793 = lo0950 & ~new_n14005 ;
  assign new_n22794 = ~lo0950 & ~new_n7761 ;
  assign new_n22795 = ~new_n22793 & ~new_n22794 ;
  assign new_n22796 = ~lo0949 & ~new_n22795 ;
  assign new_n22797 = ~new_n22792 & ~new_n22796 ;
  assign new_n22798 = new_n20794 & ~new_n22797 ;
  assign new_n22799 = ~new_n22791 & ~new_n22798 ;
  assign new_n22800 = lo1227 & ~new_n20794 ;
  assign new_n22801 = lo0949 & new_n2990 ;
  assign new_n22802 = lo0950 & ~new_n14128 ;
  assign new_n22803 = ~lo0950 & ~new_n4003 ;
  assign new_n22804 = ~new_n22802 & ~new_n22803 ;
  assign new_n22805 = ~lo0949 & ~new_n22804 ;
  assign new_n22806 = ~new_n22801 & ~new_n22805 ;
  assign new_n22807 = new_n20794 & ~new_n22806 ;
  assign new_n22808 = ~new_n22800 & ~new_n22807 ;
  assign new_n22809 = lo1228 & ~new_n20794 ;
  assign new_n22810 = lo0949 & ~new_n3372 ;
  assign new_n22811 = lo0950 & ~new_n14499 ;
  assign new_n22812 = ~lo0950 & ~new_n7637 ;
  assign new_n22813 = ~new_n22811 & ~new_n22812 ;
  assign new_n22814 = ~lo0949 & ~new_n22813 ;
  assign new_n22815 = ~new_n22810 & ~new_n22814 ;
  assign new_n22816 = new_n20794 & ~new_n22815 ;
  assign new_n22817 = ~new_n22809 & ~new_n22816 ;
  assign new_n22818 = lo1229 & ~new_n20794 ;
  assign new_n22819 = lo0949 & new_n3081 ;
  assign new_n22820 = lo0950 & ~new_n14101 ;
  assign new_n22821 = ~lo0950 & ~new_n3639 ;
  assign new_n22822 = ~new_n22820 & ~new_n22821 ;
  assign new_n22823 = ~lo0949 & ~new_n22822 ;
  assign new_n22824 = ~new_n22819 & ~new_n22823 ;
  assign new_n22825 = new_n20794 & ~new_n22824 ;
  assign new_n22826 = ~new_n22818 & ~new_n22825 ;
  assign new_n22827 = lo1230 & ~new_n20863 ;
  assign new_n22828 = lo1238 & ~new_n14656 ;
  assign new_n22829 = ~lo0977 & lo1241 ;
  assign new_n22830 = ~lo0980 & new_n22829 ;
  assign new_n22831 = ~lo0977 & lo1240 ;
  assign new_n22832 = lo0980 & new_n22831 ;
  assign new_n22833 = ~new_n20868 & ~new_n22832 ;
  assign new_n22834 = ~new_n22830 & new_n22833 ;
  assign new_n22835 = ~lo0977 & ~new_n22834 ;
  assign new_n22836 = lo0977 & new_n22834 ;
  assign new_n22837 = ~new_n22835 & ~new_n22836 ;
  assign new_n22838 = lo1239 & ~new_n22837 ;
  assign new_n22839 = ~lo1239 & new_n22835 ;
  assign new_n22840 = lo0977 & lo1242 ;
  assign new_n22841 = ~new_n22834 & new_n22840 ;
  assign new_n22842 = ~new_n22839 & ~new_n22841 ;
  assign new_n22843 = ~new_n22838 & new_n22842 ;
  assign new_n22844 = new_n14656 & ~new_n22843 ;
  assign new_n22845 = ~new_n22828 & ~new_n22844 ;
  assign new_n22846 = new_n20863 & ~new_n22845 ;
  assign new_n22847 = ~new_n22827 & ~new_n22846 ;
  assign new_n22848 = lo1231 & ~new_n21751 ;
  assign new_n22849 = lo1243 & new_n21751 ;
  assign new_n22850 = ~new_n22848 & ~new_n22849 ;
  assign new_n22851 = lo1232 & ~new_n21746 ;
  assign new_n22852 = lo1243 & new_n21746 ;
  assign new_n22853 = ~new_n22851 & ~new_n22852 ;
  assign new_n22854 = lo1233 & ~new_n21755 ;
  assign new_n22855 = lo1243 & new_n21755 ;
  assign new_n22856 = ~new_n22854 & ~new_n22855 ;
  assign new_n22857 = lo1234 & ~new_n21759 ;
  assign new_n22858 = lo1243 & new_n21759 ;
  assign new_n22859 = ~new_n22857 & ~new_n22858 ;
  assign new_n22860 = lo1235 & ~new_n21248 ;
  assign new_n22861 = lo1274 & new_n21248 ;
  assign new_n22862 = ~new_n22860 & ~new_n22861 ;
  assign new_n22863 = lo1236 & ~lo1245 ;
  assign new_n22864 = lo1244 & ~lo1468 ;
  assign new_n22865 = lo1245 & ~new_n22864 ;
  assign new_n22866 = ~new_n22863 & ~new_n22865 ;
  assign new_n22867 = lo1237 & new_n2252 ;
  assign new_n22868 = lo1246 & ~new_n2252 ;
  assign new_n22869 = ~new_n22867 & ~new_n22868 ;
  assign new_n22870 = lo1238 & ~new_n20863 ;
  assign new_n22871 = lo1247 & ~new_n14656 ;
  assign new_n22872 = ~lo0980 & lo1250 ;
  assign new_n22873 = ~lo0977 & new_n22872 ;
  assign new_n22874 = ~lo0980 & lo1249 ;
  assign new_n22875 = lo0977 & new_n22874 ;
  assign new_n22876 = ~new_n20868 & ~new_n22875 ;
  assign new_n22877 = ~new_n22873 & new_n22876 ;
  assign new_n22878 = ~lo0980 & ~new_n22877 ;
  assign new_n22879 = lo0980 & new_n22877 ;
  assign new_n22880 = ~new_n22878 & ~new_n22879 ;
  assign new_n22881 = lo1248 & ~new_n22880 ;
  assign new_n22882 = ~lo1248 & new_n22878 ;
  assign new_n22883 = lo0980 & lo1251 ;
  assign new_n22884 = ~new_n22877 & new_n22883 ;
  assign new_n22885 = ~new_n22882 & ~new_n22884 ;
  assign new_n22886 = ~new_n22881 & new_n22885 ;
  assign new_n22887 = new_n14656 & ~new_n22886 ;
  assign new_n22888 = ~new_n22871 & ~new_n22887 ;
  assign new_n22889 = new_n20863 & ~new_n22888 ;
  assign new_n22890 = ~new_n22870 & ~new_n22889 ;
  assign new_n22891 = lo1239 & ~new_n21746 ;
  assign new_n22892 = lo1252 & new_n21746 ;
  assign new_n22893 = ~new_n22891 & ~new_n22892 ;
  assign new_n22894 = lo1240 & ~new_n21751 ;
  assign new_n22895 = lo1252 & new_n21751 ;
  assign new_n22896 = ~new_n22894 & ~new_n22895 ;
  assign new_n22897 = lo1241 & ~new_n21755 ;
  assign new_n22898 = lo1252 & new_n21755 ;
  assign new_n22899 = ~new_n22897 & ~new_n22898 ;
  assign new_n22900 = lo1242 & ~new_n21759 ;
  assign new_n22901 = lo1252 & new_n21759 ;
  assign new_n22902 = ~new_n22900 & ~new_n22901 ;
  assign new_n22903 = lo1243 & ~new_n21248 ;
  assign new_n22904 = lo1275 & new_n21248 ;
  assign new_n22905 = ~new_n22903 & ~new_n22904 ;
  assign new_n22906 = lo1244 & ~lo1245 ;
  assign new_n22907 = ~lo1244 & ~lo1254 ;
  assign new_n22908 = lo1468 & ~new_n22907 ;
  assign new_n22909 = ~lo1253 & ~new_n22908 ;
  assign new_n22910 = lo1245 & ~new_n22909 ;
  assign new_n22911 = ~new_n22906 & ~new_n22910 ;
  assign new_n22912 = lo1246 & new_n2252 ;
  assign new_n22913 = new_n15611 & new_n22051 ;
  assign new_n22914 = ~new_n22912 & ~new_n22913 ;
  assign new_n22915 = lo1247 & ~new_n20863 ;
  assign new_n22916 = lo1256 & ~new_n14656 ;
  assign new_n22917 = ~lo0977 & lo1259 ;
  assign new_n22918 = ~lo0980 & new_n22917 ;
  assign new_n22919 = ~lo0977 & lo1258 ;
  assign new_n22920 = lo0980 & new_n22919 ;
  assign new_n22921 = ~new_n20868 & ~new_n22920 ;
  assign new_n22922 = ~new_n22918 & new_n22921 ;
  assign new_n22923 = ~lo0977 & ~new_n22922 ;
  assign new_n22924 = lo0977 & new_n22922 ;
  assign new_n22925 = ~new_n22923 & ~new_n22924 ;
  assign new_n22926 = lo1257 & ~new_n22925 ;
  assign new_n22927 = ~lo1257 & new_n22923 ;
  assign new_n22928 = lo0977 & lo1260 ;
  assign new_n22929 = ~new_n22922 & new_n22928 ;
  assign new_n22930 = ~new_n22927 & ~new_n22929 ;
  assign new_n22931 = ~new_n22926 & new_n22930 ;
  assign new_n22932 = new_n14656 & ~new_n22931 ;
  assign new_n22933 = ~new_n22916 & ~new_n22932 ;
  assign new_n22934 = new_n20863 & ~new_n22933 ;
  assign new_n22935 = ~new_n22915 & ~new_n22934 ;
  assign new_n22936 = lo1248 & ~new_n21751 ;
  assign new_n22937 = lo1261 & new_n21751 ;
  assign new_n22938 = ~new_n22936 & ~new_n22937 ;
  assign new_n22939 = lo1249 & ~new_n21746 ;
  assign new_n22940 = lo1261 & new_n21746 ;
  assign new_n22941 = ~new_n22939 & ~new_n22940 ;
  assign new_n22942 = lo1250 & ~new_n21755 ;
  assign new_n22943 = lo1261 & new_n21755 ;
  assign new_n22944 = ~new_n22942 & ~new_n22943 ;
  assign new_n22945 = lo1251 & ~new_n21759 ;
  assign new_n22946 = lo1261 & new_n21759 ;
  assign new_n22947 = ~new_n22945 & ~new_n22946 ;
  assign new_n22948 = lo1252 & ~new_n21248 ;
  assign new_n22949 = lo1276 & new_n21248 ;
  assign new_n22950 = ~new_n22948 & ~new_n22949 ;
  assign new_n22951 = ~lo1245 & lo1253 ;
  assign new_n22952 = ~lo1236 & lo1468 ;
  assign new_n22953 = lo1254 & ~lo1468 ;
  assign new_n22954 = ~new_n22952 & ~new_n22953 ;
  assign new_n22955 = lo1245 & ~new_n22954 ;
  assign new_n22956 = ~new_n22951 & ~new_n22955 ;
  assign new_n22957 = ~lo1245 & lo1254 ;
  assign new_n22958 = lo1245 & ~lo1468 ;
  assign new_n22959 = ~lo1236 & new_n22958 ;
  assign new_n22960 = ~new_n22957 & ~new_n22959 ;
  assign new_n22961 = lo1074 & ~lo1075 ;
  assign new_n22962 = lo1256 & ~new_n20863 ;
  assign new_n22963 = ~lo0980 & lo1264 ;
  assign new_n22964 = ~lo0977 & new_n22963 ;
  assign new_n22965 = ~lo0980 & lo1263 ;
  assign new_n22966 = lo0977 & new_n22965 ;
  assign new_n22967 = ~new_n20868 & ~new_n22966 ;
  assign new_n22968 = ~new_n22964 & new_n22967 ;
  assign new_n22969 = ~lo0980 & ~new_n22968 ;
  assign new_n22970 = lo0980 & new_n22968 ;
  assign new_n22971 = ~new_n22969 & ~new_n22970 ;
  assign new_n22972 = lo1262 & ~new_n22971 ;
  assign new_n22973 = ~lo1262 & new_n22969 ;
  assign new_n22974 = lo0980 & lo1265 ;
  assign new_n22975 = ~new_n22968 & new_n22974 ;
  assign new_n22976 = new_n14656 & ~new_n22975 ;
  assign new_n22977 = ~new_n22973 & new_n22976 ;
  assign new_n22978 = ~new_n22972 & new_n22977 ;
  assign new_n22979 = new_n20863 & ~new_n22978 ;
  assign new_n22980 = ~new_n22962 & ~new_n22979 ;
  assign new_n22981 = lo1257 & ~new_n21746 ;
  assign new_n22982 = lo1266 & new_n21746 ;
  assign new_n22983 = ~new_n22981 & ~new_n22982 ;
  assign new_n22984 = lo1258 & ~new_n21751 ;
  assign new_n22985 = lo1266 & new_n21751 ;
  assign new_n22986 = ~new_n22984 & ~new_n22985 ;
  assign new_n22987 = lo1259 & ~new_n21755 ;
  assign new_n22988 = lo1266 & new_n21755 ;
  assign new_n22989 = ~new_n22987 & ~new_n22988 ;
  assign new_n22990 = lo1260 & ~new_n21759 ;
  assign new_n22991 = lo1266 & new_n21759 ;
  assign new_n22992 = ~new_n22990 & ~new_n22991 ;
  assign new_n22993 = lo1261 & ~new_n21248 ;
  assign new_n22994 = lo1277 & new_n21248 ;
  assign new_n22995 = ~new_n22993 & ~new_n22994 ;
  assign new_n22996 = lo1262 & ~new_n21751 ;
  assign new_n22997 = lo1267 & new_n21751 ;
  assign new_n22998 = ~new_n22996 & ~new_n22997 ;
  assign new_n22999 = lo1263 & ~new_n21746 ;
  assign new_n23000 = lo1267 & new_n21746 ;
  assign new_n23001 = ~new_n22999 & ~new_n23000 ;
  assign new_n23002 = lo1264 & ~new_n21755 ;
  assign new_n23003 = lo1267 & new_n21755 ;
  assign new_n23004 = ~new_n23002 & ~new_n23003 ;
  assign new_n23005 = lo1265 & ~new_n21759 ;
  assign new_n23006 = lo1267 & new_n21759 ;
  assign new_n23007 = ~new_n23005 & ~new_n23006 ;
  assign new_n23008 = lo1266 & ~new_n21248 ;
  assign new_n23009 = lo1278 & new_n21248 ;
  assign new_n23010 = ~new_n23008 & ~new_n23009 ;
  assign new_n23011 = lo1267 & ~new_n21248 ;
  assign new_n23012 = lo1279 & new_n21248 ;
  assign new_n23013 = ~new_n23011 & ~new_n23012 ;
  assign new_n23014 = ~lo0048 & ~lo0049 ;
  assign new_n23015 = ~lo0047 & ~new_n23014 ;
  assign new_n23016 = lo0050 & ~lo1268 ;
  assign new_n23017 = ~lo1268 & ~new_n23016 ;
  assign new_n23018 = ~new_n23015 & ~new_n23017 ;
  assign new_n23019 = ~lo0050 & lo1268 ;
  assign new_n23020 = new_n23015 & new_n23019 ;
  assign new_n23021 = ~new_n23018 & ~new_n23020 ;
  assign new_n23022 = ~lo0017 & ~new_n23021 ;
  assign new_n23023 = ~lo0017 & ~new_n23022 ;
  assign new_n23024 = lo1269 & ~new_n21479 ;
  assign new_n23025 = lo1474 & ~new_n14601 ;
  assign new_n23026 = new_n14601 & ~new_n21847 ;
  assign new_n23027 = ~new_n23025 & ~new_n23026 ;
  assign new_n23028 = new_n21479 & ~new_n23027 ;
  assign new_n23029 = ~new_n23024 & ~new_n23028 ;
  assign new_n23030 = lo1270 & ~new_n21479 ;
  assign new_n23031 = lo1475 & ~new_n14601 ;
  assign new_n23032 = new_n14601 & ~new_n21909 ;
  assign new_n23033 = ~new_n23031 & ~new_n23032 ;
  assign new_n23034 = new_n21479 & ~new_n23033 ;
  assign new_n23035 = ~new_n23030 & ~new_n23034 ;
  assign new_n23036 = lo1271 & ~new_n21479 ;
  assign new_n23037 = lo1476 & ~new_n14601 ;
  assign new_n23038 = new_n14601 & ~new_n21932 ;
  assign new_n23039 = ~new_n23037 & ~new_n23038 ;
  assign new_n23040 = new_n21479 & ~new_n23039 ;
  assign new_n23041 = ~new_n23036 & ~new_n23040 ;
  assign new_n23042 = lo1272 & ~new_n21479 ;
  assign new_n23043 = lo0113 & lo0114 ;
  assign new_n23044 = ~new_n21847 & ~new_n23043 ;
  assign new_n23045 = lo1474 & new_n23043 ;
  assign new_n23046 = ~new_n23044 & ~new_n23045 ;
  assign new_n23047 = new_n21479 & ~new_n23046 ;
  assign new_n23048 = ~new_n23042 & ~new_n23047 ;
  assign new_n23049 = lo1273 & ~new_n21479 ;
  assign new_n23050 = ~new_n21909 & ~new_n23043 ;
  assign new_n23051 = lo1475 & new_n23043 ;
  assign new_n23052 = ~new_n23050 & ~new_n23051 ;
  assign new_n23053 = new_n21479 & ~new_n23052 ;
  assign new_n23054 = ~new_n23049 & ~new_n23053 ;
  assign new_n23055 = lo1274 & ~new_n21479 ;
  assign new_n23056 = ~new_n21932 & ~new_n23043 ;
  assign new_n23057 = lo1476 & new_n23043 ;
  assign new_n23058 = ~new_n23056 & ~new_n23057 ;
  assign new_n23059 = new_n21479 & ~new_n23058 ;
  assign new_n23060 = ~new_n23055 & ~new_n23059 ;
  assign new_n23061 = lo1275 & ~new_n21479 ;
  assign new_n23062 = ~new_n21514 & ~new_n23043 ;
  assign new_n23063 = lo1470 & new_n23043 ;
  assign new_n23064 = ~new_n23062 & ~new_n23063 ;
  assign new_n23065 = new_n21479 & ~new_n23064 ;
  assign new_n23066 = ~new_n23061 & ~new_n23065 ;
  assign new_n23067 = lo1276 & ~new_n21479 ;
  assign new_n23068 = ~new_n21537 & ~new_n23043 ;
  assign new_n23069 = lo1471 & new_n23043 ;
  assign new_n23070 = ~new_n23068 & ~new_n23069 ;
  assign new_n23071 = new_n21479 & ~new_n23070 ;
  assign new_n23072 = ~new_n23067 & ~new_n23071 ;
  assign new_n23073 = lo1277 & ~new_n21479 ;
  assign new_n23074 = ~new_n21491 & ~new_n23043 ;
  assign new_n23075 = lo1469 & new_n23043 ;
  assign new_n23076 = ~new_n23074 & ~new_n23075 ;
  assign new_n23077 = new_n21479 & ~new_n23076 ;
  assign new_n23078 = ~new_n23073 & ~new_n23077 ;
  assign new_n23079 = lo1278 & ~new_n21479 ;
  assign new_n23080 = ~new_n21560 & ~new_n23043 ;
  assign new_n23081 = lo1472 & new_n23043 ;
  assign new_n23082 = ~new_n23080 & ~new_n23081 ;
  assign new_n23083 = new_n21479 & ~new_n23082 ;
  assign new_n23084 = ~new_n23079 & ~new_n23083 ;
  assign new_n23085 = lo1279 & ~new_n21479 ;
  assign new_n23086 = ~new_n21671 & ~new_n23043 ;
  assign new_n23087 = lo1473 & new_n23043 ;
  assign new_n23088 = ~new_n23086 & ~new_n23087 ;
  assign new_n23089 = new_n21479 & ~new_n23088 ;
  assign new_n23090 = ~new_n23085 & ~new_n23089 ;
  assign new_n23091 = lo1280 & ~new_n21479 ;
  assign new_n23092 = lo0112 & new_n14036 ;
  assign new_n23093 = new_n14036 & ~new_n23092 ;
  assign new_n23094 = ~new_n7374 & ~new_n23093 ;
  assign new_n23095 = ~lo0112 & new_n7374 ;
  assign new_n23096 = ~new_n14036 & new_n23095 ;
  assign new_n23097 = ~new_n23094 & ~new_n23096 ;
  assign new_n23098 = lo0113 & ~new_n23097 ;
  assign new_n23099 = ~new_n21848 & ~new_n23098 ;
  assign new_n23100 = new_n21479 & ~new_n23099 ;
  assign new_n23101 = ~new_n23091 & ~new_n23100 ;
  assign new_n23102 = lo1281 & ~new_n21479 ;
  assign new_n23103 = lo0112 & new_n14446 ;
  assign new_n23104 = new_n14446 & ~new_n23103 ;
  assign new_n23105 = ~new_n7249 & ~new_n23104 ;
  assign new_n23106 = ~lo0112 & new_n7249 ;
  assign new_n23107 = ~new_n14446 & new_n23106 ;
  assign new_n23108 = ~new_n23105 & ~new_n23107 ;
  assign new_n23109 = lo0113 & ~new_n23108 ;
  assign new_n23110 = ~new_n21910 & ~new_n23109 ;
  assign new_n23111 = new_n21479 & ~new_n23110 ;
  assign new_n23112 = ~new_n23102 & ~new_n23111 ;
  assign new_n23113 = lo1282 & ~new_n21479 ;
  assign new_n23114 = lo0112 & new_n14419 ;
  assign new_n23115 = new_n14419 & ~new_n23114 ;
  assign new_n23116 = ~new_n7026 & ~new_n23115 ;
  assign new_n23117 = ~lo0112 & new_n7026 ;
  assign new_n23118 = ~new_n14419 & new_n23117 ;
  assign new_n23119 = ~new_n23116 & ~new_n23118 ;
  assign new_n23120 = lo0113 & ~new_n23119 ;
  assign new_n23121 = ~new_n21933 & ~new_n23120 ;
  assign new_n23122 = new_n21479 & ~new_n23121 ;
  assign new_n23123 = ~new_n23113 & ~new_n23122 ;
  assign new_n23124 = lo1283 & ~new_n21479 ;
  assign new_n23125 = lo0112 & new_n14393 ;
  assign new_n23126 = new_n14393 & ~new_n23125 ;
  assign new_n23127 = ~new_n6801 & ~new_n23126 ;
  assign new_n23128 = ~lo0112 & new_n6801 ;
  assign new_n23129 = ~new_n14393 & new_n23128 ;
  assign new_n23130 = ~new_n23127 & ~new_n23129 ;
  assign new_n23131 = lo0113 & ~new_n23130 ;
  assign new_n23132 = ~new_n21515 & ~new_n23131 ;
  assign new_n23133 = new_n21479 & ~new_n23132 ;
  assign new_n23134 = ~new_n23124 & ~new_n23133 ;
  assign new_n23135 = lo1284 & ~new_n21479 ;
  assign new_n23136 = lo0112 & new_n14366 ;
  assign new_n23137 = new_n14366 & ~new_n23136 ;
  assign new_n23138 = ~new_n6571 & ~new_n23137 ;
  assign new_n23139 = ~lo0112 & new_n6571 ;
  assign new_n23140 = ~new_n14366 & new_n23139 ;
  assign new_n23141 = ~new_n23138 & ~new_n23140 ;
  assign new_n23142 = lo0113 & ~new_n23141 ;
  assign new_n23143 = ~new_n21538 & ~new_n23142 ;
  assign new_n23144 = new_n21479 & ~new_n23143 ;
  assign new_n23145 = ~new_n23135 & ~new_n23144 ;
  assign new_n23146 = lo0051 & new_n14680 ;
  assign new_n23147 = ~lo0051 & ~new_n14680 ;
  assign new_n23148 = ~new_n2241 & ~new_n23147 ;
  assign new_n23149 = ~new_n23146 & new_n23148 ;
  assign new_n23150 = new_n14677 & new_n23149 ;
  assign new_n23151 = lo0899 & lo1285 ;
  assign new_n23152 = ~new_n23150 & new_n23151 ;
  assign new_n23153 = new_n14670 & new_n23152 ;
  assign new_n23154 = ~lo0899 & lo1285 ;
  assign new_n23155 = ~new_n23150 & new_n23154 ;
  assign new_n23156 = ~new_n23150 & ~new_n23155 ;
  assign new_n23157 = ~new_n23153 & new_n23156 ;
  assign new_n23158 = ~lo0017 & ~new_n23157 ;
  assign new_n23159 = ~lo0066 & ~lo0932 ;
  assign new_n23160 = ~lo0931 & new_n23159 ;
  assign new_n23161 = ~new_n2252 & ~new_n23160 ;
  assign new_n23162 = lo1286 & ~new_n23161 ;
  assign new_n23163 = lo0931 & new_n5455 ;
  assign new_n23164 = new_n5455 & ~new_n23163 ;
  assign new_n23165 = ~new_n13936 & ~new_n23164 ;
  assign new_n23166 = ~lo0931 & ~new_n5455 ;
  assign new_n23167 = new_n13936 & new_n23166 ;
  assign new_n23168 = ~new_n23165 & ~new_n23167 ;
  assign new_n23169 = ~lo0932 & ~new_n23168 ;
  assign new_n23170 = lo0111 & lo0932 ;
  assign new_n23171 = ~new_n23169 & ~new_n23170 ;
  assign new_n23172 = new_n23161 & ~new_n23171 ;
  assign new_n23173 = ~new_n23162 & ~new_n23172 ;
  assign new_n23174 = new_n20794 & ~new_n22028 ;
  assign new_n23175 = lo0951 & ~new_n2252 ;
  assign new_n23176 = ~lo0938 & ~new_n23175 ;
  assign new_n23177 = ~new_n23174 & new_n23176 ;
  assign new_n23178 = lo1287 & new_n23177 ;
  assign new_n23179 = pi425 & new_n2138 ;
  assign new_n23180 = pi424 & new_n2138 ;
  assign new_n23181 = pi423 & new_n2138 ;
  assign new_n23182 = pi422 & new_n2138 ;
  assign new_n23183 = pi421 & new_n2138 ;
  assign new_n23184 = pi420 & new_n2138 ;
  assign new_n23185 = pi419 & new_n2138 ;
  assign new_n23186 = pi418 & new_n2138 ;
  assign new_n23187 = pi417 & new_n2138 ;
  assign new_n23188 = lo1361 & new_n23187 ;
  assign new_n23189 = ~lo1382 & new_n23188 ;
  assign new_n23190 = ~lo1382 & ~new_n23189 ;
  assign new_n23191 = new_n23186 & ~new_n23190 ;
  assign new_n23192 = lo1382 & new_n23188 ;
  assign new_n23193 = ~new_n23186 & new_n23192 ;
  assign new_n23194 = ~new_n23191 & ~new_n23193 ;
  assign new_n23195 = ~lo1370 & ~new_n23194 ;
  assign new_n23196 = ~lo1370 & ~new_n23195 ;
  assign new_n23197 = new_n23185 & ~new_n23196 ;
  assign new_n23198 = lo1370 & ~new_n23194 ;
  assign new_n23199 = ~new_n23185 & new_n23198 ;
  assign new_n23200 = ~new_n23197 & ~new_n23199 ;
  assign new_n23201 = ~lo1376 & ~new_n23200 ;
  assign new_n23202 = ~lo1376 & ~new_n23201 ;
  assign new_n23203 = new_n23184 & ~new_n23202 ;
  assign new_n23204 = lo1376 & ~new_n23200 ;
  assign new_n23205 = ~new_n23184 & new_n23204 ;
  assign new_n23206 = ~new_n23203 & ~new_n23205 ;
  assign new_n23207 = ~lo1298 & ~new_n23206 ;
  assign new_n23208 = ~lo1298 & ~new_n23207 ;
  assign new_n23209 = new_n23183 & ~new_n23208 ;
  assign new_n23210 = lo1298 & ~new_n23206 ;
  assign new_n23211 = ~new_n23183 & new_n23210 ;
  assign new_n23212 = ~new_n23209 & ~new_n23211 ;
  assign new_n23213 = ~lo1337 & ~new_n23212 ;
  assign new_n23214 = ~lo1337 & ~new_n23213 ;
  assign new_n23215 = new_n23182 & ~new_n23214 ;
  assign new_n23216 = lo1337 & ~new_n23212 ;
  assign new_n23217 = ~new_n23182 & new_n23216 ;
  assign new_n23218 = ~new_n23215 & ~new_n23217 ;
  assign new_n23219 = ~lo1321 & ~new_n23218 ;
  assign new_n23220 = ~lo1321 & ~new_n23219 ;
  assign new_n23221 = new_n23181 & ~new_n23220 ;
  assign new_n23222 = lo1321 & ~new_n23218 ;
  assign new_n23223 = ~new_n23181 & new_n23222 ;
  assign new_n23224 = ~new_n23221 & ~new_n23223 ;
  assign new_n23225 = ~lo1310 & ~new_n23224 ;
  assign new_n23226 = ~lo1310 & ~new_n23225 ;
  assign new_n23227 = new_n23180 & ~new_n23226 ;
  assign new_n23228 = lo1310 & ~new_n23224 ;
  assign new_n23229 = ~new_n23180 & new_n23228 ;
  assign new_n23230 = ~new_n23227 & ~new_n23229 ;
  assign new_n23231 = lo1287 & ~new_n23230 ;
  assign new_n23232 = ~lo1287 & new_n23230 ;
  assign new_n23233 = ~new_n23231 & ~new_n23232 ;
  assign new_n23234 = new_n23179 & ~new_n23233 ;
  assign new_n23235 = ~lo1287 & ~new_n23230 ;
  assign new_n23236 = lo1287 & new_n23230 ;
  assign new_n23237 = ~new_n23235 & ~new_n23236 ;
  assign new_n23238 = ~new_n23179 & ~new_n23237 ;
  assign new_n23239 = ~new_n23234 & ~new_n23238 ;
  assign new_n23240 = ~new_n2071 & new_n2138 ;
  assign new_n23241 = lo0938 & ~lo0939 ;
  assign new_n23242 = new_n21023 & new_n23241 ;
  assign new_n23243 = pi463 & new_n2138 ;
  assign new_n23244 = lo1112 & ~new_n2138 ;
  assign new_n23245 = lo1113 & ~new_n2022 ;
  assign new_n23246 = lo1114 & new_n2022 ;
  assign new_n23247 = ~new_n23245 & ~new_n23246 ;
  assign new_n23248 = new_n23244 & ~new_n23247 ;
  assign new_n23249 = ~new_n23243 & ~new_n23248 ;
  assign new_n23250 = new_n2071 & ~new_n23249 ;
  assign new_n23251 = ~new_n2134 & new_n23244 ;
  assign new_n23252 = ~new_n2138 & ~new_n23247 ;
  assign new_n23253 = lo1229 & new_n23252 ;
  assign new_n23254 = ~new_n2130 & new_n23244 ;
  assign new_n23255 = lo1227 & new_n23252 ;
  assign new_n23256 = ~new_n2126 & new_n23244 ;
  assign new_n23257 = lo1225 & new_n23252 ;
  assign new_n23258 = ~new_n2122 & new_n23244 ;
  assign new_n23259 = lo1223 & new_n23252 ;
  assign new_n23260 = ~new_n2118 & new_n23244 ;
  assign new_n23261 = lo1221 & new_n23252 ;
  assign new_n23262 = ~new_n2114 & new_n23244 ;
  assign new_n23263 = lo1219 & new_n23252 ;
  assign new_n23264 = ~new_n2110 & new_n23244 ;
  assign new_n23265 = lo1217 & new_n23252 ;
  assign new_n23266 = ~new_n2106 & new_n23244 ;
  assign new_n23267 = lo1215 & new_n23252 ;
  assign new_n23268 = ~new_n2102 & new_n23244 ;
  assign new_n23269 = lo1213 & new_n23252 ;
  assign new_n23270 = ~new_n2098 & new_n23244 ;
  assign new_n23271 = lo1211 & new_n23252 ;
  assign new_n23272 = ~new_n2094 & new_n23244 ;
  assign new_n23273 = lo1209 & new_n23252 ;
  assign new_n23274 = ~new_n2090 & new_n23244 ;
  assign new_n23275 = lo1207 & new_n23252 ;
  assign new_n23276 = ~new_n2086 & new_n23244 ;
  assign new_n23277 = lo1205 & new_n23252 ;
  assign new_n23278 = ~new_n2082 & new_n23244 ;
  assign new_n23279 = lo1203 & new_n23252 ;
  assign new_n23280 = ~new_n2078 & new_n23244 ;
  assign new_n23281 = lo1122 & new_n23252 ;
  assign new_n23282 = ~new_n2074 & new_n23244 ;
  assign new_n23283 = lo1123 & new_n23252 ;
  assign new_n23284 = ~new_n2074 & new_n23240 ;
  assign new_n23285 = ~new_n2185 & new_n23252 ;
  assign new_n23286 = ~new_n23284 & ~new_n23285 ;
  assign new_n23287 = lo1228 & ~new_n23286 ;
  assign new_n23288 = lo1123 & new_n23240 ;
  assign new_n23289 = ~new_n2185 & new_n23244 ;
  assign new_n23290 = ~new_n23288 & ~new_n23289 ;
  assign new_n23291 = ~new_n2067 & ~new_n23290 ;
  assign new_n23292 = lo1226 & ~new_n23286 ;
  assign new_n23293 = ~new_n2064 & ~new_n23290 ;
  assign new_n23294 = lo1224 & ~new_n23286 ;
  assign new_n23295 = ~new_n2061 & ~new_n23290 ;
  assign new_n23296 = lo1222 & ~new_n23286 ;
  assign new_n23297 = ~new_n2058 & ~new_n23290 ;
  assign new_n23298 = lo1220 & ~new_n23286 ;
  assign new_n23299 = ~new_n2055 & ~new_n23290 ;
  assign new_n23300 = lo1218 & ~new_n23286 ;
  assign new_n23301 = ~new_n2052 & ~new_n23290 ;
  assign new_n23302 = lo1216 & ~new_n23286 ;
  assign new_n23303 = ~new_n2049 & ~new_n23290 ;
  assign new_n23304 = lo1214 & ~new_n23286 ;
  assign new_n23305 = ~new_n2046 & ~new_n23290 ;
  assign new_n23306 = lo1212 & ~new_n23286 ;
  assign new_n23307 = ~new_n2043 & ~new_n23290 ;
  assign new_n23308 = lo1210 & ~new_n23286 ;
  assign new_n23309 = ~new_n2040 & ~new_n23290 ;
  assign new_n23310 = lo1208 & ~new_n23286 ;
  assign new_n23311 = ~new_n2037 & ~new_n23290 ;
  assign new_n23312 = lo1206 & ~new_n23286 ;
  assign new_n23313 = ~new_n2034 & ~new_n23290 ;
  assign new_n23314 = lo1204 & ~new_n23286 ;
  assign new_n23315 = ~new_n2031 & ~new_n23290 ;
  assign new_n23316 = lo1202 & ~new_n23286 ;
  assign new_n23317 = ~new_n2028 & ~new_n23290 ;
  assign new_n23318 = lo1126 & ~new_n23286 ;
  assign new_n23319 = ~new_n2025 & ~new_n23290 ;
  assign new_n23320 = new_n23318 & new_n23319 ;
  assign new_n23321 = ~new_n23317 & new_n23320 ;
  assign new_n23322 = ~new_n23317 & ~new_n23321 ;
  assign new_n23323 = new_n23316 & ~new_n23322 ;
  assign new_n23324 = new_n23317 & new_n23320 ;
  assign new_n23325 = ~new_n23316 & new_n23324 ;
  assign new_n23326 = ~new_n23323 & ~new_n23325 ;
  assign new_n23327 = ~new_n23315 & ~new_n23326 ;
  assign new_n23328 = ~new_n23315 & ~new_n23327 ;
  assign new_n23329 = new_n23314 & ~new_n23328 ;
  assign new_n23330 = new_n23315 & ~new_n23326 ;
  assign new_n23331 = ~new_n23314 & new_n23330 ;
  assign new_n23332 = ~new_n23329 & ~new_n23331 ;
  assign new_n23333 = ~new_n23313 & ~new_n23332 ;
  assign new_n23334 = ~new_n23313 & ~new_n23333 ;
  assign new_n23335 = new_n23312 & ~new_n23334 ;
  assign new_n23336 = new_n23313 & ~new_n23332 ;
  assign new_n23337 = ~new_n23312 & new_n23336 ;
  assign new_n23338 = ~new_n23335 & ~new_n23337 ;
  assign new_n23339 = ~new_n23311 & ~new_n23338 ;
  assign new_n23340 = ~new_n23311 & ~new_n23339 ;
  assign new_n23341 = new_n23310 & ~new_n23340 ;
  assign new_n23342 = new_n23311 & ~new_n23338 ;
  assign new_n23343 = ~new_n23310 & new_n23342 ;
  assign new_n23344 = ~new_n23341 & ~new_n23343 ;
  assign new_n23345 = ~new_n23309 & ~new_n23344 ;
  assign new_n23346 = ~new_n23309 & ~new_n23345 ;
  assign new_n23347 = new_n23308 & ~new_n23346 ;
  assign new_n23348 = new_n23309 & ~new_n23344 ;
  assign new_n23349 = ~new_n23308 & new_n23348 ;
  assign new_n23350 = ~new_n23347 & ~new_n23349 ;
  assign new_n23351 = ~new_n23307 & ~new_n23350 ;
  assign new_n23352 = ~new_n23307 & ~new_n23351 ;
  assign new_n23353 = new_n23306 & ~new_n23352 ;
  assign new_n23354 = new_n23307 & ~new_n23350 ;
  assign new_n23355 = ~new_n23306 & new_n23354 ;
  assign new_n23356 = ~new_n23353 & ~new_n23355 ;
  assign new_n23357 = ~new_n23305 & ~new_n23356 ;
  assign new_n23358 = ~new_n23305 & ~new_n23357 ;
  assign new_n23359 = new_n23304 & ~new_n23358 ;
  assign new_n23360 = new_n23305 & ~new_n23356 ;
  assign new_n23361 = ~new_n23304 & new_n23360 ;
  assign new_n23362 = ~new_n23359 & ~new_n23361 ;
  assign new_n23363 = ~new_n23303 & ~new_n23362 ;
  assign new_n23364 = ~new_n23303 & ~new_n23363 ;
  assign new_n23365 = new_n23302 & ~new_n23364 ;
  assign new_n23366 = new_n23303 & ~new_n23362 ;
  assign new_n23367 = ~new_n23302 & new_n23366 ;
  assign new_n23368 = ~new_n23365 & ~new_n23367 ;
  assign new_n23369 = ~new_n23301 & ~new_n23368 ;
  assign new_n23370 = ~new_n23301 & ~new_n23369 ;
  assign new_n23371 = new_n23300 & ~new_n23370 ;
  assign new_n23372 = new_n23301 & ~new_n23368 ;
  assign new_n23373 = ~new_n23300 & new_n23372 ;
  assign new_n23374 = ~new_n23371 & ~new_n23373 ;
  assign new_n23375 = ~new_n23299 & ~new_n23374 ;
  assign new_n23376 = ~new_n23299 & ~new_n23375 ;
  assign new_n23377 = new_n23298 & ~new_n23376 ;
  assign new_n23378 = new_n23299 & ~new_n23374 ;
  assign new_n23379 = ~new_n23298 & new_n23378 ;
  assign new_n23380 = ~new_n23377 & ~new_n23379 ;
  assign new_n23381 = ~new_n23297 & ~new_n23380 ;
  assign new_n23382 = ~new_n23297 & ~new_n23381 ;
  assign new_n23383 = new_n23296 & ~new_n23382 ;
  assign new_n23384 = new_n23297 & ~new_n23380 ;
  assign new_n23385 = ~new_n23296 & new_n23384 ;
  assign new_n23386 = ~new_n23383 & ~new_n23385 ;
  assign new_n23387 = ~new_n23295 & ~new_n23386 ;
  assign new_n23388 = ~new_n23295 & ~new_n23387 ;
  assign new_n23389 = new_n23294 & ~new_n23388 ;
  assign new_n23390 = new_n23295 & ~new_n23386 ;
  assign new_n23391 = ~new_n23294 & new_n23390 ;
  assign new_n23392 = ~new_n23389 & ~new_n23391 ;
  assign new_n23393 = ~new_n23293 & ~new_n23392 ;
  assign new_n23394 = ~new_n23293 & ~new_n23393 ;
  assign new_n23395 = new_n23292 & ~new_n23394 ;
  assign new_n23396 = new_n23293 & ~new_n23392 ;
  assign new_n23397 = ~new_n23292 & new_n23396 ;
  assign new_n23398 = ~new_n23395 & ~new_n23397 ;
  assign new_n23399 = ~new_n23291 & ~new_n23398 ;
  assign new_n23400 = ~new_n23291 & ~new_n23399 ;
  assign new_n23401 = new_n23287 & ~new_n23400 ;
  assign new_n23402 = new_n23291 & ~new_n23398 ;
  assign new_n23403 = ~new_n23287 & new_n23402 ;
  assign new_n23404 = ~new_n23401 & ~new_n23403 ;
  assign new_n23405 = ~new_n23283 & ~new_n23404 ;
  assign new_n23406 = ~new_n23283 & ~new_n23405 ;
  assign new_n23407 = new_n23282 & ~new_n23406 ;
  assign new_n23408 = new_n23283 & ~new_n23404 ;
  assign new_n23409 = ~new_n23282 & new_n23408 ;
  assign new_n23410 = ~new_n23407 & ~new_n23409 ;
  assign new_n23411 = ~new_n23281 & ~new_n23410 ;
  assign new_n23412 = ~new_n23281 & ~new_n23411 ;
  assign new_n23413 = new_n23280 & ~new_n23412 ;
  assign new_n23414 = new_n23281 & ~new_n23410 ;
  assign new_n23415 = ~new_n23280 & new_n23414 ;
  assign new_n23416 = ~new_n23413 & ~new_n23415 ;
  assign new_n23417 = ~new_n23279 & ~new_n23416 ;
  assign new_n23418 = ~new_n23279 & ~new_n23417 ;
  assign new_n23419 = new_n23278 & ~new_n23418 ;
  assign new_n23420 = new_n23279 & ~new_n23416 ;
  assign new_n23421 = ~new_n23278 & new_n23420 ;
  assign new_n23422 = ~new_n23419 & ~new_n23421 ;
  assign new_n23423 = ~new_n23277 & ~new_n23422 ;
  assign new_n23424 = ~new_n23277 & ~new_n23423 ;
  assign new_n23425 = new_n23276 & ~new_n23424 ;
  assign new_n23426 = new_n23277 & ~new_n23422 ;
  assign new_n23427 = ~new_n23276 & new_n23426 ;
  assign new_n23428 = ~new_n23425 & ~new_n23427 ;
  assign new_n23429 = ~new_n23275 & ~new_n23428 ;
  assign new_n23430 = ~new_n23275 & ~new_n23429 ;
  assign new_n23431 = new_n23274 & ~new_n23430 ;
  assign new_n23432 = new_n23275 & ~new_n23428 ;
  assign new_n23433 = ~new_n23274 & new_n23432 ;
  assign new_n23434 = ~new_n23431 & ~new_n23433 ;
  assign new_n23435 = ~new_n23273 & ~new_n23434 ;
  assign new_n23436 = ~new_n23273 & ~new_n23435 ;
  assign new_n23437 = new_n23272 & ~new_n23436 ;
  assign new_n23438 = new_n23273 & ~new_n23434 ;
  assign new_n23439 = ~new_n23272 & new_n23438 ;
  assign new_n23440 = ~new_n23437 & ~new_n23439 ;
  assign new_n23441 = ~new_n23271 & ~new_n23440 ;
  assign new_n23442 = ~new_n23271 & ~new_n23441 ;
  assign new_n23443 = new_n23270 & ~new_n23442 ;
  assign new_n23444 = new_n23271 & ~new_n23440 ;
  assign new_n23445 = ~new_n23270 & new_n23444 ;
  assign new_n23446 = ~new_n23443 & ~new_n23445 ;
  assign new_n23447 = ~new_n23269 & ~new_n23446 ;
  assign new_n23448 = ~new_n23269 & ~new_n23447 ;
  assign new_n23449 = new_n23268 & ~new_n23448 ;
  assign new_n23450 = new_n23269 & ~new_n23446 ;
  assign new_n23451 = ~new_n23268 & new_n23450 ;
  assign new_n23452 = ~new_n23449 & ~new_n23451 ;
  assign new_n23453 = ~new_n23267 & ~new_n23452 ;
  assign new_n23454 = ~new_n23267 & ~new_n23453 ;
  assign new_n23455 = new_n23266 & ~new_n23454 ;
  assign new_n23456 = new_n23267 & ~new_n23452 ;
  assign new_n23457 = ~new_n23266 & new_n23456 ;
  assign new_n23458 = ~new_n23455 & ~new_n23457 ;
  assign new_n23459 = ~new_n23265 & ~new_n23458 ;
  assign new_n23460 = ~new_n23265 & ~new_n23459 ;
  assign new_n23461 = new_n23264 & ~new_n23460 ;
  assign new_n23462 = new_n23265 & ~new_n23458 ;
  assign new_n23463 = ~new_n23264 & new_n23462 ;
  assign new_n23464 = ~new_n23461 & ~new_n23463 ;
  assign new_n23465 = ~new_n23263 & ~new_n23464 ;
  assign new_n23466 = ~new_n23263 & ~new_n23465 ;
  assign new_n23467 = new_n23262 & ~new_n23466 ;
  assign new_n23468 = new_n23263 & ~new_n23464 ;
  assign new_n23469 = ~new_n23262 & new_n23468 ;
  assign new_n23470 = ~new_n23467 & ~new_n23469 ;
  assign new_n23471 = ~new_n23261 & ~new_n23470 ;
  assign new_n23472 = ~new_n23261 & ~new_n23471 ;
  assign new_n23473 = new_n23260 & ~new_n23472 ;
  assign new_n23474 = new_n23261 & ~new_n23470 ;
  assign new_n23475 = ~new_n23260 & new_n23474 ;
  assign new_n23476 = ~new_n23473 & ~new_n23475 ;
  assign new_n23477 = ~new_n23259 & ~new_n23476 ;
  assign new_n23478 = ~new_n23259 & ~new_n23477 ;
  assign new_n23479 = new_n23258 & ~new_n23478 ;
  assign new_n23480 = new_n23259 & ~new_n23476 ;
  assign new_n23481 = ~new_n23258 & new_n23480 ;
  assign new_n23482 = ~new_n23479 & ~new_n23481 ;
  assign new_n23483 = ~new_n23257 & ~new_n23482 ;
  assign new_n23484 = ~new_n23257 & ~new_n23483 ;
  assign new_n23485 = new_n23256 & ~new_n23484 ;
  assign new_n23486 = new_n23257 & ~new_n23482 ;
  assign new_n23487 = ~new_n23256 & new_n23486 ;
  assign new_n23488 = ~new_n23485 & ~new_n23487 ;
  assign new_n23489 = ~new_n23255 & ~new_n23488 ;
  assign new_n23490 = ~new_n23255 & ~new_n23489 ;
  assign new_n23491 = new_n23254 & ~new_n23490 ;
  assign new_n23492 = new_n23255 & ~new_n23488 ;
  assign new_n23493 = ~new_n23254 & new_n23492 ;
  assign new_n23494 = ~new_n23491 & ~new_n23493 ;
  assign new_n23495 = ~new_n23253 & ~new_n23494 ;
  assign new_n23496 = ~new_n23253 & ~new_n23495 ;
  assign new_n23497 = new_n23251 & ~new_n23496 ;
  assign new_n23498 = new_n23253 & ~new_n23494 ;
  assign new_n23499 = ~new_n23251 & new_n23498 ;
  assign new_n23500 = ~new_n23497 & ~new_n23499 ;
  assign new_n23501 = ~new_n23242 & new_n23500 ;
  assign new_n23502 = new_n23242 & ~new_n23500 ;
  assign new_n23503 = ~new_n23501 & ~new_n23502 ;
  assign new_n23504 = pi462 & new_n2071 ;
  assign new_n23505 = ~new_n23253 & new_n23494 ;
  assign new_n23506 = ~new_n23498 & ~new_n23505 ;
  assign new_n23507 = new_n23251 & ~new_n23506 ;
  assign new_n23508 = new_n23253 & new_n23494 ;
  assign new_n23509 = ~new_n23495 & ~new_n23508 ;
  assign new_n23510 = ~new_n23251 & ~new_n23509 ;
  assign new_n23511 = ~new_n23507 & ~new_n23510 ;
  assign new_n23512 = ~new_n23242 & new_n23511 ;
  assign new_n23513 = new_n23242 & ~new_n23511 ;
  assign new_n23514 = ~new_n23512 & ~new_n23513 ;
  assign new_n23515 = pi461 & new_n2071 ;
  assign new_n23516 = ~new_n23255 & new_n23488 ;
  assign new_n23517 = ~new_n23492 & ~new_n23516 ;
  assign new_n23518 = new_n23254 & ~new_n23517 ;
  assign new_n23519 = new_n23255 & new_n23488 ;
  assign new_n23520 = ~new_n23489 & ~new_n23519 ;
  assign new_n23521 = ~new_n23254 & ~new_n23520 ;
  assign new_n23522 = ~new_n23518 & ~new_n23521 ;
  assign new_n23523 = ~new_n23242 & new_n23522 ;
  assign new_n23524 = new_n23242 & ~new_n23522 ;
  assign new_n23525 = ~new_n23523 & ~new_n23524 ;
  assign new_n23526 = pi460 & new_n2071 ;
  assign new_n23527 = ~new_n23257 & new_n23482 ;
  assign new_n23528 = ~new_n23486 & ~new_n23527 ;
  assign new_n23529 = new_n23256 & ~new_n23528 ;
  assign new_n23530 = new_n23257 & new_n23482 ;
  assign new_n23531 = ~new_n23483 & ~new_n23530 ;
  assign new_n23532 = ~new_n23256 & ~new_n23531 ;
  assign new_n23533 = ~new_n23529 & ~new_n23532 ;
  assign new_n23534 = ~new_n23242 & new_n23533 ;
  assign new_n23535 = new_n23242 & ~new_n23533 ;
  assign new_n23536 = ~new_n23534 & ~new_n23535 ;
  assign new_n23537 = pi459 & new_n2071 ;
  assign new_n23538 = ~new_n23259 & new_n23476 ;
  assign new_n23539 = ~new_n23480 & ~new_n23538 ;
  assign new_n23540 = new_n23258 & ~new_n23539 ;
  assign new_n23541 = new_n23259 & new_n23476 ;
  assign new_n23542 = ~new_n23477 & ~new_n23541 ;
  assign new_n23543 = ~new_n23258 & ~new_n23542 ;
  assign new_n23544 = ~new_n23540 & ~new_n23543 ;
  assign new_n23545 = ~new_n23242 & new_n23544 ;
  assign new_n23546 = new_n23242 & ~new_n23544 ;
  assign new_n23547 = ~new_n23545 & ~new_n23546 ;
  assign new_n23548 = pi458 & new_n2071 ;
  assign new_n23549 = ~new_n23261 & new_n23470 ;
  assign new_n23550 = ~new_n23474 & ~new_n23549 ;
  assign new_n23551 = new_n23260 & ~new_n23550 ;
  assign new_n23552 = new_n23261 & new_n23470 ;
  assign new_n23553 = ~new_n23471 & ~new_n23552 ;
  assign new_n23554 = ~new_n23260 & ~new_n23553 ;
  assign new_n23555 = ~new_n23551 & ~new_n23554 ;
  assign new_n23556 = ~new_n23242 & new_n23555 ;
  assign new_n23557 = new_n23242 & ~new_n23555 ;
  assign new_n23558 = ~new_n23556 & ~new_n23557 ;
  assign new_n23559 = pi457 & new_n2071 ;
  assign new_n23560 = ~new_n23263 & new_n23464 ;
  assign new_n23561 = ~new_n23468 & ~new_n23560 ;
  assign new_n23562 = new_n23262 & ~new_n23561 ;
  assign new_n23563 = new_n23263 & new_n23464 ;
  assign new_n23564 = ~new_n23465 & ~new_n23563 ;
  assign new_n23565 = ~new_n23262 & ~new_n23564 ;
  assign new_n23566 = ~new_n23562 & ~new_n23565 ;
  assign new_n23567 = ~new_n23242 & new_n23566 ;
  assign new_n23568 = new_n23242 & ~new_n23566 ;
  assign new_n23569 = ~new_n23567 & ~new_n23568 ;
  assign new_n23570 = pi456 & new_n2071 ;
  assign new_n23571 = ~new_n23265 & new_n23458 ;
  assign new_n23572 = ~new_n23462 & ~new_n23571 ;
  assign new_n23573 = new_n23264 & ~new_n23572 ;
  assign new_n23574 = new_n23265 & new_n23458 ;
  assign new_n23575 = ~new_n23459 & ~new_n23574 ;
  assign new_n23576 = ~new_n23264 & ~new_n23575 ;
  assign new_n23577 = ~new_n23573 & ~new_n23576 ;
  assign new_n23578 = ~new_n23242 & new_n23577 ;
  assign new_n23579 = new_n23242 & ~new_n23577 ;
  assign new_n23580 = ~new_n23578 & ~new_n23579 ;
  assign new_n23581 = pi455 & new_n2071 ;
  assign new_n23582 = ~new_n23267 & new_n23452 ;
  assign new_n23583 = ~new_n23456 & ~new_n23582 ;
  assign new_n23584 = new_n23266 & ~new_n23583 ;
  assign new_n23585 = new_n23267 & new_n23452 ;
  assign new_n23586 = ~new_n23453 & ~new_n23585 ;
  assign new_n23587 = ~new_n23266 & ~new_n23586 ;
  assign new_n23588 = ~new_n23584 & ~new_n23587 ;
  assign new_n23589 = ~new_n23242 & new_n23588 ;
  assign new_n23590 = new_n23242 & ~new_n23588 ;
  assign new_n23591 = ~new_n23589 & ~new_n23590 ;
  assign new_n23592 = pi454 & new_n2071 ;
  assign new_n23593 = ~new_n23269 & new_n23446 ;
  assign new_n23594 = ~new_n23450 & ~new_n23593 ;
  assign new_n23595 = new_n23268 & ~new_n23594 ;
  assign new_n23596 = new_n23269 & new_n23446 ;
  assign new_n23597 = ~new_n23447 & ~new_n23596 ;
  assign new_n23598 = ~new_n23268 & ~new_n23597 ;
  assign new_n23599 = ~new_n23595 & ~new_n23598 ;
  assign new_n23600 = ~new_n23242 & new_n23599 ;
  assign new_n23601 = new_n23242 & ~new_n23599 ;
  assign new_n23602 = ~new_n23600 & ~new_n23601 ;
  assign new_n23603 = pi453 & new_n2071 ;
  assign new_n23604 = ~new_n23271 & new_n23440 ;
  assign new_n23605 = ~new_n23444 & ~new_n23604 ;
  assign new_n23606 = new_n23270 & ~new_n23605 ;
  assign new_n23607 = new_n23271 & new_n23440 ;
  assign new_n23608 = ~new_n23441 & ~new_n23607 ;
  assign new_n23609 = ~new_n23270 & ~new_n23608 ;
  assign new_n23610 = ~new_n23606 & ~new_n23609 ;
  assign new_n23611 = ~new_n23242 & new_n23610 ;
  assign new_n23612 = new_n23242 & ~new_n23610 ;
  assign new_n23613 = ~new_n23611 & ~new_n23612 ;
  assign new_n23614 = pi452 & new_n2071 ;
  assign new_n23615 = ~new_n23273 & new_n23434 ;
  assign new_n23616 = ~new_n23438 & ~new_n23615 ;
  assign new_n23617 = new_n23272 & ~new_n23616 ;
  assign new_n23618 = new_n23273 & new_n23434 ;
  assign new_n23619 = ~new_n23435 & ~new_n23618 ;
  assign new_n23620 = ~new_n23272 & ~new_n23619 ;
  assign new_n23621 = ~new_n23617 & ~new_n23620 ;
  assign new_n23622 = ~new_n23242 & new_n23621 ;
  assign new_n23623 = new_n23242 & ~new_n23621 ;
  assign new_n23624 = ~new_n23622 & ~new_n23623 ;
  assign new_n23625 = pi451 & new_n2071 ;
  assign new_n23626 = ~new_n23275 & new_n23428 ;
  assign new_n23627 = ~new_n23432 & ~new_n23626 ;
  assign new_n23628 = new_n23274 & ~new_n23627 ;
  assign new_n23629 = new_n23275 & new_n23428 ;
  assign new_n23630 = ~new_n23429 & ~new_n23629 ;
  assign new_n23631 = ~new_n23274 & ~new_n23630 ;
  assign new_n23632 = ~new_n23628 & ~new_n23631 ;
  assign new_n23633 = ~new_n23242 & new_n23632 ;
  assign new_n23634 = new_n23242 & ~new_n23632 ;
  assign new_n23635 = ~new_n23633 & ~new_n23634 ;
  assign new_n23636 = pi450 & new_n2071 ;
  assign new_n23637 = ~new_n23277 & new_n23422 ;
  assign new_n23638 = ~new_n23426 & ~new_n23637 ;
  assign new_n23639 = new_n23276 & ~new_n23638 ;
  assign new_n23640 = new_n23277 & new_n23422 ;
  assign new_n23641 = ~new_n23423 & ~new_n23640 ;
  assign new_n23642 = ~new_n23276 & ~new_n23641 ;
  assign new_n23643 = ~new_n23639 & ~new_n23642 ;
  assign new_n23644 = ~new_n23242 & new_n23643 ;
  assign new_n23645 = new_n23242 & ~new_n23643 ;
  assign new_n23646 = ~new_n23644 & ~new_n23645 ;
  assign new_n23647 = pi449 & new_n2071 ;
  assign new_n23648 = ~new_n23279 & new_n23416 ;
  assign new_n23649 = ~new_n23420 & ~new_n23648 ;
  assign new_n23650 = new_n23278 & ~new_n23649 ;
  assign new_n23651 = new_n23279 & new_n23416 ;
  assign new_n23652 = ~new_n23417 & ~new_n23651 ;
  assign new_n23653 = ~new_n23278 & ~new_n23652 ;
  assign new_n23654 = ~new_n23650 & ~new_n23653 ;
  assign new_n23655 = ~new_n23242 & new_n23654 ;
  assign new_n23656 = new_n23242 & ~new_n23654 ;
  assign new_n23657 = ~new_n23655 & ~new_n23656 ;
  assign new_n23658 = pi448 & new_n2071 ;
  assign new_n23659 = ~new_n23281 & new_n23410 ;
  assign new_n23660 = ~new_n23414 & ~new_n23659 ;
  assign new_n23661 = new_n23280 & ~new_n23660 ;
  assign new_n23662 = new_n23281 & new_n23410 ;
  assign new_n23663 = ~new_n23411 & ~new_n23662 ;
  assign new_n23664 = ~new_n23280 & ~new_n23663 ;
  assign new_n23665 = ~new_n23661 & ~new_n23664 ;
  assign new_n23666 = ~new_n23242 & new_n23665 ;
  assign new_n23667 = new_n23242 & ~new_n23665 ;
  assign new_n23668 = ~new_n23666 & ~new_n23667 ;
  assign new_n23669 = ~new_n23283 & new_n23404 ;
  assign new_n23670 = ~new_n23408 & ~new_n23669 ;
  assign new_n23671 = new_n23282 & ~new_n23670 ;
  assign new_n23672 = new_n23283 & new_n23404 ;
  assign new_n23673 = ~new_n23405 & ~new_n23672 ;
  assign new_n23674 = ~new_n23282 & ~new_n23673 ;
  assign new_n23675 = ~new_n23671 & ~new_n23674 ;
  assign new_n23676 = ~new_n23242 & new_n23675 ;
  assign new_n23677 = new_n23242 & ~new_n23675 ;
  assign new_n23678 = ~new_n23676 & ~new_n23677 ;
  assign new_n23679 = lo1123 & ~new_n2071 ;
  assign new_n23680 = ~new_n2074 & new_n23679 ;
  assign new_n23681 = pi447 & new_n2071 ;
  assign new_n23682 = ~new_n23680 & ~new_n23681 ;
  assign new_n23683 = ~new_n23291 & new_n23398 ;
  assign new_n23684 = ~new_n23402 & ~new_n23683 ;
  assign new_n23685 = new_n23287 & ~new_n23684 ;
  assign new_n23686 = new_n23291 & new_n23398 ;
  assign new_n23687 = ~new_n23399 & ~new_n23686 ;
  assign new_n23688 = ~new_n23287 & ~new_n23687 ;
  assign new_n23689 = ~new_n23685 & ~new_n23688 ;
  assign new_n23690 = ~new_n23242 & new_n23689 ;
  assign new_n23691 = new_n23242 & ~new_n23689 ;
  assign new_n23692 = ~new_n23690 & ~new_n23691 ;
  assign new_n23693 = ~new_n23293 & new_n23392 ;
  assign new_n23694 = ~new_n23396 & ~new_n23693 ;
  assign new_n23695 = new_n23292 & ~new_n23694 ;
  assign new_n23696 = new_n23293 & new_n23392 ;
  assign new_n23697 = ~new_n23393 & ~new_n23696 ;
  assign new_n23698 = ~new_n23292 & ~new_n23697 ;
  assign new_n23699 = ~new_n23695 & ~new_n23698 ;
  assign new_n23700 = ~new_n23242 & new_n23699 ;
  assign new_n23701 = new_n23242 & ~new_n23699 ;
  assign new_n23702 = ~new_n23700 & ~new_n23701 ;
  assign new_n23703 = ~new_n23295 & new_n23386 ;
  assign new_n23704 = ~new_n23390 & ~new_n23703 ;
  assign new_n23705 = new_n23294 & ~new_n23704 ;
  assign new_n23706 = new_n23295 & new_n23386 ;
  assign new_n23707 = ~new_n23387 & ~new_n23706 ;
  assign new_n23708 = ~new_n23294 & ~new_n23707 ;
  assign new_n23709 = ~new_n23705 & ~new_n23708 ;
  assign new_n23710 = ~new_n23242 & new_n23709 ;
  assign new_n23711 = new_n23242 & ~new_n23709 ;
  assign new_n23712 = ~new_n23710 & ~new_n23711 ;
  assign new_n23713 = ~new_n23297 & new_n23380 ;
  assign new_n23714 = ~new_n23384 & ~new_n23713 ;
  assign new_n23715 = new_n23296 & ~new_n23714 ;
  assign new_n23716 = new_n23297 & new_n23380 ;
  assign new_n23717 = ~new_n23381 & ~new_n23716 ;
  assign new_n23718 = ~new_n23296 & ~new_n23717 ;
  assign new_n23719 = ~new_n23715 & ~new_n23718 ;
  assign new_n23720 = ~new_n23242 & new_n23719 ;
  assign new_n23721 = new_n23242 & ~new_n23719 ;
  assign new_n23722 = ~new_n23720 & ~new_n23721 ;
  assign new_n23723 = ~new_n23299 & new_n23374 ;
  assign new_n23724 = ~new_n23378 & ~new_n23723 ;
  assign new_n23725 = new_n23298 & ~new_n23724 ;
  assign new_n23726 = new_n23299 & new_n23374 ;
  assign new_n23727 = ~new_n23375 & ~new_n23726 ;
  assign new_n23728 = ~new_n23298 & ~new_n23727 ;
  assign new_n23729 = ~new_n23725 & ~new_n23728 ;
  assign new_n23730 = ~new_n23242 & new_n23729 ;
  assign new_n23731 = new_n23242 & ~new_n23729 ;
  assign new_n23732 = ~new_n23730 & ~new_n23731 ;
  assign new_n23733 = ~new_n23301 & new_n23368 ;
  assign new_n23734 = ~new_n23372 & ~new_n23733 ;
  assign new_n23735 = new_n23300 & ~new_n23734 ;
  assign new_n23736 = new_n23301 & new_n23368 ;
  assign new_n23737 = ~new_n23369 & ~new_n23736 ;
  assign new_n23738 = ~new_n23300 & ~new_n23737 ;
  assign new_n23739 = ~new_n23735 & ~new_n23738 ;
  assign new_n23740 = ~new_n23242 & new_n23739 ;
  assign new_n23741 = new_n23242 & ~new_n23739 ;
  assign new_n23742 = ~new_n23740 & ~new_n23741 ;
  assign new_n23743 = ~new_n23303 & new_n23362 ;
  assign new_n23744 = ~new_n23366 & ~new_n23743 ;
  assign new_n23745 = new_n23302 & ~new_n23744 ;
  assign new_n23746 = new_n23303 & new_n23362 ;
  assign new_n23747 = ~new_n23363 & ~new_n23746 ;
  assign new_n23748 = ~new_n23302 & ~new_n23747 ;
  assign new_n23749 = ~new_n23745 & ~new_n23748 ;
  assign new_n23750 = ~new_n23242 & new_n23749 ;
  assign new_n23751 = new_n23242 & ~new_n23749 ;
  assign new_n23752 = ~new_n23750 & ~new_n23751 ;
  assign new_n23753 = ~new_n23305 & new_n23356 ;
  assign new_n23754 = ~new_n23360 & ~new_n23753 ;
  assign new_n23755 = new_n23304 & ~new_n23754 ;
  assign new_n23756 = new_n23305 & new_n23356 ;
  assign new_n23757 = ~new_n23357 & ~new_n23756 ;
  assign new_n23758 = ~new_n23304 & ~new_n23757 ;
  assign new_n23759 = ~new_n23755 & ~new_n23758 ;
  assign new_n23760 = ~new_n23242 & new_n23759 ;
  assign new_n23761 = new_n23242 & ~new_n23759 ;
  assign new_n23762 = ~new_n23760 & ~new_n23761 ;
  assign new_n23763 = ~new_n23307 & new_n23350 ;
  assign new_n23764 = ~new_n23354 & ~new_n23763 ;
  assign new_n23765 = new_n23306 & ~new_n23764 ;
  assign new_n23766 = new_n23307 & new_n23350 ;
  assign new_n23767 = ~new_n23351 & ~new_n23766 ;
  assign new_n23768 = ~new_n23306 & ~new_n23767 ;
  assign new_n23769 = ~new_n23765 & ~new_n23768 ;
  assign new_n23770 = ~new_n23242 & new_n23769 ;
  assign new_n23771 = new_n23242 & ~new_n23769 ;
  assign new_n23772 = ~new_n23770 & ~new_n23771 ;
  assign new_n23773 = ~new_n23309 & new_n23344 ;
  assign new_n23774 = ~new_n23348 & ~new_n23773 ;
  assign new_n23775 = new_n23308 & ~new_n23774 ;
  assign new_n23776 = new_n23309 & new_n23344 ;
  assign new_n23777 = ~new_n23345 & ~new_n23776 ;
  assign new_n23778 = ~new_n23308 & ~new_n23777 ;
  assign new_n23779 = ~new_n23775 & ~new_n23778 ;
  assign new_n23780 = ~new_n23242 & new_n23779 ;
  assign new_n23781 = new_n23242 & ~new_n23779 ;
  assign new_n23782 = ~new_n23780 & ~new_n23781 ;
  assign new_n23783 = ~new_n23311 & new_n23338 ;
  assign new_n23784 = ~new_n23342 & ~new_n23783 ;
  assign new_n23785 = new_n23310 & ~new_n23784 ;
  assign new_n23786 = new_n23311 & new_n23338 ;
  assign new_n23787 = ~new_n23339 & ~new_n23786 ;
  assign new_n23788 = ~new_n23310 & ~new_n23787 ;
  assign new_n23789 = ~new_n23785 & ~new_n23788 ;
  assign new_n23790 = ~new_n23242 & new_n23789 ;
  assign new_n23791 = new_n23242 & ~new_n23789 ;
  assign new_n23792 = ~new_n23790 & ~new_n23791 ;
  assign new_n23793 = ~new_n23313 & new_n23332 ;
  assign new_n23794 = ~new_n23336 & ~new_n23793 ;
  assign new_n23795 = new_n23312 & ~new_n23794 ;
  assign new_n23796 = new_n23313 & new_n23332 ;
  assign new_n23797 = ~new_n23333 & ~new_n23796 ;
  assign new_n23798 = ~new_n23312 & ~new_n23797 ;
  assign new_n23799 = ~new_n23795 & ~new_n23798 ;
  assign new_n23800 = ~new_n23242 & new_n23799 ;
  assign new_n23801 = new_n23242 & ~new_n23799 ;
  assign new_n23802 = ~new_n23800 & ~new_n23801 ;
  assign new_n23803 = ~new_n23315 & new_n23326 ;
  assign new_n23804 = ~new_n23330 & ~new_n23803 ;
  assign new_n23805 = new_n23314 & ~new_n23804 ;
  assign new_n23806 = new_n23315 & new_n23326 ;
  assign new_n23807 = ~new_n23327 & ~new_n23806 ;
  assign new_n23808 = ~new_n23314 & ~new_n23807 ;
  assign new_n23809 = ~new_n23805 & ~new_n23808 ;
  assign new_n23810 = ~new_n23242 & new_n23809 ;
  assign new_n23811 = new_n23242 & ~new_n23809 ;
  assign new_n23812 = ~new_n23810 & ~new_n23811 ;
  assign new_n23813 = ~new_n23317 & ~new_n23320 ;
  assign new_n23814 = ~new_n23324 & ~new_n23813 ;
  assign new_n23815 = new_n23316 & ~new_n23814 ;
  assign new_n23816 = new_n23317 & ~new_n23320 ;
  assign new_n23817 = ~new_n23321 & ~new_n23816 ;
  assign new_n23818 = ~new_n23316 & ~new_n23817 ;
  assign new_n23819 = ~new_n23815 & ~new_n23818 ;
  assign new_n23820 = ~new_n23242 & new_n23819 ;
  assign new_n23821 = new_n23242 & ~new_n23819 ;
  assign new_n23822 = ~new_n23820 & ~new_n23821 ;
  assign new_n23823 = new_n23318 & ~new_n23319 ;
  assign new_n23824 = ~new_n23318 & new_n23319 ;
  assign new_n23825 = ~new_n23823 & ~new_n23824 ;
  assign new_n23826 = ~new_n23242 & new_n23825 ;
  assign new_n23827 = new_n23242 & ~new_n23825 ;
  assign new_n23828 = ~new_n23826 & ~new_n23827 ;
  assign new_n23829 = ~pi432 & new_n23242 ;
  assign new_n23830 = ~pi432 & ~new_n23829 ;
  assign new_n23831 = new_n23828 & ~new_n23830 ;
  assign new_n23832 = pi432 & new_n23242 ;
  assign new_n23833 = ~new_n23828 & new_n23832 ;
  assign new_n23834 = ~new_n23831 & ~new_n23833 ;
  assign new_n23835 = ~pi433 & ~new_n23834 ;
  assign new_n23836 = ~pi433 & ~new_n23835 ;
  assign new_n23837 = new_n23822 & ~new_n23836 ;
  assign new_n23838 = pi433 & ~new_n23834 ;
  assign new_n23839 = ~new_n23822 & new_n23838 ;
  assign new_n23840 = ~new_n23837 & ~new_n23839 ;
  assign new_n23841 = ~pi434 & ~new_n23840 ;
  assign new_n23842 = ~pi434 & ~new_n23841 ;
  assign new_n23843 = new_n23812 & ~new_n23842 ;
  assign new_n23844 = pi434 & ~new_n23840 ;
  assign new_n23845 = ~new_n23812 & new_n23844 ;
  assign new_n23846 = ~new_n23843 & ~new_n23845 ;
  assign new_n23847 = ~pi435 & ~new_n23846 ;
  assign new_n23848 = ~pi435 & ~new_n23847 ;
  assign new_n23849 = new_n23802 & ~new_n23848 ;
  assign new_n23850 = pi435 & ~new_n23846 ;
  assign new_n23851 = ~new_n23802 & new_n23850 ;
  assign new_n23852 = ~new_n23849 & ~new_n23851 ;
  assign new_n23853 = ~pi436 & ~new_n23852 ;
  assign new_n23854 = ~pi436 & ~new_n23853 ;
  assign new_n23855 = new_n23792 & ~new_n23854 ;
  assign new_n23856 = pi436 & ~new_n23852 ;
  assign new_n23857 = ~new_n23792 & new_n23856 ;
  assign new_n23858 = ~new_n23855 & ~new_n23857 ;
  assign new_n23859 = ~pi437 & ~new_n23858 ;
  assign new_n23860 = ~pi437 & ~new_n23859 ;
  assign new_n23861 = new_n23782 & ~new_n23860 ;
  assign new_n23862 = pi437 & ~new_n23858 ;
  assign new_n23863 = ~new_n23782 & new_n23862 ;
  assign new_n23864 = ~new_n23861 & ~new_n23863 ;
  assign new_n23865 = ~pi438 & ~new_n23864 ;
  assign new_n23866 = ~pi438 & ~new_n23865 ;
  assign new_n23867 = new_n23772 & ~new_n23866 ;
  assign new_n23868 = pi438 & ~new_n23864 ;
  assign new_n23869 = ~new_n23772 & new_n23868 ;
  assign new_n23870 = ~new_n23867 & ~new_n23869 ;
  assign new_n23871 = ~pi439 & ~new_n23870 ;
  assign new_n23872 = ~pi439 & ~new_n23871 ;
  assign new_n23873 = new_n23762 & ~new_n23872 ;
  assign new_n23874 = pi439 & ~new_n23870 ;
  assign new_n23875 = ~new_n23762 & new_n23874 ;
  assign new_n23876 = ~new_n23873 & ~new_n23875 ;
  assign new_n23877 = ~pi440 & ~new_n23876 ;
  assign new_n23878 = ~pi440 & ~new_n23877 ;
  assign new_n23879 = new_n23752 & ~new_n23878 ;
  assign new_n23880 = pi440 & ~new_n23876 ;
  assign new_n23881 = ~new_n23752 & new_n23880 ;
  assign new_n23882 = ~new_n23879 & ~new_n23881 ;
  assign new_n23883 = ~pi441 & ~new_n23882 ;
  assign new_n23884 = ~pi441 & ~new_n23883 ;
  assign new_n23885 = new_n23742 & ~new_n23884 ;
  assign new_n23886 = pi441 & ~new_n23882 ;
  assign new_n23887 = ~new_n23742 & new_n23886 ;
  assign new_n23888 = ~new_n23885 & ~new_n23887 ;
  assign new_n23889 = ~pi442 & ~new_n23888 ;
  assign new_n23890 = ~pi442 & ~new_n23889 ;
  assign new_n23891 = new_n23732 & ~new_n23890 ;
  assign new_n23892 = pi442 & ~new_n23888 ;
  assign new_n23893 = ~new_n23732 & new_n23892 ;
  assign new_n23894 = ~new_n23891 & ~new_n23893 ;
  assign new_n23895 = ~pi443 & ~new_n23894 ;
  assign new_n23896 = ~pi443 & ~new_n23895 ;
  assign new_n23897 = new_n23722 & ~new_n23896 ;
  assign new_n23898 = pi443 & ~new_n23894 ;
  assign new_n23899 = ~new_n23722 & new_n23898 ;
  assign new_n23900 = ~new_n23897 & ~new_n23899 ;
  assign new_n23901 = ~pi444 & ~new_n23900 ;
  assign new_n23902 = ~pi444 & ~new_n23901 ;
  assign new_n23903 = new_n23712 & ~new_n23902 ;
  assign new_n23904 = pi444 & ~new_n23900 ;
  assign new_n23905 = ~new_n23712 & new_n23904 ;
  assign new_n23906 = ~new_n23903 & ~new_n23905 ;
  assign new_n23907 = ~pi445 & ~new_n23906 ;
  assign new_n23908 = ~pi445 & ~new_n23907 ;
  assign new_n23909 = new_n23702 & ~new_n23908 ;
  assign new_n23910 = pi445 & ~new_n23906 ;
  assign new_n23911 = ~new_n23702 & new_n23910 ;
  assign new_n23912 = ~new_n23909 & ~new_n23911 ;
  assign new_n23913 = ~pi446 & ~new_n23912 ;
  assign new_n23914 = ~pi446 & ~new_n23913 ;
  assign new_n23915 = new_n23692 & ~new_n23914 ;
  assign new_n23916 = pi446 & ~new_n23912 ;
  assign new_n23917 = ~new_n23692 & new_n23916 ;
  assign new_n23918 = ~new_n23915 & ~new_n23917 ;
  assign new_n23919 = new_n23682 & ~new_n23918 ;
  assign new_n23920 = new_n23682 & ~new_n23919 ;
  assign new_n23921 = new_n23678 & ~new_n23920 ;
  assign new_n23922 = ~new_n23682 & ~new_n23918 ;
  assign new_n23923 = ~new_n23678 & new_n23922 ;
  assign new_n23924 = ~new_n23921 & ~new_n23923 ;
  assign new_n23925 = ~new_n23668 & ~new_n23924 ;
  assign new_n23926 = ~new_n23668 & ~new_n23925 ;
  assign new_n23927 = new_n23658 & ~new_n23926 ;
  assign new_n23928 = new_n23668 & ~new_n23924 ;
  assign new_n23929 = ~new_n23658 & new_n23928 ;
  assign new_n23930 = ~new_n23927 & ~new_n23929 ;
  assign new_n23931 = ~new_n23657 & ~new_n23930 ;
  assign new_n23932 = ~new_n23657 & ~new_n23931 ;
  assign new_n23933 = new_n23647 & ~new_n23932 ;
  assign new_n23934 = new_n23657 & ~new_n23930 ;
  assign new_n23935 = ~new_n23647 & new_n23934 ;
  assign new_n23936 = ~new_n23933 & ~new_n23935 ;
  assign new_n23937 = ~new_n23646 & ~new_n23936 ;
  assign new_n23938 = ~new_n23646 & ~new_n23937 ;
  assign new_n23939 = new_n23636 & ~new_n23938 ;
  assign new_n23940 = new_n23646 & ~new_n23936 ;
  assign new_n23941 = ~new_n23636 & new_n23940 ;
  assign new_n23942 = ~new_n23939 & ~new_n23941 ;
  assign new_n23943 = ~new_n23635 & ~new_n23942 ;
  assign new_n23944 = ~new_n23635 & ~new_n23943 ;
  assign new_n23945 = new_n23625 & ~new_n23944 ;
  assign new_n23946 = new_n23635 & ~new_n23942 ;
  assign new_n23947 = ~new_n23625 & new_n23946 ;
  assign new_n23948 = ~new_n23945 & ~new_n23947 ;
  assign new_n23949 = ~new_n23624 & ~new_n23948 ;
  assign new_n23950 = ~new_n23624 & ~new_n23949 ;
  assign new_n23951 = new_n23614 & ~new_n23950 ;
  assign new_n23952 = new_n23624 & ~new_n23948 ;
  assign new_n23953 = ~new_n23614 & new_n23952 ;
  assign new_n23954 = ~new_n23951 & ~new_n23953 ;
  assign new_n23955 = ~new_n23613 & ~new_n23954 ;
  assign new_n23956 = ~new_n23613 & ~new_n23955 ;
  assign new_n23957 = new_n23603 & ~new_n23956 ;
  assign new_n23958 = new_n23613 & ~new_n23954 ;
  assign new_n23959 = ~new_n23603 & new_n23958 ;
  assign new_n23960 = ~new_n23957 & ~new_n23959 ;
  assign new_n23961 = ~new_n23602 & ~new_n23960 ;
  assign new_n23962 = ~new_n23602 & ~new_n23961 ;
  assign new_n23963 = new_n23592 & ~new_n23962 ;
  assign new_n23964 = new_n23602 & ~new_n23960 ;
  assign new_n23965 = ~new_n23592 & new_n23964 ;
  assign new_n23966 = ~new_n23963 & ~new_n23965 ;
  assign new_n23967 = ~new_n23591 & ~new_n23966 ;
  assign new_n23968 = ~new_n23591 & ~new_n23967 ;
  assign new_n23969 = new_n23581 & ~new_n23968 ;
  assign new_n23970 = new_n23591 & ~new_n23966 ;
  assign new_n23971 = ~new_n23581 & new_n23970 ;
  assign new_n23972 = ~new_n23969 & ~new_n23971 ;
  assign new_n23973 = ~new_n23580 & ~new_n23972 ;
  assign new_n23974 = ~new_n23580 & ~new_n23973 ;
  assign new_n23975 = new_n23570 & ~new_n23974 ;
  assign new_n23976 = new_n23580 & ~new_n23972 ;
  assign new_n23977 = ~new_n23570 & new_n23976 ;
  assign new_n23978 = ~new_n23975 & ~new_n23977 ;
  assign new_n23979 = ~new_n23569 & ~new_n23978 ;
  assign new_n23980 = ~new_n23569 & ~new_n23979 ;
  assign new_n23981 = new_n23559 & ~new_n23980 ;
  assign new_n23982 = new_n23569 & ~new_n23978 ;
  assign new_n23983 = ~new_n23559 & new_n23982 ;
  assign new_n23984 = ~new_n23981 & ~new_n23983 ;
  assign new_n23985 = ~new_n23558 & ~new_n23984 ;
  assign new_n23986 = ~new_n23558 & ~new_n23985 ;
  assign new_n23987 = new_n23548 & ~new_n23986 ;
  assign new_n23988 = new_n23558 & ~new_n23984 ;
  assign new_n23989 = ~new_n23548 & new_n23988 ;
  assign new_n23990 = ~new_n23987 & ~new_n23989 ;
  assign new_n23991 = ~new_n23547 & ~new_n23990 ;
  assign new_n23992 = ~new_n23547 & ~new_n23991 ;
  assign new_n23993 = new_n23537 & ~new_n23992 ;
  assign new_n23994 = new_n23547 & ~new_n23990 ;
  assign new_n23995 = ~new_n23537 & new_n23994 ;
  assign new_n23996 = ~new_n23993 & ~new_n23995 ;
  assign new_n23997 = ~new_n23536 & ~new_n23996 ;
  assign new_n23998 = ~new_n23536 & ~new_n23997 ;
  assign new_n23999 = new_n23526 & ~new_n23998 ;
  assign new_n24000 = new_n23536 & ~new_n23996 ;
  assign new_n24001 = ~new_n23526 & new_n24000 ;
  assign new_n24002 = ~new_n23999 & ~new_n24001 ;
  assign new_n24003 = ~new_n23525 & ~new_n24002 ;
  assign new_n24004 = ~new_n23525 & ~new_n24003 ;
  assign new_n24005 = new_n23515 & ~new_n24004 ;
  assign new_n24006 = new_n23525 & ~new_n24002 ;
  assign new_n24007 = ~new_n23515 & new_n24006 ;
  assign new_n24008 = ~new_n24005 & ~new_n24007 ;
  assign new_n24009 = ~new_n23514 & ~new_n24008 ;
  assign new_n24010 = ~new_n23514 & ~new_n24009 ;
  assign new_n24011 = new_n23504 & ~new_n24010 ;
  assign new_n24012 = new_n23514 & ~new_n24008 ;
  assign new_n24013 = ~new_n23504 & new_n24012 ;
  assign new_n24014 = ~new_n24011 & ~new_n24013 ;
  assign new_n24015 = ~new_n23503 & ~new_n24014 ;
  assign new_n24016 = ~new_n23503 & ~new_n24015 ;
  assign new_n24017 = new_n23250 & ~new_n24016 ;
  assign new_n24018 = new_n23503 & ~new_n24014 ;
  assign new_n24019 = ~new_n23250 & new_n24018 ;
  assign new_n24020 = ~new_n24017 & ~new_n24019 ;
  assign new_n24021 = new_n23242 & new_n24020 ;
  assign new_n24022 = ~new_n23242 & ~new_n24020 ;
  assign new_n24023 = ~new_n24021 & ~new_n24022 ;
  assign new_n24024 = new_n23240 & ~new_n24023 ;
  assign new_n24025 = ~new_n2138 & ~new_n24023 ;
  assign new_n24026 = ~new_n24024 & ~new_n24025 ;
  assign new_n24027 = ~lo1408 & ~new_n24026 ;
  assign new_n24028 = new_n2069 & new_n21021 ;
  assign new_n24029 = lo1408 & new_n24028 ;
  assign new_n24030 = lo1330 & new_n24028 ;
  assign new_n24031 = ~new_n23503 & new_n24014 ;
  assign new_n24032 = ~new_n24018 & ~new_n24031 ;
  assign new_n24033 = new_n23250 & ~new_n24032 ;
  assign new_n24034 = new_n23503 & new_n24014 ;
  assign new_n24035 = ~new_n24015 & ~new_n24034 ;
  assign new_n24036 = ~new_n23250 & ~new_n24035 ;
  assign new_n24037 = ~new_n24033 & ~new_n24036 ;
  assign new_n24038 = ~new_n2138 & ~new_n24037 ;
  assign new_n24039 = ~new_n24024 & ~new_n24038 ;
  assign new_n24040 = lo1405 & new_n24028 ;
  assign new_n24041 = ~new_n23514 & new_n24008 ;
  assign new_n24042 = ~new_n24012 & ~new_n24041 ;
  assign new_n24043 = new_n23504 & ~new_n24042 ;
  assign new_n24044 = new_n23514 & new_n24008 ;
  assign new_n24045 = ~new_n24009 & ~new_n24044 ;
  assign new_n24046 = ~new_n23504 & ~new_n24045 ;
  assign new_n24047 = ~new_n24043 & ~new_n24046 ;
  assign new_n24048 = ~new_n2138 & ~new_n24047 ;
  assign new_n24049 = ~new_n24024 & ~new_n24048 ;
  assign new_n24050 = lo1353 & new_n24028 ;
  assign new_n24051 = ~new_n23525 & new_n24002 ;
  assign new_n24052 = ~new_n24006 & ~new_n24051 ;
  assign new_n24053 = new_n23515 & ~new_n24052 ;
  assign new_n24054 = new_n23525 & new_n24002 ;
  assign new_n24055 = ~new_n24003 & ~new_n24054 ;
  assign new_n24056 = ~new_n23515 & ~new_n24055 ;
  assign new_n24057 = ~new_n24053 & ~new_n24056 ;
  assign new_n24058 = ~new_n2138 & ~new_n24057 ;
  assign new_n24059 = ~new_n24024 & ~new_n24058 ;
  assign new_n24060 = lo1399 & new_n24028 ;
  assign new_n24061 = ~new_n23536 & new_n23996 ;
  assign new_n24062 = ~new_n24000 & ~new_n24061 ;
  assign new_n24063 = new_n23526 & ~new_n24062 ;
  assign new_n24064 = new_n23536 & new_n23996 ;
  assign new_n24065 = ~new_n23997 & ~new_n24064 ;
  assign new_n24066 = ~new_n23526 & ~new_n24065 ;
  assign new_n24067 = ~new_n24063 & ~new_n24066 ;
  assign new_n24068 = ~new_n2138 & ~new_n24067 ;
  assign new_n24069 = ~new_n24024 & ~new_n24068 ;
  assign new_n24070 = lo1414 & new_n24028 ;
  assign new_n24071 = ~new_n23547 & new_n23990 ;
  assign new_n24072 = ~new_n23994 & ~new_n24071 ;
  assign new_n24073 = new_n23537 & ~new_n24072 ;
  assign new_n24074 = new_n23547 & new_n23990 ;
  assign new_n24075 = ~new_n23991 & ~new_n24074 ;
  assign new_n24076 = ~new_n23537 & ~new_n24075 ;
  assign new_n24077 = ~new_n24073 & ~new_n24076 ;
  assign new_n24078 = ~new_n2138 & ~new_n24077 ;
  assign new_n24079 = ~new_n24024 & ~new_n24078 ;
  assign new_n24080 = lo1402 & new_n24028 ;
  assign new_n24081 = ~new_n23558 & new_n23984 ;
  assign new_n24082 = ~new_n23988 & ~new_n24081 ;
  assign new_n24083 = new_n23548 & ~new_n24082 ;
  assign new_n24084 = new_n23558 & new_n23984 ;
  assign new_n24085 = ~new_n23985 & ~new_n24084 ;
  assign new_n24086 = ~new_n23548 & ~new_n24085 ;
  assign new_n24087 = ~new_n24083 & ~new_n24086 ;
  assign new_n24088 = ~new_n2138 & ~new_n24087 ;
  assign new_n24089 = ~new_n24024 & ~new_n24088 ;
  assign new_n24090 = lo1417 & new_n24028 ;
  assign new_n24091 = ~new_n23569 & new_n23978 ;
  assign new_n24092 = ~new_n23982 & ~new_n24091 ;
  assign new_n24093 = new_n23559 & ~new_n24092 ;
  assign new_n24094 = new_n23569 & new_n23978 ;
  assign new_n24095 = ~new_n23979 & ~new_n24094 ;
  assign new_n24096 = ~new_n23559 & ~new_n24095 ;
  assign new_n24097 = ~new_n24093 & ~new_n24096 ;
  assign new_n24098 = ~new_n2138 & ~new_n24097 ;
  assign new_n24099 = ~new_n24024 & ~new_n24098 ;
  assign new_n24100 = lo1393 & new_n24028 ;
  assign new_n24101 = ~new_n23580 & new_n23972 ;
  assign new_n24102 = ~new_n23976 & ~new_n24101 ;
  assign new_n24103 = new_n23570 & ~new_n24102 ;
  assign new_n24104 = new_n23580 & new_n23972 ;
  assign new_n24105 = ~new_n23973 & ~new_n24104 ;
  assign new_n24106 = ~new_n23570 & ~new_n24105 ;
  assign new_n24107 = ~new_n24103 & ~new_n24106 ;
  assign new_n24108 = ~new_n2138 & ~new_n24107 ;
  assign new_n24109 = ~new_n24024 & ~new_n24108 ;
  assign new_n24110 = lo1356 & new_n24028 ;
  assign new_n24111 = ~new_n23591 & new_n23966 ;
  assign new_n24112 = ~new_n23970 & ~new_n24111 ;
  assign new_n24113 = new_n23581 & ~new_n24112 ;
  assign new_n24114 = new_n23591 & new_n23966 ;
  assign new_n24115 = ~new_n23967 & ~new_n24114 ;
  assign new_n24116 = ~new_n23581 & ~new_n24115 ;
  assign new_n24117 = ~new_n24113 & ~new_n24116 ;
  assign new_n24118 = ~new_n2138 & ~new_n24117 ;
  assign new_n24119 = ~new_n24024 & ~new_n24118 ;
  assign new_n24120 = lo1341 & new_n24028 ;
  assign new_n24121 = ~new_n23602 & new_n23960 ;
  assign new_n24122 = ~new_n23964 & ~new_n24121 ;
  assign new_n24123 = new_n23592 & ~new_n24122 ;
  assign new_n24124 = new_n23602 & new_n23960 ;
  assign new_n24125 = ~new_n23961 & ~new_n24124 ;
  assign new_n24126 = ~new_n23592 & ~new_n24125 ;
  assign new_n24127 = ~new_n24123 & ~new_n24126 ;
  assign new_n24128 = ~new_n2138 & ~new_n24127 ;
  assign new_n24129 = ~new_n24024 & ~new_n24128 ;
  assign new_n24130 = lo1299 & new_n24028 ;
  assign new_n24131 = ~new_n23613 & new_n23954 ;
  assign new_n24132 = ~new_n23958 & ~new_n24131 ;
  assign new_n24133 = new_n23603 & ~new_n24132 ;
  assign new_n24134 = new_n23613 & new_n23954 ;
  assign new_n24135 = ~new_n23955 & ~new_n24134 ;
  assign new_n24136 = ~new_n23603 & ~new_n24135 ;
  assign new_n24137 = ~new_n24133 & ~new_n24136 ;
  assign new_n24138 = ~new_n2138 & ~new_n24137 ;
  assign new_n24139 = ~new_n24024 & ~new_n24138 ;
  assign new_n24140 = lo1377 & new_n24028 ;
  assign new_n24141 = ~new_n23624 & new_n23948 ;
  assign new_n24142 = ~new_n23952 & ~new_n24141 ;
  assign new_n24143 = new_n23614 & ~new_n24142 ;
  assign new_n24144 = new_n23624 & new_n23948 ;
  assign new_n24145 = ~new_n23949 & ~new_n24144 ;
  assign new_n24146 = ~new_n23614 & ~new_n24145 ;
  assign new_n24147 = ~new_n24143 & ~new_n24146 ;
  assign new_n24148 = ~new_n2138 & ~new_n24147 ;
  assign new_n24149 = ~new_n24024 & ~new_n24148 ;
  assign new_n24150 = lo1371 & new_n24028 ;
  assign new_n24151 = ~new_n23635 & new_n23942 ;
  assign new_n24152 = ~new_n23946 & ~new_n24151 ;
  assign new_n24153 = new_n23625 & ~new_n24152 ;
  assign new_n24154 = new_n23635 & new_n23942 ;
  assign new_n24155 = ~new_n23943 & ~new_n24154 ;
  assign new_n24156 = ~new_n23625 & ~new_n24155 ;
  assign new_n24157 = ~new_n24153 & ~new_n24156 ;
  assign new_n24158 = ~new_n2138 & ~new_n24157 ;
  assign new_n24159 = ~new_n24024 & ~new_n24158 ;
  assign new_n24160 = lo1389 & new_n24028 ;
  assign new_n24161 = ~new_n23646 & new_n23936 ;
  assign new_n24162 = ~new_n23940 & ~new_n24161 ;
  assign new_n24163 = new_n23636 & ~new_n24162 ;
  assign new_n24164 = new_n23646 & new_n23936 ;
  assign new_n24165 = ~new_n23937 & ~new_n24164 ;
  assign new_n24166 = ~new_n23636 & ~new_n24165 ;
  assign new_n24167 = ~new_n24163 & ~new_n24166 ;
  assign new_n24168 = ~new_n2138 & ~new_n24167 ;
  assign new_n24169 = ~new_n24024 & ~new_n24168 ;
  assign new_n24170 = lo1364 & new_n24028 ;
  assign new_n24171 = ~new_n23657 & new_n23930 ;
  assign new_n24172 = ~new_n23934 & ~new_n24171 ;
  assign new_n24173 = new_n23647 & ~new_n24172 ;
  assign new_n24174 = new_n23657 & new_n23930 ;
  assign new_n24175 = ~new_n23931 & ~new_n24174 ;
  assign new_n24176 = ~new_n23647 & ~new_n24175 ;
  assign new_n24177 = ~new_n24173 & ~new_n24176 ;
  assign new_n24178 = ~new_n2138 & ~new_n24177 ;
  assign new_n24179 = ~new_n24024 & ~new_n24178 ;
  assign new_n24180 = lo1313 & new_n24028 ;
  assign new_n24181 = new_n2138 & ~new_n24023 ;
  assign new_n24182 = ~new_n23668 & new_n23924 ;
  assign new_n24183 = ~new_n23928 & ~new_n24182 ;
  assign new_n24184 = new_n23658 & ~new_n24183 ;
  assign new_n24185 = new_n23668 & new_n23924 ;
  assign new_n24186 = ~new_n23925 & ~new_n24185 ;
  assign new_n24187 = ~new_n23658 & ~new_n24186 ;
  assign new_n24188 = ~new_n24184 & ~new_n24187 ;
  assign new_n24189 = ~new_n2138 & ~new_n24188 ;
  assign new_n24190 = ~new_n24181 & ~new_n24189 ;
  assign new_n24191 = lo1325 & new_n24028 ;
  assign new_n24192 = new_n2138 & ~new_n24037 ;
  assign new_n24193 = ~new_n23682 & new_n23918 ;
  assign new_n24194 = ~new_n23919 & ~new_n24193 ;
  assign new_n24195 = ~new_n23678 & ~new_n24194 ;
  assign new_n24196 = new_n23682 & new_n23918 ;
  assign new_n24197 = ~new_n23922 & ~new_n24196 ;
  assign new_n24198 = new_n23678 & ~new_n24197 ;
  assign new_n24199 = ~new_n24195 & ~new_n24198 ;
  assign new_n24200 = ~new_n2138 & ~new_n24199 ;
  assign new_n24201 = ~new_n24192 & ~new_n24200 ;
  assign new_n24202 = lo1338 & new_n24028 ;
  assign new_n24203 = new_n2138 & ~new_n24047 ;
  assign new_n24204 = pi446 & new_n23912 ;
  assign new_n24205 = ~new_n23913 & ~new_n24204 ;
  assign new_n24206 = ~new_n23692 & ~new_n24205 ;
  assign new_n24207 = ~pi446 & new_n23912 ;
  assign new_n24208 = ~new_n23916 & ~new_n24207 ;
  assign new_n24209 = new_n23692 & ~new_n24208 ;
  assign new_n24210 = ~new_n24206 & ~new_n24209 ;
  assign new_n24211 = ~new_n2138 & ~new_n24210 ;
  assign new_n24212 = ~new_n24203 & ~new_n24211 ;
  assign new_n24213 = lo1345 & new_n24028 ;
  assign new_n24214 = new_n2138 & ~new_n24057 ;
  assign new_n24215 = pi445 & new_n23906 ;
  assign new_n24216 = ~new_n23907 & ~new_n24215 ;
  assign new_n24217 = ~new_n23702 & ~new_n24216 ;
  assign new_n24218 = ~pi445 & new_n23906 ;
  assign new_n24219 = ~new_n23910 & ~new_n24218 ;
  assign new_n24220 = new_n23702 & ~new_n24219 ;
  assign new_n24221 = ~new_n24217 & ~new_n24220 ;
  assign new_n24222 = ~new_n2138 & ~new_n24221 ;
  assign new_n24223 = ~new_n24214 & ~new_n24222 ;
  assign new_n24224 = lo1398 & new_n24028 ;
  assign new_n24225 = new_n2138 & ~new_n24067 ;
  assign new_n24226 = pi444 & new_n23900 ;
  assign new_n24227 = ~new_n23901 & ~new_n24226 ;
  assign new_n24228 = ~new_n23712 & ~new_n24227 ;
  assign new_n24229 = ~pi444 & new_n23900 ;
  assign new_n24230 = ~new_n23904 & ~new_n24229 ;
  assign new_n24231 = new_n23712 & ~new_n24230 ;
  assign new_n24232 = ~new_n24228 & ~new_n24231 ;
  assign new_n24233 = ~new_n2138 & ~new_n24232 ;
  assign new_n24234 = ~new_n24225 & ~new_n24233 ;
  assign new_n24235 = lo1413 & new_n24028 ;
  assign new_n24236 = new_n2138 & ~new_n24077 ;
  assign new_n24237 = pi443 & new_n23894 ;
  assign new_n24238 = ~new_n23895 & ~new_n24237 ;
  assign new_n24239 = ~new_n23722 & ~new_n24238 ;
  assign new_n24240 = ~pi443 & new_n23894 ;
  assign new_n24241 = ~new_n23898 & ~new_n24240 ;
  assign new_n24242 = new_n23722 & ~new_n24241 ;
  assign new_n24243 = ~new_n24239 & ~new_n24242 ;
  assign new_n24244 = ~new_n2138 & ~new_n24243 ;
  assign new_n24245 = ~new_n24236 & ~new_n24244 ;
  assign new_n24246 = lo1387 & new_n24028 ;
  assign new_n24247 = new_n2138 & ~new_n24087 ;
  assign new_n24248 = pi442 & new_n23888 ;
  assign new_n24249 = ~new_n23889 & ~new_n24248 ;
  assign new_n24250 = ~new_n23732 & ~new_n24249 ;
  assign new_n24251 = ~pi442 & new_n23888 ;
  assign new_n24252 = ~new_n23892 & ~new_n24251 ;
  assign new_n24253 = new_n23732 & ~new_n24252 ;
  assign new_n24254 = ~new_n24250 & ~new_n24253 ;
  assign new_n24255 = ~new_n2138 & ~new_n24254 ;
  assign new_n24256 = ~new_n24247 & ~new_n24255 ;
  assign new_n24257 = lo1289 & new_n24028 ;
  assign new_n24258 = new_n2138 & ~new_n24097 ;
  assign new_n24259 = pi441 & new_n23882 ;
  assign new_n24260 = ~new_n23883 & ~new_n24259 ;
  assign new_n24261 = ~new_n23742 & ~new_n24260 ;
  assign new_n24262 = ~pi441 & new_n23882 ;
  assign new_n24263 = ~new_n23886 & ~new_n24262 ;
  assign new_n24264 = new_n23742 & ~new_n24263 ;
  assign new_n24265 = ~new_n24261 & ~new_n24264 ;
  assign new_n24266 = ~new_n2138 & ~new_n24265 ;
  assign new_n24267 = ~new_n24258 & ~new_n24266 ;
  assign new_n24268 = lo1311 & new_n24028 ;
  assign new_n24269 = new_n2138 & ~new_n24107 ;
  assign new_n24270 = pi440 & new_n23876 ;
  assign new_n24271 = ~new_n23877 & ~new_n24270 ;
  assign new_n24272 = ~new_n23752 & ~new_n24271 ;
  assign new_n24273 = ~pi440 & new_n23876 ;
  assign new_n24274 = ~new_n23880 & ~new_n24273 ;
  assign new_n24275 = new_n23752 & ~new_n24274 ;
  assign new_n24276 = ~new_n24272 & ~new_n24275 ;
  assign new_n24277 = ~new_n2138 & ~new_n24276 ;
  assign new_n24278 = ~new_n24269 & ~new_n24277 ;
  assign new_n24279 = lo1323 & new_n24028 ;
  assign new_n24280 = new_n2138 & ~new_n24117 ;
  assign new_n24281 = pi439 & new_n23870 ;
  assign new_n24282 = ~new_n23871 & ~new_n24281 ;
  assign new_n24283 = ~new_n23762 & ~new_n24282 ;
  assign new_n24284 = ~pi439 & new_n23870 ;
  assign new_n24285 = ~new_n23874 & ~new_n24284 ;
  assign new_n24286 = new_n23762 & ~new_n24285 ;
  assign new_n24287 = ~new_n24283 & ~new_n24286 ;
  assign new_n24288 = ~new_n2138 & ~new_n24287 ;
  assign new_n24289 = ~new_n24280 & ~new_n24288 ;
  assign new_n24290 = lo1335 & new_n24028 ;
  assign new_n24291 = new_n2138 & ~new_n24127 ;
  assign new_n24292 = pi438 & new_n23864 ;
  assign new_n24293 = ~new_n23865 & ~new_n24292 ;
  assign new_n24294 = ~new_n23772 & ~new_n24293 ;
  assign new_n24295 = ~pi438 & new_n23864 ;
  assign new_n24296 = ~new_n23868 & ~new_n24295 ;
  assign new_n24297 = new_n23772 & ~new_n24296 ;
  assign new_n24298 = ~new_n24294 & ~new_n24297 ;
  assign new_n24299 = ~new_n2138 & ~new_n24298 ;
  assign new_n24300 = ~new_n24291 & ~new_n24299 ;
  assign new_n24301 = lo1296 & new_n24028 ;
  assign new_n24302 = new_n2138 & ~new_n24137 ;
  assign new_n24303 = pi437 & new_n23858 ;
  assign new_n24304 = ~new_n23859 & ~new_n24303 ;
  assign new_n24305 = ~new_n23782 & ~new_n24304 ;
  assign new_n24306 = ~pi437 & new_n23858 ;
  assign new_n24307 = ~new_n23862 & ~new_n24306 ;
  assign new_n24308 = new_n23782 & ~new_n24307 ;
  assign new_n24309 = ~new_n24305 & ~new_n24308 ;
  assign new_n24310 = ~new_n2138 & ~new_n24309 ;
  assign new_n24311 = ~new_n24302 & ~new_n24310 ;
  assign new_n24312 = lo1374 & new_n24028 ;
  assign new_n24313 = new_n2138 & ~new_n24147 ;
  assign new_n24314 = pi436 & new_n23852 ;
  assign new_n24315 = ~new_n23853 & ~new_n24314 ;
  assign new_n24316 = ~new_n23792 & ~new_n24315 ;
  assign new_n24317 = ~pi436 & new_n23852 ;
  assign new_n24318 = ~new_n23856 & ~new_n24317 ;
  assign new_n24319 = new_n23792 & ~new_n24318 ;
  assign new_n24320 = ~new_n24316 & ~new_n24319 ;
  assign new_n24321 = ~new_n2138 & ~new_n24320 ;
  assign new_n24322 = ~new_n24313 & ~new_n24321 ;
  assign new_n24323 = lo1368 & new_n24028 ;
  assign new_n24324 = new_n2138 & ~new_n24157 ;
  assign new_n24325 = pi435 & new_n23846 ;
  assign new_n24326 = ~new_n23847 & ~new_n24325 ;
  assign new_n24327 = ~new_n23802 & ~new_n24326 ;
  assign new_n24328 = ~pi435 & new_n23846 ;
  assign new_n24329 = ~new_n23850 & ~new_n24328 ;
  assign new_n24330 = new_n23802 & ~new_n24329 ;
  assign new_n24331 = ~new_n24327 & ~new_n24330 ;
  assign new_n24332 = ~new_n2138 & ~new_n24331 ;
  assign new_n24333 = ~new_n24324 & ~new_n24332 ;
  assign new_n24334 = lo1383 & new_n24028 ;
  assign new_n24335 = new_n2138 & ~new_n24167 ;
  assign new_n24336 = pi434 & new_n23840 ;
  assign new_n24337 = ~new_n23841 & ~new_n24336 ;
  assign new_n24338 = ~new_n23812 & ~new_n24337 ;
  assign new_n24339 = ~pi434 & new_n23840 ;
  assign new_n24340 = ~new_n23844 & ~new_n24339 ;
  assign new_n24341 = new_n23812 & ~new_n24340 ;
  assign new_n24342 = ~new_n24338 & ~new_n24341 ;
  assign new_n24343 = ~new_n2138 & ~new_n24342 ;
  assign new_n24344 = ~new_n24335 & ~new_n24343 ;
  assign new_n24345 = lo1362 & new_n24028 ;
  assign new_n24346 = new_n2138 & ~new_n24177 ;
  assign new_n24347 = pi433 & new_n23834 ;
  assign new_n24348 = ~new_n23835 & ~new_n24347 ;
  assign new_n24349 = ~new_n23822 & ~new_n24348 ;
  assign new_n24350 = ~pi433 & new_n23834 ;
  assign new_n24351 = ~new_n23838 & ~new_n24350 ;
  assign new_n24352 = new_n23822 & ~new_n24351 ;
  assign new_n24353 = ~new_n24349 & ~new_n24352 ;
  assign new_n24354 = ~new_n2138 & ~new_n24353 ;
  assign new_n24355 = ~new_n24346 & ~new_n24354 ;
  assign new_n24356 = new_n2138 & ~new_n24188 ;
  assign new_n24357 = pi432 & ~new_n23242 ;
  assign new_n24358 = ~new_n23829 & ~new_n24357 ;
  assign new_n24359 = ~new_n23828 & ~new_n24358 ;
  assign new_n24360 = ~pi432 & ~new_n23242 ;
  assign new_n24361 = ~new_n23832 & ~new_n24360 ;
  assign new_n24362 = new_n23828 & ~new_n24361 ;
  assign new_n24363 = ~new_n24359 & ~new_n24362 ;
  assign new_n24364 = ~new_n2138 & ~new_n24363 ;
  assign new_n24365 = ~new_n24356 & ~new_n24364 ;
  assign new_n24366 = new_n2138 & ~new_n24199 ;
  assign new_n24367 = pi431 & ~new_n2138 ;
  assign new_n24368 = ~new_n24366 & ~new_n24367 ;
  assign new_n24369 = new_n2138 & ~new_n24210 ;
  assign new_n24370 = pi430 & ~new_n2138 ;
  assign new_n24371 = ~new_n24369 & ~new_n24370 ;
  assign new_n24372 = new_n2138 & ~new_n24221 ;
  assign new_n24373 = pi429 & ~new_n2138 ;
  assign new_n24374 = ~new_n24372 & ~new_n24373 ;
  assign new_n24375 = new_n2138 & ~new_n24232 ;
  assign new_n24376 = pi428 & ~new_n2138 ;
  assign new_n24377 = ~new_n24375 & ~new_n24376 ;
  assign new_n24378 = new_n2138 & ~new_n24243 ;
  assign new_n24379 = pi427 & ~new_n2138 ;
  assign new_n24380 = ~new_n24378 & ~new_n24379 ;
  assign new_n24381 = new_n2138 & ~new_n24254 ;
  assign new_n24382 = pi426 & ~new_n2138 ;
  assign new_n24383 = ~new_n24381 & ~new_n24382 ;
  assign new_n24384 = new_n2138 & ~new_n24265 ;
  assign new_n24385 = pi425 & ~new_n2138 ;
  assign new_n24386 = ~new_n24384 & ~new_n24385 ;
  assign new_n24387 = new_n2138 & ~new_n24276 ;
  assign new_n24388 = pi424 & ~new_n2138 ;
  assign new_n24389 = ~new_n24387 & ~new_n24388 ;
  assign new_n24390 = new_n2138 & ~new_n24287 ;
  assign new_n24391 = pi423 & ~new_n2138 ;
  assign new_n24392 = ~new_n24390 & ~new_n24391 ;
  assign new_n24393 = new_n2138 & ~new_n24298 ;
  assign new_n24394 = pi422 & ~new_n2138 ;
  assign new_n24395 = ~new_n24393 & ~new_n24394 ;
  assign new_n24396 = new_n2138 & ~new_n24309 ;
  assign new_n24397 = pi421 & ~new_n2138 ;
  assign new_n24398 = ~new_n24396 & ~new_n24397 ;
  assign new_n24399 = new_n2138 & ~new_n24320 ;
  assign new_n24400 = pi420 & ~new_n2138 ;
  assign new_n24401 = ~new_n24399 & ~new_n24400 ;
  assign new_n24402 = new_n2138 & ~new_n24331 ;
  assign new_n24403 = pi419 & ~new_n2138 ;
  assign new_n24404 = ~new_n24402 & ~new_n24403 ;
  assign new_n24405 = new_n2138 & ~new_n24342 ;
  assign new_n24406 = pi418 & ~new_n2138 ;
  assign new_n24407 = ~new_n24405 & ~new_n24406 ;
  assign new_n24408 = new_n2138 & ~new_n24353 ;
  assign new_n24409 = pi417 & ~new_n2138 ;
  assign new_n24410 = ~new_n24408 & ~new_n24409 ;
  assign new_n24411 = new_n2138 & ~new_n24363 ;
  assign new_n24412 = pi431 & new_n2138 ;
  assign new_n24413 = pi430 & new_n2138 ;
  assign new_n24414 = pi429 & new_n2138 ;
  assign new_n24415 = pi428 & new_n2138 ;
  assign new_n24416 = pi427 & new_n2138 ;
  assign new_n24417 = pi426 & new_n2138 ;
  assign new_n24418 = ~lo1287 & ~new_n23235 ;
  assign new_n24419 = new_n23179 & ~new_n24418 ;
  assign new_n24420 = ~new_n23179 & new_n23231 ;
  assign new_n24421 = ~new_n24419 & ~new_n24420 ;
  assign new_n24422 = ~lo1386 & ~new_n24421 ;
  assign new_n24423 = ~lo1386 & ~new_n24422 ;
  assign new_n24424 = new_n24417 & ~new_n24423 ;
  assign new_n24425 = lo1386 & ~new_n24421 ;
  assign new_n24426 = ~new_n24417 & new_n24425 ;
  assign new_n24427 = ~new_n24424 & ~new_n24426 ;
  assign new_n24428 = ~lo1411 & ~new_n24427 ;
  assign new_n24429 = ~lo1411 & ~new_n24428 ;
  assign new_n24430 = new_n24416 & ~new_n24429 ;
  assign new_n24431 = lo1411 & ~new_n24427 ;
  assign new_n24432 = ~new_n24416 & new_n24431 ;
  assign new_n24433 = ~new_n24430 & ~new_n24432 ;
  assign new_n24434 = ~lo1396 & ~new_n24433 ;
  assign new_n24435 = ~lo1396 & ~new_n24434 ;
  assign new_n24436 = new_n24415 & ~new_n24435 ;
  assign new_n24437 = lo1396 & ~new_n24433 ;
  assign new_n24438 = ~new_n24415 & new_n24437 ;
  assign new_n24439 = ~new_n24436 & ~new_n24438 ;
  assign new_n24440 = ~lo1347 & ~new_n24439 ;
  assign new_n24441 = ~lo1347 & ~new_n24440 ;
  assign new_n24442 = new_n24414 & ~new_n24441 ;
  assign new_n24443 = lo1347 & ~new_n24439 ;
  assign new_n24444 = ~new_n24414 & new_n24443 ;
  assign new_n24445 = ~new_n24442 & ~new_n24444 ;
  assign new_n24446 = ~lo1340 & ~new_n24445 ;
  assign new_n24447 = ~lo1340 & ~new_n24446 ;
  assign new_n24448 = new_n24413 & ~new_n24447 ;
  assign new_n24449 = lo1340 & ~new_n24445 ;
  assign new_n24450 = ~new_n24413 & new_n24449 ;
  assign new_n24451 = ~new_n24448 & ~new_n24450 ;
  assign new_n24452 = ~lo1327 & ~new_n24451 ;
  assign new_n24453 = ~lo1327 & ~new_n24452 ;
  assign new_n24454 = new_n24412 & ~new_n24453 ;
  assign new_n24455 = lo1327 & ~new_n24451 ;
  assign new_n24456 = ~new_n24412 & new_n24455 ;
  assign new_n24457 = ~new_n24454 & ~new_n24456 ;
  assign new_n24458 = ~lo1316 & ~new_n24457 ;
  assign new_n24459 = ~lo1316 & ~new_n24458 ;
  assign new_n24460 = new_n24411 & ~new_n24459 ;
  assign new_n24461 = lo1316 & ~new_n24457 ;
  assign new_n24462 = ~new_n24411 & new_n24461 ;
  assign new_n24463 = ~new_n24460 & ~new_n24462 ;
  assign new_n24464 = ~lo1366 & ~new_n24463 ;
  assign new_n24465 = ~lo1366 & ~new_n24464 ;
  assign new_n24466 = ~new_n24410 & ~new_n24465 ;
  assign new_n24467 = lo1366 & ~new_n24463 ;
  assign new_n24468 = new_n24410 & new_n24467 ;
  assign new_n24469 = ~new_n24466 & ~new_n24468 ;
  assign new_n24470 = ~lo1391 & ~new_n24469 ;
  assign new_n24471 = ~lo1391 & ~new_n24470 ;
  assign new_n24472 = ~new_n24407 & ~new_n24471 ;
  assign new_n24473 = lo1391 & ~new_n24469 ;
  assign new_n24474 = new_n24407 & new_n24473 ;
  assign new_n24475 = ~new_n24472 & ~new_n24474 ;
  assign new_n24476 = ~lo1373 & ~new_n24475 ;
  assign new_n24477 = ~lo1373 & ~new_n24476 ;
  assign new_n24478 = ~new_n24404 & ~new_n24477 ;
  assign new_n24479 = lo1373 & ~new_n24475 ;
  assign new_n24480 = new_n24404 & new_n24479 ;
  assign new_n24481 = ~new_n24478 & ~new_n24480 ;
  assign new_n24482 = ~lo1379 & ~new_n24481 ;
  assign new_n24483 = ~lo1379 & ~new_n24482 ;
  assign new_n24484 = ~new_n24401 & ~new_n24483 ;
  assign new_n24485 = lo1379 & ~new_n24481 ;
  assign new_n24486 = new_n24401 & new_n24485 ;
  assign new_n24487 = ~new_n24484 & ~new_n24486 ;
  assign new_n24488 = ~lo1302 & ~new_n24487 ;
  assign new_n24489 = ~lo1302 & ~new_n24488 ;
  assign new_n24490 = ~new_n24398 & ~new_n24489 ;
  assign new_n24491 = lo1302 & ~new_n24487 ;
  assign new_n24492 = new_n24398 & new_n24491 ;
  assign new_n24493 = ~new_n24490 & ~new_n24492 ;
  assign new_n24494 = ~lo1343 & ~new_n24493 ;
  assign new_n24495 = ~lo1343 & ~new_n24494 ;
  assign new_n24496 = ~new_n24395 & ~new_n24495 ;
  assign new_n24497 = lo1343 & ~new_n24493 ;
  assign new_n24498 = new_n24395 & new_n24497 ;
  assign new_n24499 = ~new_n24496 & ~new_n24498 ;
  assign new_n24500 = ~lo1358 & ~new_n24499 ;
  assign new_n24501 = ~lo1358 & ~new_n24500 ;
  assign new_n24502 = ~new_n24392 & ~new_n24501 ;
  assign new_n24503 = lo1358 & ~new_n24499 ;
  assign new_n24504 = new_n24392 & new_n24503 ;
  assign new_n24505 = ~new_n24502 & ~new_n24504 ;
  assign new_n24506 = ~lo1395 & ~new_n24505 ;
  assign new_n24507 = ~lo1395 & ~new_n24506 ;
  assign new_n24508 = ~new_n24389 & ~new_n24507 ;
  assign new_n24509 = lo1395 & ~new_n24505 ;
  assign new_n24510 = new_n24389 & new_n24509 ;
  assign new_n24511 = ~new_n24508 & ~new_n24510 ;
  assign new_n24512 = ~lo1419 & ~new_n24511 ;
  assign new_n24513 = ~lo1419 & ~new_n24512 ;
  assign new_n24514 = ~new_n24386 & ~new_n24513 ;
  assign new_n24515 = lo1419 & ~new_n24511 ;
  assign new_n24516 = new_n24386 & new_n24515 ;
  assign new_n24517 = ~new_n24514 & ~new_n24516 ;
  assign new_n24518 = ~lo1404 & ~new_n24517 ;
  assign new_n24519 = ~lo1404 & ~new_n24518 ;
  assign new_n24520 = ~new_n24383 & ~new_n24519 ;
  assign new_n24521 = lo1404 & ~new_n24517 ;
  assign new_n24522 = new_n24383 & new_n24521 ;
  assign new_n24523 = ~new_n24520 & ~new_n24522 ;
  assign new_n24524 = ~lo1416 & ~new_n24523 ;
  assign new_n24525 = ~lo1416 & ~new_n24524 ;
  assign new_n24526 = ~new_n24380 & ~new_n24525 ;
  assign new_n24527 = lo1416 & ~new_n24523 ;
  assign new_n24528 = new_n24380 & new_n24527 ;
  assign new_n24529 = ~new_n24526 & ~new_n24528 ;
  assign new_n24530 = ~lo1401 & ~new_n24529 ;
  assign new_n24531 = ~lo1401 & ~new_n24530 ;
  assign new_n24532 = ~new_n24377 & ~new_n24531 ;
  assign new_n24533 = lo1401 & ~new_n24529 ;
  assign new_n24534 = new_n24377 & new_n24533 ;
  assign new_n24535 = ~new_n24532 & ~new_n24534 ;
  assign new_n24536 = ~lo1355 & ~new_n24535 ;
  assign new_n24537 = ~lo1355 & ~new_n24536 ;
  assign new_n24538 = ~new_n24374 & ~new_n24537 ;
  assign new_n24539 = lo1355 & ~new_n24535 ;
  assign new_n24540 = new_n24374 & new_n24539 ;
  assign new_n24541 = ~new_n24538 & ~new_n24540 ;
  assign new_n24542 = ~lo1407 & ~new_n24541 ;
  assign new_n24543 = ~lo1407 & ~new_n24542 ;
  assign new_n24544 = ~new_n24371 & ~new_n24543 ;
  assign new_n24545 = lo1407 & ~new_n24541 ;
  assign new_n24546 = new_n24371 & new_n24545 ;
  assign new_n24547 = ~new_n24544 & ~new_n24546 ;
  assign new_n24548 = ~lo1332 & ~new_n24547 ;
  assign new_n24549 = ~lo1332 & ~new_n24548 ;
  assign new_n24550 = ~new_n24368 & ~new_n24549 ;
  assign new_n24551 = lo1332 & ~new_n24547 ;
  assign new_n24552 = new_n24368 & new_n24551 ;
  assign new_n24553 = ~new_n24550 & ~new_n24552 ;
  assign new_n24554 = ~lo1410 & ~new_n24553 ;
  assign new_n24555 = ~lo1410 & ~new_n24554 ;
  assign new_n24556 = ~new_n24365 & ~new_n24555 ;
  assign new_n24557 = lo1410 & ~new_n24553 ;
  assign new_n24558 = new_n24365 & new_n24557 ;
  assign new_n24559 = ~new_n24556 & ~new_n24558 ;
  assign new_n24560 = new_n24355 & ~new_n24559 ;
  assign new_n24561 = new_n24355 & ~new_n24560 ;
  assign new_n24562 = new_n24345 & ~new_n24561 ;
  assign new_n24563 = ~new_n24355 & ~new_n24559 ;
  assign new_n24564 = ~new_n24345 & new_n24563 ;
  assign new_n24565 = ~new_n24562 & ~new_n24564 ;
  assign new_n24566 = new_n24344 & ~new_n24565 ;
  assign new_n24567 = new_n24344 & ~new_n24566 ;
  assign new_n24568 = new_n24334 & ~new_n24567 ;
  assign new_n24569 = ~new_n24344 & ~new_n24565 ;
  assign new_n24570 = ~new_n24334 & new_n24569 ;
  assign new_n24571 = ~new_n24568 & ~new_n24570 ;
  assign new_n24572 = new_n24333 & ~new_n24571 ;
  assign new_n24573 = new_n24333 & ~new_n24572 ;
  assign new_n24574 = new_n24323 & ~new_n24573 ;
  assign new_n24575 = ~new_n24333 & ~new_n24571 ;
  assign new_n24576 = ~new_n24323 & new_n24575 ;
  assign new_n24577 = ~new_n24574 & ~new_n24576 ;
  assign new_n24578 = new_n24322 & ~new_n24577 ;
  assign new_n24579 = new_n24322 & ~new_n24578 ;
  assign new_n24580 = new_n24312 & ~new_n24579 ;
  assign new_n24581 = ~new_n24322 & ~new_n24577 ;
  assign new_n24582 = ~new_n24312 & new_n24581 ;
  assign new_n24583 = ~new_n24580 & ~new_n24582 ;
  assign new_n24584 = new_n24311 & ~new_n24583 ;
  assign new_n24585 = new_n24311 & ~new_n24584 ;
  assign new_n24586 = new_n24301 & ~new_n24585 ;
  assign new_n24587 = ~new_n24311 & ~new_n24583 ;
  assign new_n24588 = ~new_n24301 & new_n24587 ;
  assign new_n24589 = ~new_n24586 & ~new_n24588 ;
  assign new_n24590 = new_n24300 & ~new_n24589 ;
  assign new_n24591 = new_n24300 & ~new_n24590 ;
  assign new_n24592 = new_n24290 & ~new_n24591 ;
  assign new_n24593 = ~new_n24300 & ~new_n24589 ;
  assign new_n24594 = ~new_n24290 & new_n24593 ;
  assign new_n24595 = ~new_n24592 & ~new_n24594 ;
  assign new_n24596 = new_n24289 & ~new_n24595 ;
  assign new_n24597 = new_n24289 & ~new_n24596 ;
  assign new_n24598 = new_n24279 & ~new_n24597 ;
  assign new_n24599 = ~new_n24289 & ~new_n24595 ;
  assign new_n24600 = ~new_n24279 & new_n24599 ;
  assign new_n24601 = ~new_n24598 & ~new_n24600 ;
  assign new_n24602 = new_n24278 & ~new_n24601 ;
  assign new_n24603 = new_n24278 & ~new_n24602 ;
  assign new_n24604 = new_n24268 & ~new_n24603 ;
  assign new_n24605 = ~new_n24278 & ~new_n24601 ;
  assign new_n24606 = ~new_n24268 & new_n24605 ;
  assign new_n24607 = ~new_n24604 & ~new_n24606 ;
  assign new_n24608 = new_n24267 & ~new_n24607 ;
  assign new_n24609 = new_n24267 & ~new_n24608 ;
  assign new_n24610 = new_n24257 & ~new_n24609 ;
  assign new_n24611 = ~new_n24267 & ~new_n24607 ;
  assign new_n24612 = ~new_n24257 & new_n24611 ;
  assign new_n24613 = ~new_n24610 & ~new_n24612 ;
  assign new_n24614 = new_n24256 & ~new_n24613 ;
  assign new_n24615 = new_n24256 & ~new_n24614 ;
  assign new_n24616 = new_n24246 & ~new_n24615 ;
  assign new_n24617 = ~new_n24256 & ~new_n24613 ;
  assign new_n24618 = ~new_n24246 & new_n24617 ;
  assign new_n24619 = ~new_n24616 & ~new_n24618 ;
  assign new_n24620 = new_n24245 & ~new_n24619 ;
  assign new_n24621 = new_n24245 & ~new_n24620 ;
  assign new_n24622 = new_n24235 & ~new_n24621 ;
  assign new_n24623 = ~new_n24245 & ~new_n24619 ;
  assign new_n24624 = ~new_n24235 & new_n24623 ;
  assign new_n24625 = ~new_n24622 & ~new_n24624 ;
  assign new_n24626 = new_n24234 & ~new_n24625 ;
  assign new_n24627 = new_n24234 & ~new_n24626 ;
  assign new_n24628 = new_n24224 & ~new_n24627 ;
  assign new_n24629 = ~new_n24234 & ~new_n24625 ;
  assign new_n24630 = ~new_n24224 & new_n24629 ;
  assign new_n24631 = ~new_n24628 & ~new_n24630 ;
  assign new_n24632 = new_n24223 & ~new_n24631 ;
  assign new_n24633 = new_n24223 & ~new_n24632 ;
  assign new_n24634 = new_n24213 & ~new_n24633 ;
  assign new_n24635 = ~new_n24223 & ~new_n24631 ;
  assign new_n24636 = ~new_n24213 & new_n24635 ;
  assign new_n24637 = ~new_n24634 & ~new_n24636 ;
  assign new_n24638 = new_n24212 & ~new_n24637 ;
  assign new_n24639 = new_n24212 & ~new_n24638 ;
  assign new_n24640 = new_n24202 & ~new_n24639 ;
  assign new_n24641 = ~new_n24212 & ~new_n24637 ;
  assign new_n24642 = ~new_n24202 & new_n24641 ;
  assign new_n24643 = ~new_n24640 & ~new_n24642 ;
  assign new_n24644 = new_n24201 & ~new_n24643 ;
  assign new_n24645 = new_n24201 & ~new_n24644 ;
  assign new_n24646 = new_n24191 & ~new_n24645 ;
  assign new_n24647 = ~new_n24201 & ~new_n24643 ;
  assign new_n24648 = ~new_n24191 & new_n24647 ;
  assign new_n24649 = ~new_n24646 & ~new_n24648 ;
  assign new_n24650 = new_n24190 & ~new_n24649 ;
  assign new_n24651 = new_n24190 & ~new_n24650 ;
  assign new_n24652 = new_n24180 & ~new_n24651 ;
  assign new_n24653 = ~new_n24190 & ~new_n24649 ;
  assign new_n24654 = ~new_n24180 & new_n24653 ;
  assign new_n24655 = ~new_n24652 & ~new_n24654 ;
  assign new_n24656 = new_n24179 & ~new_n24655 ;
  assign new_n24657 = new_n24179 & ~new_n24656 ;
  assign new_n24658 = new_n24170 & ~new_n24657 ;
  assign new_n24659 = ~new_n24179 & ~new_n24655 ;
  assign new_n24660 = ~new_n24170 & new_n24659 ;
  assign new_n24661 = ~new_n24658 & ~new_n24660 ;
  assign new_n24662 = new_n24169 & ~new_n24661 ;
  assign new_n24663 = new_n24169 & ~new_n24662 ;
  assign new_n24664 = new_n24160 & ~new_n24663 ;
  assign new_n24665 = ~new_n24169 & ~new_n24661 ;
  assign new_n24666 = ~new_n24160 & new_n24665 ;
  assign new_n24667 = ~new_n24664 & ~new_n24666 ;
  assign new_n24668 = new_n24159 & ~new_n24667 ;
  assign new_n24669 = new_n24159 & ~new_n24668 ;
  assign new_n24670 = new_n24150 & ~new_n24669 ;
  assign new_n24671 = ~new_n24159 & ~new_n24667 ;
  assign new_n24672 = ~new_n24150 & new_n24671 ;
  assign new_n24673 = ~new_n24670 & ~new_n24672 ;
  assign new_n24674 = new_n24149 & ~new_n24673 ;
  assign new_n24675 = new_n24149 & ~new_n24674 ;
  assign new_n24676 = new_n24140 & ~new_n24675 ;
  assign new_n24677 = ~new_n24149 & ~new_n24673 ;
  assign new_n24678 = ~new_n24140 & new_n24677 ;
  assign new_n24679 = ~new_n24676 & ~new_n24678 ;
  assign new_n24680 = new_n24139 & ~new_n24679 ;
  assign new_n24681 = new_n24139 & ~new_n24680 ;
  assign new_n24682 = new_n24130 & ~new_n24681 ;
  assign new_n24683 = ~new_n24139 & ~new_n24679 ;
  assign new_n24684 = ~new_n24130 & new_n24683 ;
  assign new_n24685 = ~new_n24682 & ~new_n24684 ;
  assign new_n24686 = new_n24129 & ~new_n24685 ;
  assign new_n24687 = new_n24129 & ~new_n24686 ;
  assign new_n24688 = new_n24120 & ~new_n24687 ;
  assign new_n24689 = ~new_n24129 & ~new_n24685 ;
  assign new_n24690 = ~new_n24120 & new_n24689 ;
  assign new_n24691 = ~new_n24688 & ~new_n24690 ;
  assign new_n24692 = new_n24119 & ~new_n24691 ;
  assign new_n24693 = new_n24119 & ~new_n24692 ;
  assign new_n24694 = new_n24110 & ~new_n24693 ;
  assign new_n24695 = ~new_n24119 & ~new_n24691 ;
  assign new_n24696 = ~new_n24110 & new_n24695 ;
  assign new_n24697 = ~new_n24694 & ~new_n24696 ;
  assign new_n24698 = new_n24109 & ~new_n24697 ;
  assign new_n24699 = new_n24109 & ~new_n24698 ;
  assign new_n24700 = new_n24100 & ~new_n24699 ;
  assign new_n24701 = ~new_n24109 & ~new_n24697 ;
  assign new_n24702 = ~new_n24100 & new_n24701 ;
  assign new_n24703 = ~new_n24700 & ~new_n24702 ;
  assign new_n24704 = new_n24099 & ~new_n24703 ;
  assign new_n24705 = new_n24099 & ~new_n24704 ;
  assign new_n24706 = new_n24090 & ~new_n24705 ;
  assign new_n24707 = ~new_n24099 & ~new_n24703 ;
  assign new_n24708 = ~new_n24090 & new_n24707 ;
  assign new_n24709 = ~new_n24706 & ~new_n24708 ;
  assign new_n24710 = new_n24089 & ~new_n24709 ;
  assign new_n24711 = new_n24089 & ~new_n24710 ;
  assign new_n24712 = new_n24080 & ~new_n24711 ;
  assign new_n24713 = ~new_n24089 & ~new_n24709 ;
  assign new_n24714 = ~new_n24080 & new_n24713 ;
  assign new_n24715 = ~new_n24712 & ~new_n24714 ;
  assign new_n24716 = new_n24079 & ~new_n24715 ;
  assign new_n24717 = new_n24079 & ~new_n24716 ;
  assign new_n24718 = new_n24070 & ~new_n24717 ;
  assign new_n24719 = ~new_n24079 & ~new_n24715 ;
  assign new_n24720 = ~new_n24070 & new_n24719 ;
  assign new_n24721 = ~new_n24718 & ~new_n24720 ;
  assign new_n24722 = new_n24069 & ~new_n24721 ;
  assign new_n24723 = new_n24069 & ~new_n24722 ;
  assign new_n24724 = new_n24060 & ~new_n24723 ;
  assign new_n24725 = ~new_n24069 & ~new_n24721 ;
  assign new_n24726 = ~new_n24060 & new_n24725 ;
  assign new_n24727 = ~new_n24724 & ~new_n24726 ;
  assign new_n24728 = new_n24059 & ~new_n24727 ;
  assign new_n24729 = new_n24059 & ~new_n24728 ;
  assign new_n24730 = new_n24050 & ~new_n24729 ;
  assign new_n24731 = ~new_n24059 & ~new_n24727 ;
  assign new_n24732 = ~new_n24050 & new_n24731 ;
  assign new_n24733 = ~new_n24730 & ~new_n24732 ;
  assign new_n24734 = new_n24049 & ~new_n24733 ;
  assign new_n24735 = new_n24049 & ~new_n24734 ;
  assign new_n24736 = new_n24040 & ~new_n24735 ;
  assign new_n24737 = ~new_n24049 & ~new_n24733 ;
  assign new_n24738 = ~new_n24040 & new_n24737 ;
  assign new_n24739 = ~new_n24736 & ~new_n24738 ;
  assign new_n24740 = new_n24039 & ~new_n24739 ;
  assign new_n24741 = new_n24039 & ~new_n24740 ;
  assign new_n24742 = new_n24030 & ~new_n24741 ;
  assign new_n24743 = ~new_n24039 & ~new_n24739 ;
  assign new_n24744 = ~new_n24030 & new_n24743 ;
  assign new_n24745 = ~new_n24742 & ~new_n24744 ;
  assign new_n24746 = new_n24026 & ~new_n24745 ;
  assign new_n24747 = ~new_n24026 & new_n24745 ;
  assign new_n24748 = ~new_n24746 & ~new_n24747 ;
  assign new_n24749 = new_n24029 & ~new_n24748 ;
  assign new_n24750 = ~new_n24026 & ~new_n24745 ;
  assign new_n24751 = new_n24026 & new_n24745 ;
  assign new_n24752 = ~new_n24750 & ~new_n24751 ;
  assign new_n24753 = ~new_n24029 & ~new_n24752 ;
  assign new_n24754 = ~new_n24749 & ~new_n24753 ;
  assign new_n24755 = ~lo1408 & new_n24754 ;
  assign new_n24756 = new_n24026 & ~new_n24755 ;
  assign new_n24757 = ~new_n24027 & ~new_n24756 ;
  assign new_n24758 = ~new_n21027 & ~new_n24757 ;
  assign new_n24759 = ~lo0941 & ~new_n24758 ;
  assign new_n24760 = ~new_n24026 & new_n24759 ;
  assign new_n24761 = lo0941 & ~new_n24365 ;
  assign new_n24762 = ~lo1408 & new_n24026 ;
  assign new_n24763 = new_n24754 & ~new_n24762 ;
  assign new_n24764 = ~lo0941 & ~new_n21027 ;
  assign new_n24765 = new_n24763 & new_n24764 ;
  assign new_n24766 = ~new_n24761 & ~new_n24765 ;
  assign new_n24767 = ~new_n23174 & new_n24766 ;
  assign new_n24768 = ~new_n24760 & new_n24767 ;
  assign new_n24769 = ~lo1410 & new_n24553 ;
  assign new_n24770 = ~new_n24557 & ~new_n24769 ;
  assign new_n24771 = ~new_n24365 & ~new_n24770 ;
  assign new_n24772 = lo1410 & new_n24553 ;
  assign new_n24773 = ~new_n24554 & ~new_n24772 ;
  assign new_n24774 = new_n24365 & ~new_n24773 ;
  assign new_n24775 = ~new_n24771 & ~new_n24774 ;
  assign new_n24776 = lo1410 & new_n24775 ;
  assign new_n24777 = ~new_n24766 & ~new_n24776 ;
  assign new_n24778 = lo1410 & new_n24766 ;
  assign new_n24779 = ~lo1410 & new_n24775 ;
  assign new_n24780 = ~new_n24778 & ~new_n24779 ;
  assign new_n24781 = ~new_n24777 & new_n24780 ;
  assign new_n24782 = lo0941 & ~new_n24781 ;
  assign new_n24783 = new_n24039 & new_n24739 ;
  assign new_n24784 = ~new_n24743 & ~new_n24783 ;
  assign new_n24785 = new_n24030 & ~new_n24784 ;
  assign new_n24786 = ~new_n24039 & new_n24739 ;
  assign new_n24787 = ~new_n24740 & ~new_n24786 ;
  assign new_n24788 = ~new_n24030 & ~new_n24787 ;
  assign new_n24789 = ~new_n24785 & ~new_n24788 ;
  assign new_n24790 = new_n24049 & new_n24733 ;
  assign new_n24791 = ~new_n24737 & ~new_n24790 ;
  assign new_n24792 = new_n24040 & ~new_n24791 ;
  assign new_n24793 = ~new_n24049 & new_n24733 ;
  assign new_n24794 = ~new_n24734 & ~new_n24793 ;
  assign new_n24795 = ~new_n24040 & ~new_n24794 ;
  assign new_n24796 = ~new_n24792 & ~new_n24795 ;
  assign new_n24797 = new_n24059 & new_n24727 ;
  assign new_n24798 = ~new_n24731 & ~new_n24797 ;
  assign new_n24799 = new_n24050 & ~new_n24798 ;
  assign new_n24800 = ~new_n24059 & new_n24727 ;
  assign new_n24801 = ~new_n24728 & ~new_n24800 ;
  assign new_n24802 = ~new_n24050 & ~new_n24801 ;
  assign new_n24803 = ~new_n24799 & ~new_n24802 ;
  assign new_n24804 = new_n24069 & new_n24721 ;
  assign new_n24805 = ~new_n24725 & ~new_n24804 ;
  assign new_n24806 = new_n24060 & ~new_n24805 ;
  assign new_n24807 = ~new_n24069 & new_n24721 ;
  assign new_n24808 = ~new_n24722 & ~new_n24807 ;
  assign new_n24809 = ~new_n24060 & ~new_n24808 ;
  assign new_n24810 = ~new_n24806 & ~new_n24809 ;
  assign new_n24811 = new_n24079 & new_n24715 ;
  assign new_n24812 = ~new_n24719 & ~new_n24811 ;
  assign new_n24813 = new_n24070 & ~new_n24812 ;
  assign new_n24814 = ~new_n24079 & new_n24715 ;
  assign new_n24815 = ~new_n24716 & ~new_n24814 ;
  assign new_n24816 = ~new_n24070 & ~new_n24815 ;
  assign new_n24817 = ~new_n24813 & ~new_n24816 ;
  assign new_n24818 = new_n24089 & new_n24709 ;
  assign new_n24819 = ~new_n24713 & ~new_n24818 ;
  assign new_n24820 = new_n24080 & ~new_n24819 ;
  assign new_n24821 = ~new_n24089 & new_n24709 ;
  assign new_n24822 = ~new_n24710 & ~new_n24821 ;
  assign new_n24823 = ~new_n24080 & ~new_n24822 ;
  assign new_n24824 = ~new_n24820 & ~new_n24823 ;
  assign new_n24825 = new_n24099 & new_n24703 ;
  assign new_n24826 = ~new_n24707 & ~new_n24825 ;
  assign new_n24827 = new_n24090 & ~new_n24826 ;
  assign new_n24828 = ~new_n24099 & new_n24703 ;
  assign new_n24829 = ~new_n24704 & ~new_n24828 ;
  assign new_n24830 = ~new_n24090 & ~new_n24829 ;
  assign new_n24831 = ~new_n24827 & ~new_n24830 ;
  assign new_n24832 = new_n24109 & new_n24697 ;
  assign new_n24833 = ~new_n24701 & ~new_n24832 ;
  assign new_n24834 = new_n24100 & ~new_n24833 ;
  assign new_n24835 = ~new_n24109 & new_n24697 ;
  assign new_n24836 = ~new_n24698 & ~new_n24835 ;
  assign new_n24837 = ~new_n24100 & ~new_n24836 ;
  assign new_n24838 = ~new_n24834 & ~new_n24837 ;
  assign new_n24839 = new_n24119 & new_n24691 ;
  assign new_n24840 = ~new_n24695 & ~new_n24839 ;
  assign new_n24841 = new_n24110 & ~new_n24840 ;
  assign new_n24842 = ~new_n24119 & new_n24691 ;
  assign new_n24843 = ~new_n24692 & ~new_n24842 ;
  assign new_n24844 = ~new_n24110 & ~new_n24843 ;
  assign new_n24845 = ~new_n24841 & ~new_n24844 ;
  assign new_n24846 = new_n24129 & new_n24685 ;
  assign new_n24847 = ~new_n24689 & ~new_n24846 ;
  assign new_n24848 = new_n24120 & ~new_n24847 ;
  assign new_n24849 = ~new_n24129 & new_n24685 ;
  assign new_n24850 = ~new_n24686 & ~new_n24849 ;
  assign new_n24851 = ~new_n24120 & ~new_n24850 ;
  assign new_n24852 = ~new_n24848 & ~new_n24851 ;
  assign new_n24853 = new_n24139 & new_n24679 ;
  assign new_n24854 = ~new_n24683 & ~new_n24853 ;
  assign new_n24855 = new_n24130 & ~new_n24854 ;
  assign new_n24856 = ~new_n24139 & new_n24679 ;
  assign new_n24857 = ~new_n24680 & ~new_n24856 ;
  assign new_n24858 = ~new_n24130 & ~new_n24857 ;
  assign new_n24859 = ~new_n24855 & ~new_n24858 ;
  assign new_n24860 = new_n24149 & new_n24673 ;
  assign new_n24861 = ~new_n24677 & ~new_n24860 ;
  assign new_n24862 = new_n24140 & ~new_n24861 ;
  assign new_n24863 = ~new_n24149 & new_n24673 ;
  assign new_n24864 = ~new_n24674 & ~new_n24863 ;
  assign new_n24865 = ~new_n24140 & ~new_n24864 ;
  assign new_n24866 = ~new_n24862 & ~new_n24865 ;
  assign new_n24867 = new_n24159 & new_n24667 ;
  assign new_n24868 = ~new_n24671 & ~new_n24867 ;
  assign new_n24869 = new_n24150 & ~new_n24868 ;
  assign new_n24870 = ~new_n24159 & new_n24667 ;
  assign new_n24871 = ~new_n24668 & ~new_n24870 ;
  assign new_n24872 = ~new_n24150 & ~new_n24871 ;
  assign new_n24873 = ~new_n24869 & ~new_n24872 ;
  assign new_n24874 = new_n24169 & new_n24661 ;
  assign new_n24875 = ~new_n24665 & ~new_n24874 ;
  assign new_n24876 = new_n24160 & ~new_n24875 ;
  assign new_n24877 = ~new_n24169 & new_n24661 ;
  assign new_n24878 = ~new_n24662 & ~new_n24877 ;
  assign new_n24879 = ~new_n24160 & ~new_n24878 ;
  assign new_n24880 = ~new_n24876 & ~new_n24879 ;
  assign new_n24881 = new_n24190 & new_n24649 ;
  assign new_n24882 = ~new_n24653 & ~new_n24881 ;
  assign new_n24883 = new_n24180 & ~new_n24882 ;
  assign new_n24884 = ~new_n24190 & new_n24649 ;
  assign new_n24885 = ~new_n24650 & ~new_n24884 ;
  assign new_n24886 = ~new_n24180 & ~new_n24885 ;
  assign new_n24887 = ~new_n24883 & ~new_n24886 ;
  assign new_n24888 = new_n24179 & new_n24655 ;
  assign new_n24889 = ~new_n24659 & ~new_n24888 ;
  assign new_n24890 = new_n24170 & ~new_n24889 ;
  assign new_n24891 = ~new_n24179 & new_n24655 ;
  assign new_n24892 = ~new_n24656 & ~new_n24891 ;
  assign new_n24893 = ~new_n24170 & ~new_n24892 ;
  assign new_n24894 = ~new_n24890 & ~new_n24893 ;
  assign new_n24895 = new_n24887 & new_n24894 ;
  assign new_n24896 = new_n24880 & new_n24895 ;
  assign new_n24897 = new_n24873 & new_n24896 ;
  assign new_n24898 = new_n24866 & new_n24897 ;
  assign new_n24899 = new_n24859 & new_n24898 ;
  assign new_n24900 = new_n24852 & new_n24899 ;
  assign new_n24901 = new_n24845 & new_n24900 ;
  assign new_n24902 = new_n24838 & new_n24901 ;
  assign new_n24903 = new_n24831 & new_n24902 ;
  assign new_n24904 = new_n24824 & new_n24903 ;
  assign new_n24905 = new_n24817 & new_n24904 ;
  assign new_n24906 = new_n24810 & new_n24905 ;
  assign new_n24907 = new_n24803 & new_n24906 ;
  assign new_n24908 = new_n24796 & new_n24907 ;
  assign new_n24909 = new_n24789 & new_n24908 ;
  assign new_n24910 = ~new_n24754 & new_n24909 ;
  assign new_n24911 = ~new_n24754 & ~new_n24910 ;
  assign new_n24912 = ~new_n24887 & ~new_n24894 ;
  assign new_n24913 = ~new_n24880 & new_n24912 ;
  assign new_n24914 = ~new_n24873 & new_n24913 ;
  assign new_n24915 = ~new_n24866 & new_n24914 ;
  assign new_n24916 = ~new_n24859 & new_n24915 ;
  assign new_n24917 = ~new_n24852 & new_n24916 ;
  assign new_n24918 = ~new_n24845 & new_n24917 ;
  assign new_n24919 = ~new_n24838 & new_n24918 ;
  assign new_n24920 = ~new_n24831 & new_n24919 ;
  assign new_n24921 = ~new_n24824 & new_n24920 ;
  assign new_n24922 = ~new_n24817 & new_n24921 ;
  assign new_n24923 = ~new_n24810 & new_n24922 ;
  assign new_n24924 = ~new_n24803 & new_n24923 ;
  assign new_n24925 = ~new_n24796 & new_n24924 ;
  assign new_n24926 = ~new_n24789 & new_n24925 ;
  assign new_n24927 = new_n24754 & ~new_n24926 ;
  assign new_n24928 = ~new_n24911 & ~new_n24927 ;
  assign new_n24929 = new_n24759 & new_n24766 ;
  assign new_n24930 = new_n24928 & ~new_n24929 ;
  assign new_n24931 = ~new_n21027 & ~new_n24930 ;
  assign new_n24932 = ~lo0941 & ~new_n24931 ;
  assign new_n24933 = ~new_n24782 & ~new_n24932 ;
  assign new_n24934 = ~new_n23174 & ~new_n24933 ;
  assign new_n24935 = ~new_n24768 & new_n24934 ;
  assign new_n24936 = ~new_n24768 & ~new_n24935 ;
  assign new_n24937 = ~new_n23239 & ~new_n24936 ;
  assign new_n24938 = new_n23239 & new_n24768 ;
  assign new_n24939 = ~new_n24934 & new_n24938 ;
  assign new_n24940 = ~new_n24937 & ~new_n24939 ;
  assign new_n24941 = ~new_n23175 & ~new_n24940 ;
  assign new_n24942 = ~new_n22707 & new_n23175 ;
  assign new_n24943 = ~new_n24941 & ~new_n24942 ;
  assign new_n24944 = ~new_n23177 & ~new_n24943 ;
  assign new_n24945 = ~new_n23178 & ~new_n24944 ;
  assign new_n24946 = lo1288 & ~new_n17706 ;
  assign new_n24947 = lo0955 & ~new_n13936 ;
  assign new_n24948 = ~lo0955 & ~new_n5455 ;
  assign new_n24949 = ~new_n24947 & ~new_n24948 ;
  assign new_n24950 = new_n17706 & ~new_n24949 ;
  assign new_n24951 = ~new_n24946 & ~new_n24950 ;
  assign new_n24952 = ~lo0944 & lo0948 ;
  assign new_n24953 = ~lo0947 & ~new_n24952 ;
  assign new_n24954 = ~lo0944 & lo0947 ;
  assign new_n24955 = lo0943 & ~lo0959 ;
  assign new_n24956 = new_n20793 & new_n24955 ;
  assign new_n24957 = ~new_n24954 & new_n24956 ;
  assign new_n24958 = ~new_n24953 & new_n24957 ;
  assign new_n24959 = new_n23174 & ~new_n24958 ;
  assign new_n24960 = lo0938 & new_n24028 ;
  assign new_n24961 = lo0962 & ~new_n2252 ;
  assign new_n24962 = ~new_n24960 & ~new_n24961 ;
  assign new_n24963 = ~new_n24959 & new_n24962 ;
  assign new_n24964 = lo1289 & new_n24963 ;
  assign new_n24965 = new_n24267 & new_n24607 ;
  assign new_n24966 = ~new_n24611 & ~new_n24965 ;
  assign new_n24967 = new_n24257 & ~new_n24966 ;
  assign new_n24968 = ~new_n24267 & new_n24607 ;
  assign new_n24969 = ~new_n24608 & ~new_n24968 ;
  assign new_n24970 = ~new_n24257 & ~new_n24969 ;
  assign new_n24971 = ~new_n24967 & ~new_n24970 ;
  assign new_n24972 = ~new_n24754 & ~new_n24757 ;
  assign new_n24973 = lo1408 & new_n24754 ;
  assign new_n24974 = new_n24026 & ~new_n24973 ;
  assign new_n24975 = ~new_n24972 & ~new_n24974 ;
  assign new_n24976 = ~lo0941 & ~new_n24975 ;
  assign new_n24977 = ~new_n24761 & ~new_n24976 ;
  assign new_n24978 = ~new_n24959 & ~new_n24977 ;
  assign new_n24979 = ~lo1410 & ~new_n24775 ;
  assign new_n24980 = new_n24365 & ~new_n24979 ;
  assign new_n24981 = ~new_n24365 & ~new_n24776 ;
  assign new_n24982 = ~new_n24980 & ~new_n24981 ;
  assign new_n24983 = lo0941 & ~new_n24982 ;
  assign new_n24984 = new_n24757 & ~new_n24763 ;
  assign new_n24985 = new_n24928 & ~new_n24984 ;
  assign new_n24986 = ~new_n21027 & ~new_n24985 ;
  assign new_n24987 = ~lo0941 & ~new_n24986 ;
  assign new_n24988 = ~new_n24983 & ~new_n24987 ;
  assign new_n24989 = ~new_n24959 & ~new_n24988 ;
  assign new_n24990 = ~new_n24978 & new_n24989 ;
  assign new_n24991 = ~new_n24978 & ~new_n24990 ;
  assign new_n24992 = ~new_n24971 & ~new_n24991 ;
  assign new_n24993 = new_n24971 & new_n24978 ;
  assign new_n24994 = ~new_n24989 & new_n24993 ;
  assign new_n24995 = ~new_n24992 & ~new_n24994 ;
  assign new_n24996 = ~new_n24961 & ~new_n24995 ;
  assign new_n24997 = ~new_n22332 & new_n24961 ;
  assign new_n24998 = ~new_n24996 & ~new_n24997 ;
  assign new_n24999 = ~new_n24963 & ~new_n24998 ;
  assign new_n25000 = ~new_n24964 & ~new_n24999 ;
  assign new_n25001 = lo1290 & new_n2252 ;
  assign new_n25002 = new_n12523 & new_n12713 ;
  assign new_n25003 = ~new_n12605 & ~new_n25002 ;
  assign new_n25004 = new_n12452 & new_n12526 ;
  assign new_n25005 = ~new_n25003 & new_n25004 ;
  assign new_n25006 = new_n15473 & ~new_n25005 ;
  assign new_n25007 = new_n2446 & ~new_n25006 ;
  assign new_n25008 = ~new_n2446 & new_n25006 ;
  assign new_n25009 = ~new_n25007 & ~new_n25008 ;
  assign new_n25010 = new_n13776 & ~new_n25009 ;
  assign new_n25011 = ~new_n13776 & new_n25007 ;
  assign new_n25012 = new_n12325 & ~new_n15481 ;
  assign new_n25013 = ~new_n12377 & ~new_n25012 ;
  assign new_n25014 = ~new_n2446 & new_n13782 ;
  assign new_n25015 = ~new_n25013 & new_n25014 ;
  assign new_n25016 = ~new_n25006 & new_n25015 ;
  assign new_n25017 = ~new_n25011 & ~new_n25016 ;
  assign new_n25018 = ~new_n25010 & new_n25017 ;
  assign new_n25019 = ~new_n2454 & new_n25018 ;
  assign new_n25020 = new_n25018 & ~new_n25019 ;
  assign new_n25021 = new_n12508 & ~new_n25020 ;
  assign new_n25022 = new_n2454 & ~new_n12508 ;
  assign new_n25023 = ~new_n25018 & new_n25022 ;
  assign new_n25024 = ~new_n25021 & ~new_n25023 ;
  assign new_n25025 = new_n2450 & ~new_n25024 ;
  assign new_n25026 = ~new_n15471 & ~new_n25025 ;
  assign new_n25027 = ~new_n2252 & ~new_n25026 ;
  assign new_n25028 = ~new_n25001 & ~new_n25027 ;
  assign new_n25029 = new_n12325 & new_n12338 ;
  assign new_n25030 = ~lo1292 & new_n12316 ;
  assign new_n25031 = lo1292 & ~new_n12325 ;
  assign new_n25032 = ~new_n25030 & ~new_n25031 ;
  assign new_n25033 = ~lo1291 & ~new_n25032 ;
  assign new_n25034 = ~new_n25029 & ~new_n25033 ;
  assign new_n25035 = new_n2262 & new_n12329 ;
  assign new_n25036 = ~new_n25034 & new_n25035 ;
  assign new_n25037 = ~new_n12377 & ~new_n12917 ;
  assign new_n25038 = ~new_n12329 & ~new_n25037 ;
  assign new_n25039 = ~new_n12375 & ~new_n25038 ;
  assign new_n25040 = ~new_n25036 & new_n25039 ;
  assign new_n25041 = new_n2455 & ~new_n25040 ;
  assign new_n25042 = ~new_n12384 & ~new_n15428 ;
  assign new_n25043 = new_n12402 & ~new_n25042 ;
  assign new_n25044 = new_n12408 & ~new_n25043 ;
  assign new_n25045 = ~new_n25041 & new_n25044 ;
  assign new_n25046 = ~new_n2446 & ~new_n25045 ;
  assign new_n25047 = ~new_n12504 & ~new_n25046 ;
  assign new_n25048 = new_n15452 & ~new_n25047 ;
  assign new_n25049 = new_n15452 & new_n25047 ;
  assign new_n25050 = lo1292 & new_n25049 ;
  assign new_n25051 = lo1291 & ~new_n25050 ;
  assign new_n25052 = ~lo1291 & new_n25050 ;
  assign new_n25053 = ~new_n25051 & ~new_n25052 ;
  assign new_n25054 = ~new_n25048 & ~new_n25053 ;
  assign new_n25055 = lo1292 & ~new_n25049 ;
  assign new_n25056 = ~lo1292 & new_n25049 ;
  assign new_n25057 = ~new_n25055 & ~new_n25056 ;
  assign new_n25058 = ~new_n25048 & ~new_n25057 ;
  assign new_n25059 = lo1291 & new_n25050 ;
  assign new_n25060 = lo1293 & ~new_n25059 ;
  assign new_n25061 = ~lo1293 & new_n25059 ;
  assign new_n25062 = ~new_n25060 & ~new_n25061 ;
  assign new_n25063 = ~new_n25048 & ~new_n25062 ;
  assign new_n25064 = lo1293 & new_n25059 ;
  assign new_n25065 = lo1294 & ~new_n25064 ;
  assign new_n25066 = ~lo1294 & new_n25064 ;
  assign new_n25067 = ~new_n25065 & ~new_n25066 ;
  assign new_n25068 = ~new_n25048 & ~new_n25067 ;
  assign new_n25069 = lo1295 & ~new_n17706 ;
  assign new_n25070 = lo0955 & ~new_n16735 ;
  assign new_n25071 = ~lo0955 & new_n6433 ;
  assign new_n25072 = ~new_n25070 & ~new_n25071 ;
  assign new_n25073 = new_n17706 & ~new_n25072 ;
  assign new_n25074 = ~new_n25069 & ~new_n25073 ;
  assign new_n25075 = lo1296 & new_n24963 ;
  assign new_n25076 = new_n24311 & new_n24583 ;
  assign new_n25077 = ~new_n24587 & ~new_n25076 ;
  assign new_n25078 = new_n24301 & ~new_n25077 ;
  assign new_n25079 = ~new_n24311 & new_n24583 ;
  assign new_n25080 = ~new_n24584 & ~new_n25079 ;
  assign new_n25081 = ~new_n24301 & ~new_n25080 ;
  assign new_n25082 = ~new_n25078 & ~new_n25081 ;
  assign new_n25083 = ~new_n24991 & ~new_n25082 ;
  assign new_n25084 = new_n24978 & new_n25082 ;
  assign new_n25085 = ~new_n24989 & new_n25084 ;
  assign new_n25086 = ~new_n25083 & ~new_n25085 ;
  assign new_n25087 = ~new_n24961 & ~new_n25086 ;
  assign new_n25088 = ~new_n22284 & new_n24961 ;
  assign new_n25089 = ~new_n25087 & ~new_n25088 ;
  assign new_n25090 = ~new_n24963 & ~new_n25089 ;
  assign new_n25091 = ~new_n25075 & ~new_n25090 ;
  assign new_n25092 = lo1297 & ~new_n23161 ;
  assign new_n25093 = lo0931 & ~new_n6433 ;
  assign new_n25094 = ~new_n6433 & ~new_n25093 ;
  assign new_n25095 = ~new_n16735 & ~new_n25094 ;
  assign new_n25096 = ~lo0931 & new_n6433 ;
  assign new_n25097 = new_n16735 & new_n25096 ;
  assign new_n25098 = ~new_n25095 & ~new_n25097 ;
  assign new_n25099 = ~lo0932 & ~new_n25098 ;
  assign new_n25100 = lo0226 & lo0932 ;
  assign new_n25101 = ~new_n25099 & ~new_n25100 ;
  assign new_n25102 = new_n23161 & ~new_n25101 ;
  assign new_n25103 = ~new_n25092 & ~new_n25102 ;
  assign new_n25104 = lo1298 & new_n23177 ;
  assign new_n25105 = ~lo1298 & new_n23206 ;
  assign new_n25106 = ~new_n23210 & ~new_n25105 ;
  assign new_n25107 = new_n23183 & ~new_n25106 ;
  assign new_n25108 = lo1298 & new_n23206 ;
  assign new_n25109 = ~new_n23207 & ~new_n25108 ;
  assign new_n25110 = ~new_n23183 & ~new_n25109 ;
  assign new_n25111 = ~new_n25107 & ~new_n25110 ;
  assign new_n25112 = ~new_n24936 & ~new_n25111 ;
  assign new_n25113 = new_n24768 & new_n25111 ;
  assign new_n25114 = ~new_n24934 & new_n25113 ;
  assign new_n25115 = ~new_n25112 & ~new_n25114 ;
  assign new_n25116 = ~new_n23175 & ~new_n25115 ;
  assign new_n25117 = ~new_n22635 & new_n23175 ;
  assign new_n25118 = ~new_n25116 & ~new_n25117 ;
  assign new_n25119 = ~new_n23177 & ~new_n25118 ;
  assign new_n25120 = ~new_n25104 & ~new_n25119 ;
  assign new_n25121 = lo1299 & new_n24963 ;
  assign new_n25122 = ~lo0941 & new_n24975 ;
  assign new_n25123 = ~new_n24761 & ~new_n25122 ;
  assign new_n25124 = ~new_n24959 & ~new_n25123 ;
  assign new_n25125 = new_n24989 & ~new_n25124 ;
  assign new_n25126 = ~new_n25124 & ~new_n25125 ;
  assign new_n25127 = ~new_n24859 & ~new_n25126 ;
  assign new_n25128 = new_n24859 & new_n25124 ;
  assign new_n25129 = ~new_n24989 & new_n25128 ;
  assign new_n25130 = ~new_n25127 & ~new_n25129 ;
  assign new_n25131 = ~new_n24961 & ~new_n25130 ;
  assign new_n25132 = ~new_n22452 & new_n24961 ;
  assign new_n25133 = ~new_n25131 & ~new_n25132 ;
  assign new_n25134 = ~new_n24963 & ~new_n25133 ;
  assign new_n25135 = ~new_n25121 & ~new_n25134 ;
  assign new_n25136 = lo1300 & ~new_n17706 ;
  assign new_n25137 = lo0955 & ~new_n14366 ;
  assign new_n25138 = ~lo0955 & new_n4257 ;
  assign new_n25139 = ~new_n25137 & ~new_n25138 ;
  assign new_n25140 = new_n17706 & ~new_n25139 ;
  assign new_n25141 = ~new_n25136 & ~new_n25140 ;
  assign new_n25142 = lo1301 & ~new_n23161 ;
  assign new_n25143 = lo0931 & ~new_n4257 ;
  assign new_n25144 = ~new_n4257 & ~new_n25143 ;
  assign new_n25145 = ~new_n14366 & ~new_n25144 ;
  assign new_n25146 = ~lo0931 & new_n4257 ;
  assign new_n25147 = new_n14366 & new_n25146 ;
  assign new_n25148 = ~new_n25145 & ~new_n25147 ;
  assign new_n25149 = ~lo0932 & ~new_n25148 ;
  assign new_n25150 = lo0245 & lo0932 ;
  assign new_n25151 = ~new_n25149 & ~new_n25150 ;
  assign new_n25152 = new_n23161 & ~new_n25151 ;
  assign new_n25153 = ~new_n25142 & ~new_n25152 ;
  assign new_n25154 = lo1302 & new_n23177 ;
  assign new_n25155 = ~lo1302 & new_n24487 ;
  assign new_n25156 = ~new_n24491 & ~new_n25155 ;
  assign new_n25157 = ~new_n24398 & ~new_n25156 ;
  assign new_n25158 = lo1302 & new_n24487 ;
  assign new_n25159 = ~new_n24488 & ~new_n25158 ;
  assign new_n25160 = new_n24398 & ~new_n25159 ;
  assign new_n25161 = ~new_n25157 & ~new_n25160 ;
  assign new_n25162 = ~new_n24936 & ~new_n25161 ;
  assign new_n25163 = new_n24768 & new_n25161 ;
  assign new_n25164 = ~new_n24934 & new_n25163 ;
  assign new_n25165 = ~new_n25162 & ~new_n25164 ;
  assign new_n25166 = ~new_n23175 & ~new_n25165 ;
  assign new_n25167 = ~new_n22644 & new_n23175 ;
  assign new_n25168 = ~new_n25166 & ~new_n25167 ;
  assign new_n25169 = ~new_n23177 & ~new_n25168 ;
  assign new_n25170 = ~new_n25154 & ~new_n25169 ;
  assign new_n25171 = lo1303 & ~new_n17706 ;
  assign new_n25172 = lo0955 & ~new_n14313 ;
  assign new_n25173 = ~lo0955 & new_n3538 ;
  assign new_n25174 = ~new_n25172 & ~new_n25173 ;
  assign new_n25175 = new_n17706 & ~new_n25174 ;
  assign new_n25176 = ~new_n25171 & ~new_n25175 ;
  assign new_n25177 = lo1304 & ~new_n17706 ;
  assign new_n25178 = lo0955 & ~new_n14154 ;
  assign new_n25179 = ~lo0955 & new_n3453 ;
  assign new_n25180 = ~new_n25178 & ~new_n25179 ;
  assign new_n25181 = new_n17706 & ~new_n25180 ;
  assign new_n25182 = ~new_n25177 & ~new_n25181 ;
  assign new_n25183 = lo1305 & ~new_n17706 ;
  assign new_n25184 = lo0955 & ~new_n14393 ;
  assign new_n25185 = ~lo0955 & new_n4619 ;
  assign new_n25186 = ~new_n25184 & ~new_n25185 ;
  assign new_n25187 = new_n17706 & ~new_n25186 ;
  assign new_n25188 = ~new_n25183 & ~new_n25187 ;
  assign new_n25189 = lo1306 & ~new_n17706 ;
  assign new_n25190 = lo0955 & ~new_n14419 ;
  assign new_n25191 = ~lo0955 & new_n4981 ;
  assign new_n25192 = ~new_n25190 & ~new_n25191 ;
  assign new_n25193 = new_n17706 & ~new_n25192 ;
  assign new_n25194 = ~new_n25189 & ~new_n25193 ;
  assign new_n25195 = lo1307 & ~new_n15033 ;
  assign new_n25196 = ~new_n14552 & new_n15036 ;
  assign new_n25197 = ~new_n4168 & ~new_n15036 ;
  assign new_n25198 = ~new_n25196 & ~new_n25197 ;
  assign new_n25199 = new_n15033 & ~new_n25198 ;
  assign new_n25200 = ~new_n25195 & ~new_n25199 ;
  assign new_n25201 = lo1308 & ~new_n17706 ;
  assign new_n25202 = lo0955 & ~new_n14340 ;
  assign new_n25203 = ~lo0955 & new_n3897 ;
  assign new_n25204 = ~new_n25202 & ~new_n25203 ;
  assign new_n25205 = new_n17706 & ~new_n25204 ;
  assign new_n25206 = ~new_n25201 & ~new_n25205 ;
  assign new_n25207 = lo1309 & ~new_n17706 ;
  assign new_n25208 = lo0955 & ~new_n16677 ;
  assign new_n25209 = ~lo0955 & ~new_n5743 ;
  assign new_n25210 = ~new_n25208 & ~new_n25209 ;
  assign new_n25211 = new_n17706 & ~new_n25210 ;
  assign new_n25212 = ~new_n25207 & ~new_n25211 ;
  assign new_n25213 = lo1310 & new_n23177 ;
  assign new_n25214 = ~lo1310 & new_n23224 ;
  assign new_n25215 = ~new_n23228 & ~new_n25214 ;
  assign new_n25216 = new_n23180 & ~new_n25215 ;
  assign new_n25217 = lo1310 & new_n23224 ;
  assign new_n25218 = ~new_n23225 & ~new_n25217 ;
  assign new_n25219 = ~new_n23180 & ~new_n25218 ;
  assign new_n25220 = ~new_n25216 & ~new_n25219 ;
  assign new_n25221 = ~new_n24936 & ~new_n25220 ;
  assign new_n25222 = new_n24768 & new_n25220 ;
  assign new_n25223 = ~new_n24934 & new_n25222 ;
  assign new_n25224 = ~new_n25221 & ~new_n25223 ;
  assign new_n25225 = ~new_n23175 & ~new_n25224 ;
  assign new_n25226 = ~new_n22689 & new_n23175 ;
  assign new_n25227 = ~new_n25225 & ~new_n25226 ;
  assign new_n25228 = ~new_n23177 & ~new_n25227 ;
  assign new_n25229 = ~new_n25213 & ~new_n25228 ;
  assign new_n25230 = lo1311 & new_n24963 ;
  assign new_n25231 = new_n24278 & new_n24601 ;
  assign new_n25232 = ~new_n24605 & ~new_n25231 ;
  assign new_n25233 = new_n24268 & ~new_n25232 ;
  assign new_n25234 = ~new_n24278 & new_n24601 ;
  assign new_n25235 = ~new_n24602 & ~new_n25234 ;
  assign new_n25236 = ~new_n24268 & ~new_n25235 ;
  assign new_n25237 = ~new_n25233 & ~new_n25236 ;
  assign new_n25238 = ~new_n24991 & ~new_n25237 ;
  assign new_n25239 = new_n24978 & new_n25237 ;
  assign new_n25240 = ~new_n24989 & new_n25239 ;
  assign new_n25241 = ~new_n25238 & ~new_n25240 ;
  assign new_n25242 = ~new_n24961 & ~new_n25241 ;
  assign new_n25243 = ~new_n22320 & new_n24961 ;
  assign new_n25244 = ~new_n25242 & ~new_n25243 ;
  assign new_n25245 = ~new_n24963 & ~new_n25244 ;
  assign new_n25246 = ~new_n25230 & ~new_n25245 ;
  assign new_n25247 = lo1312 & ~new_n23161 ;
  assign new_n25248 = lo0931 & new_n5743 ;
  assign new_n25249 = new_n5743 & ~new_n25248 ;
  assign new_n25250 = ~new_n16677 & ~new_n25249 ;
  assign new_n25251 = ~lo0931 & ~new_n5743 ;
  assign new_n25252 = new_n16677 & new_n25251 ;
  assign new_n25253 = ~new_n25250 & ~new_n25252 ;
  assign new_n25254 = ~lo0932 & ~new_n25253 ;
  assign new_n25255 = lo0399 & lo0932 ;
  assign new_n25256 = ~new_n25254 & ~new_n25255 ;
  assign new_n25257 = new_n23161 & ~new_n25256 ;
  assign new_n25258 = ~new_n25247 & ~new_n25257 ;
  assign new_n25259 = lo1313 & new_n24963 ;
  assign new_n25260 = ~new_n24887 & ~new_n25126 ;
  assign new_n25261 = new_n24887 & new_n25124 ;
  assign new_n25262 = ~new_n24989 & new_n25261 ;
  assign new_n25263 = ~new_n25260 & ~new_n25262 ;
  assign new_n25264 = ~new_n24961 & ~new_n25263 ;
  assign new_n25265 = ~new_n22103 & new_n24961 ;
  assign new_n25266 = ~new_n25264 & ~new_n25265 ;
  assign new_n25267 = ~new_n24963 & ~new_n25266 ;
  assign new_n25268 = ~new_n25259 & ~new_n25267 ;
  assign new_n25269 = lo1314 & ~new_n17706 ;
  assign new_n25270 = lo0955 & ~new_n14472 ;
  assign new_n25271 = ~lo0955 & new_n2899 ;
  assign new_n25272 = ~new_n25270 & ~new_n25271 ;
  assign new_n25273 = new_n17706 & ~new_n25272 ;
  assign new_n25274 = ~new_n25269 & ~new_n25273 ;
  assign new_n25275 = lo1315 & ~new_n23161 ;
  assign new_n25276 = lo0931 & ~new_n2899 ;
  assign new_n25277 = ~new_n2899 & ~new_n25276 ;
  assign new_n25278 = ~new_n14472 & ~new_n25277 ;
  assign new_n25279 = ~lo0931 & new_n2899 ;
  assign new_n25280 = new_n14472 & new_n25279 ;
  assign new_n25281 = ~new_n25278 & ~new_n25280 ;
  assign new_n25282 = ~lo0932 & ~new_n25281 ;
  assign new_n25283 = lo0417 & lo0932 ;
  assign new_n25284 = ~new_n25282 & ~new_n25283 ;
  assign new_n25285 = new_n23161 & ~new_n25284 ;
  assign new_n25286 = ~new_n25275 & ~new_n25285 ;
  assign new_n25287 = lo1316 & new_n23177 ;
  assign new_n25288 = ~lo1316 & new_n24457 ;
  assign new_n25289 = ~new_n24461 & ~new_n25288 ;
  assign new_n25290 = new_n24411 & ~new_n25289 ;
  assign new_n25291 = lo1316 & new_n24457 ;
  assign new_n25292 = ~new_n24458 & ~new_n25291 ;
  assign new_n25293 = ~new_n24411 & ~new_n25292 ;
  assign new_n25294 = ~new_n25290 & ~new_n25293 ;
  assign new_n25295 = ~new_n24936 & ~new_n25294 ;
  assign new_n25296 = new_n24768 & new_n25294 ;
  assign new_n25297 = ~new_n24934 & new_n25296 ;
  assign new_n25298 = ~new_n25295 & ~new_n25297 ;
  assign new_n25299 = ~new_n23175 & ~new_n25298 ;
  assign new_n25300 = ~new_n22091 & new_n23175 ;
  assign new_n25301 = ~new_n25299 & ~new_n25300 ;
  assign new_n25302 = ~new_n23177 & ~new_n25301 ;
  assign new_n25303 = ~new_n25287 & ~new_n25302 ;
  assign new_n25304 = lo1317 & ~new_n17706 ;
  assign new_n25305 = lo0955 & ~new_n14499 ;
  assign new_n25306 = ~lo0955 & ~new_n3372 ;
  assign new_n25307 = ~new_n25305 & ~new_n25306 ;
  assign new_n25308 = new_n17706 & ~new_n25307 ;
  assign new_n25309 = ~new_n25304 & ~new_n25308 ;
  assign new_n25310 = lo1318 & ~new_n17706 ;
  assign new_n25311 = lo0955 & ~new_n14128 ;
  assign new_n25312 = ~lo0955 & new_n2990 ;
  assign new_n25313 = ~new_n25311 & ~new_n25312 ;
  assign new_n25314 = new_n17706 & ~new_n25313 ;
  assign new_n25315 = ~new_n25310 & ~new_n25314 ;
  assign new_n25316 = lo1319 & ~new_n17706 ;
  assign new_n25317 = lo0955 & ~new_n14060 ;
  assign new_n25318 = ~lo0955 & new_n2718 ;
  assign new_n25319 = ~new_n25317 & ~new_n25318 ;
  assign new_n25320 = new_n17706 & ~new_n25319 ;
  assign new_n25321 = ~new_n25316 & ~new_n25320 ;
  assign new_n25322 = lo1320 & ~new_n17706 ;
  assign new_n25323 = lo0955 & ~new_n14101 ;
  assign new_n25324 = ~lo0955 & new_n3081 ;
  assign new_n25325 = ~new_n25323 & ~new_n25324 ;
  assign new_n25326 = new_n17706 & ~new_n25325 ;
  assign new_n25327 = ~new_n25322 & ~new_n25326 ;
  assign new_n25328 = lo1321 & new_n23177 ;
  assign new_n25329 = ~lo1321 & new_n23218 ;
  assign new_n25330 = ~new_n23222 & ~new_n25329 ;
  assign new_n25331 = new_n23181 & ~new_n25330 ;
  assign new_n25332 = lo1321 & new_n23218 ;
  assign new_n25333 = ~new_n23219 & ~new_n25332 ;
  assign new_n25334 = ~new_n23181 & ~new_n25333 ;
  assign new_n25335 = ~new_n25331 & ~new_n25334 ;
  assign new_n25336 = ~new_n24936 & ~new_n25335 ;
  assign new_n25337 = new_n24768 & new_n25335 ;
  assign new_n25338 = ~new_n24934 & new_n25337 ;
  assign new_n25339 = ~new_n25336 & ~new_n25338 ;
  assign new_n25340 = ~new_n23175 & ~new_n25339 ;
  assign new_n25341 = ~new_n22671 & new_n23175 ;
  assign new_n25342 = ~new_n25340 & ~new_n25341 ;
  assign new_n25343 = ~new_n23177 & ~new_n25342 ;
  assign new_n25344 = ~new_n25328 & ~new_n25343 ;
  assign new_n25345 = lo1322 & ~new_n17706 ;
  assign new_n25346 = lo0955 & ~new_n16697 ;
  assign new_n25347 = ~lo0955 & new_n5977 ;
  assign new_n25348 = ~new_n25346 & ~new_n25347 ;
  assign new_n25349 = new_n17706 & ~new_n25348 ;
  assign new_n25350 = ~new_n25345 & ~new_n25349 ;
  assign new_n25351 = lo1323 & new_n24963 ;
  assign new_n25352 = new_n24289 & new_n24595 ;
  assign new_n25353 = ~new_n24599 & ~new_n25352 ;
  assign new_n25354 = new_n24279 & ~new_n25353 ;
  assign new_n25355 = ~new_n24289 & new_n24595 ;
  assign new_n25356 = ~new_n24596 & ~new_n25355 ;
  assign new_n25357 = ~new_n24279 & ~new_n25356 ;
  assign new_n25358 = ~new_n25354 & ~new_n25357 ;
  assign new_n25359 = ~new_n24991 & ~new_n25358 ;
  assign new_n25360 = new_n24978 & new_n25358 ;
  assign new_n25361 = ~new_n24989 & new_n25360 ;
  assign new_n25362 = ~new_n25359 & ~new_n25361 ;
  assign new_n25363 = ~new_n24961 & ~new_n25362 ;
  assign new_n25364 = ~new_n22308 & new_n24961 ;
  assign new_n25365 = ~new_n25363 & ~new_n25364 ;
  assign new_n25366 = ~new_n24963 & ~new_n25365 ;
  assign new_n25367 = ~new_n25351 & ~new_n25366 ;
  assign new_n25368 = lo1324 & ~new_n23161 ;
  assign new_n25369 = lo0931 & ~new_n5977 ;
  assign new_n25370 = ~new_n5977 & ~new_n25369 ;
  assign new_n25371 = ~new_n16697 & ~new_n25370 ;
  assign new_n25372 = ~lo0931 & new_n5977 ;
  assign new_n25373 = new_n16697 & new_n25372 ;
  assign new_n25374 = ~new_n25371 & ~new_n25373 ;
  assign new_n25375 = ~lo0932 & ~new_n25374 ;
  assign new_n25376 = lo0516 & lo0932 ;
  assign new_n25377 = ~new_n25375 & ~new_n25376 ;
  assign new_n25378 = new_n23161 & ~new_n25377 ;
  assign new_n25379 = ~new_n25368 & ~new_n25378 ;
  assign new_n25380 = lo1325 & new_n24963 ;
  assign new_n25381 = new_n24201 & new_n24643 ;
  assign new_n25382 = ~new_n24647 & ~new_n25381 ;
  assign new_n25383 = new_n24191 & ~new_n25382 ;
  assign new_n25384 = ~new_n24201 & new_n24643 ;
  assign new_n25385 = ~new_n24644 & ~new_n25384 ;
  assign new_n25386 = ~new_n24191 & ~new_n25385 ;
  assign new_n25387 = ~new_n25383 & ~new_n25386 ;
  assign new_n25388 = ~new_n24991 & ~new_n25387 ;
  assign new_n25389 = new_n24978 & new_n25387 ;
  assign new_n25390 = ~new_n24989 & new_n25389 ;
  assign new_n25391 = ~new_n25388 & ~new_n25390 ;
  assign new_n25392 = ~new_n24961 & ~new_n25391 ;
  assign new_n25393 = ~new_n22404 & new_n24961 ;
  assign new_n25394 = ~new_n25392 & ~new_n25393 ;
  assign new_n25395 = ~new_n24963 & ~new_n25394 ;
  assign new_n25396 = ~new_n25380 & ~new_n25395 ;
  assign new_n25397 = lo1326 & ~new_n23161 ;
  assign new_n25398 = lo0931 & new_n3372 ;
  assign new_n25399 = new_n3372 & ~new_n25398 ;
  assign new_n25400 = ~new_n14499 & ~new_n25399 ;
  assign new_n25401 = ~lo0931 & ~new_n3372 ;
  assign new_n25402 = new_n14499 & new_n25401 ;
  assign new_n25403 = ~new_n25400 & ~new_n25402 ;
  assign new_n25404 = ~lo0932 & ~new_n25403 ;
  assign new_n25405 = lo0437 & lo0932 ;
  assign new_n25406 = ~new_n25404 & ~new_n25405 ;
  assign new_n25407 = new_n23161 & ~new_n25406 ;
  assign new_n25408 = ~new_n25397 & ~new_n25407 ;
  assign new_n25409 = lo1327 & new_n23177 ;
  assign new_n25410 = ~lo1327 & new_n24451 ;
  assign new_n25411 = ~new_n24455 & ~new_n25410 ;
  assign new_n25412 = new_n24412 & ~new_n25411 ;
  assign new_n25413 = lo1327 & new_n24451 ;
  assign new_n25414 = ~new_n24452 & ~new_n25413 ;
  assign new_n25415 = ~new_n24412 & ~new_n25414 ;
  assign new_n25416 = ~new_n25412 & ~new_n25415 ;
  assign new_n25417 = ~new_n24936 & ~new_n25416 ;
  assign new_n25418 = new_n24768 & new_n25416 ;
  assign new_n25419 = ~new_n24934 & new_n25418 ;
  assign new_n25420 = ~new_n25417 & ~new_n25419 ;
  assign new_n25421 = ~new_n23175 & ~new_n25420 ;
  assign new_n25422 = ~new_n22815 & new_n23175 ;
  assign new_n25423 = ~new_n25421 & ~new_n25422 ;
  assign new_n25424 = ~new_n23177 & ~new_n25423 ;
  assign new_n25425 = ~new_n25409 & ~new_n25424 ;
  assign new_n25426 = lo1328 & ~new_n17706 ;
  assign new_n25427 = lo0955 & ~new_n14005 ;
  assign new_n25428 = ~lo0955 & ~new_n3723 ;
  assign new_n25429 = ~new_n25427 & ~new_n25428 ;
  assign new_n25430 = new_n17706 & ~new_n25429 ;
  assign new_n25431 = ~new_n25426 & ~new_n25430 ;
  assign new_n25432 = lo1329 & ~new_n17706 ;
  assign new_n25433 = lo0955 & ~new_n14036 ;
  assign new_n25434 = ~lo0955 & new_n5549 ;
  assign new_n25435 = ~new_n25433 & ~new_n25434 ;
  assign new_n25436 = new_n17706 & ~new_n25435 ;
  assign new_n25437 = ~new_n25432 & ~new_n25436 ;
  assign new_n25438 = lo1330 & new_n24963 ;
  assign new_n25439 = ~new_n24789 & ~new_n25126 ;
  assign new_n25440 = new_n24789 & new_n25124 ;
  assign new_n25441 = ~new_n24989 & new_n25440 ;
  assign new_n25442 = ~new_n25439 & ~new_n25441 ;
  assign new_n25443 = ~new_n24961 & ~new_n25442 ;
  assign new_n25444 = ~new_n22572 & new_n24961 ;
  assign new_n25445 = ~new_n25443 & ~new_n25444 ;
  assign new_n25446 = ~new_n24963 & ~new_n25445 ;
  assign new_n25447 = ~new_n25438 & ~new_n25446 ;
  assign new_n25448 = lo1331 & ~new_n23161 ;
  assign new_n25449 = lo0931 & ~new_n3081 ;
  assign new_n25450 = ~new_n3081 & ~new_n25449 ;
  assign new_n25451 = ~new_n14101 & ~new_n25450 ;
  assign new_n25452 = ~lo0931 & new_n3081 ;
  assign new_n25453 = new_n14101 & new_n25452 ;
  assign new_n25454 = ~new_n25451 & ~new_n25453 ;
  assign new_n25455 = ~lo0932 & ~new_n25454 ;
  assign new_n25456 = lo0495 & lo0932 ;
  assign new_n25457 = ~new_n25455 & ~new_n25456 ;
  assign new_n25458 = new_n23161 & ~new_n25457 ;
  assign new_n25459 = ~new_n25448 & ~new_n25458 ;
  assign new_n25460 = lo1332 & new_n23177 ;
  assign new_n25461 = ~lo1332 & new_n24547 ;
  assign new_n25462 = ~new_n24551 & ~new_n25461 ;
  assign new_n25463 = ~new_n24368 & ~new_n25462 ;
  assign new_n25464 = lo1332 & new_n24547 ;
  assign new_n25465 = ~new_n24548 & ~new_n25464 ;
  assign new_n25466 = new_n24368 & ~new_n25465 ;
  assign new_n25467 = ~new_n25463 & ~new_n25466 ;
  assign new_n25468 = ~new_n24936 & ~new_n25467 ;
  assign new_n25469 = new_n24768 & new_n25467 ;
  assign new_n25470 = ~new_n24934 & new_n25469 ;
  assign new_n25471 = ~new_n25468 & ~new_n25470 ;
  assign new_n25472 = ~new_n23175 & ~new_n25471 ;
  assign new_n25473 = ~new_n22824 & new_n23175 ;
  assign new_n25474 = ~new_n25472 & ~new_n25473 ;
  assign new_n25475 = ~new_n23177 & ~new_n25474 ;
  assign new_n25476 = ~new_n25460 & ~new_n25475 ;
  assign new_n25477 = lo1333 & ~new_n17706 ;
  assign new_n25478 = lo0955 & ~new_n18863 ;
  assign new_n25479 = ~lo0955 & new_n6667 ;
  assign new_n25480 = ~new_n25478 & ~new_n25479 ;
  assign new_n25481 = new_n17706 & ~new_n25480 ;
  assign new_n25482 = ~new_n25477 & ~new_n25481 ;
  assign new_n25483 = lo1334 & ~new_n17706 ;
  assign new_n25484 = lo0955 & ~new_n16716 ;
  assign new_n25485 = ~lo0955 & new_n6202 ;
  assign new_n25486 = ~new_n25484 & ~new_n25485 ;
  assign new_n25487 = new_n17706 & ~new_n25486 ;
  assign new_n25488 = ~new_n25483 & ~new_n25487 ;
  assign new_n25489 = lo1335 & new_n24963 ;
  assign new_n25490 = new_n24300 & new_n24589 ;
  assign new_n25491 = ~new_n24593 & ~new_n25490 ;
  assign new_n25492 = new_n24290 & ~new_n25491 ;
  assign new_n25493 = ~new_n24300 & new_n24589 ;
  assign new_n25494 = ~new_n24590 & ~new_n25493 ;
  assign new_n25495 = ~new_n24290 & ~new_n25494 ;
  assign new_n25496 = ~new_n25492 & ~new_n25495 ;
  assign new_n25497 = ~new_n24991 & ~new_n25496 ;
  assign new_n25498 = new_n24978 & new_n25496 ;
  assign new_n25499 = ~new_n24989 & new_n25498 ;
  assign new_n25500 = ~new_n25497 & ~new_n25499 ;
  assign new_n25501 = ~new_n24961 & ~new_n25500 ;
  assign new_n25502 = ~new_n22296 & new_n24961 ;
  assign new_n25503 = ~new_n25501 & ~new_n25502 ;
  assign new_n25504 = ~new_n24963 & ~new_n25503 ;
  assign new_n25505 = ~new_n25489 & ~new_n25504 ;
  assign new_n25506 = lo1336 & ~new_n23161 ;
  assign new_n25507 = lo0931 & ~new_n6202 ;
  assign new_n25508 = ~new_n6202 & ~new_n25507 ;
  assign new_n25509 = ~new_n16716 & ~new_n25508 ;
  assign new_n25510 = ~lo0931 & new_n6202 ;
  assign new_n25511 = new_n16716 & new_n25510 ;
  assign new_n25512 = ~new_n25509 & ~new_n25511 ;
  assign new_n25513 = ~lo0932 & ~new_n25512 ;
  assign new_n25514 = lo0600 & lo0932 ;
  assign new_n25515 = ~new_n25513 & ~new_n25514 ;
  assign new_n25516 = new_n23161 & ~new_n25515 ;
  assign new_n25517 = ~new_n25506 & ~new_n25516 ;
  assign new_n25518 = lo1337 & new_n23177 ;
  assign new_n25519 = ~lo1337 & new_n23212 ;
  assign new_n25520 = ~new_n23216 & ~new_n25519 ;
  assign new_n25521 = new_n23182 & ~new_n25520 ;
  assign new_n25522 = lo1337 & new_n23212 ;
  assign new_n25523 = ~new_n23213 & ~new_n25522 ;
  assign new_n25524 = ~new_n23182 & ~new_n25523 ;
  assign new_n25525 = ~new_n25521 & ~new_n25524 ;
  assign new_n25526 = ~new_n24936 & ~new_n25525 ;
  assign new_n25527 = new_n24768 & new_n25525 ;
  assign new_n25528 = ~new_n24934 & new_n25527 ;
  assign new_n25529 = ~new_n25526 & ~new_n25528 ;
  assign new_n25530 = ~new_n23175 & ~new_n25529 ;
  assign new_n25531 = ~new_n22653 & new_n23175 ;
  assign new_n25532 = ~new_n25530 & ~new_n25531 ;
  assign new_n25533 = ~new_n23177 & ~new_n25532 ;
  assign new_n25534 = ~new_n25518 & ~new_n25533 ;
  assign new_n25535 = lo1338 & new_n24963 ;
  assign new_n25536 = new_n24212 & new_n24637 ;
  assign new_n25537 = ~new_n24641 & ~new_n25536 ;
  assign new_n25538 = new_n24202 & ~new_n25537 ;
  assign new_n25539 = ~new_n24212 & new_n24637 ;
  assign new_n25540 = ~new_n24638 & ~new_n25539 ;
  assign new_n25541 = ~new_n24202 & ~new_n25540 ;
  assign new_n25542 = ~new_n25538 & ~new_n25541 ;
  assign new_n25543 = ~new_n24991 & ~new_n25542 ;
  assign new_n25544 = new_n24978 & new_n25542 ;
  assign new_n25545 = ~new_n24989 & new_n25544 ;
  assign new_n25546 = ~new_n25543 & ~new_n25545 ;
  assign new_n25547 = ~new_n24961 & ~new_n25546 ;
  assign new_n25548 = ~new_n22392 & new_n24961 ;
  assign new_n25549 = ~new_n25547 & ~new_n25548 ;
  assign new_n25550 = ~new_n24963 & ~new_n25549 ;
  assign new_n25551 = ~new_n25535 & ~new_n25550 ;
  assign new_n25552 = lo1339 & ~new_n23161 ;
  assign new_n25553 = lo0931 & new_n3723 ;
  assign new_n25554 = new_n3723 & ~new_n25553 ;
  assign new_n25555 = ~new_n14005 & ~new_n25554 ;
  assign new_n25556 = ~lo0931 & ~new_n3723 ;
  assign new_n25557 = new_n14005 & new_n25556 ;
  assign new_n25558 = ~new_n25555 & ~new_n25557 ;
  assign new_n25559 = ~lo0932 & ~new_n25558 ;
  assign new_n25560 = lo0535 & lo0932 ;
  assign new_n25561 = ~new_n25559 & ~new_n25560 ;
  assign new_n25562 = new_n23161 & ~new_n25561 ;
  assign new_n25563 = ~new_n25552 & ~new_n25562 ;
  assign new_n25564 = lo1340 & new_n23177 ;
  assign new_n25565 = ~lo1340 & new_n24445 ;
  assign new_n25566 = ~new_n24449 & ~new_n25565 ;
  assign new_n25567 = new_n24413 & ~new_n25566 ;
  assign new_n25568 = lo1340 & new_n24445 ;
  assign new_n25569 = ~new_n24446 & ~new_n25568 ;
  assign new_n25570 = ~new_n24413 & ~new_n25569 ;
  assign new_n25571 = ~new_n25567 & ~new_n25570 ;
  assign new_n25572 = ~new_n24936 & ~new_n25571 ;
  assign new_n25573 = new_n24768 & new_n25571 ;
  assign new_n25574 = ~new_n24934 & new_n25573 ;
  assign new_n25575 = ~new_n25572 & ~new_n25574 ;
  assign new_n25576 = ~new_n23175 & ~new_n25575 ;
  assign new_n25577 = ~new_n22797 & new_n23175 ;
  assign new_n25578 = ~new_n25576 & ~new_n25577 ;
  assign new_n25579 = ~new_n23177 & ~new_n25578 ;
  assign new_n25580 = ~new_n25564 & ~new_n25579 ;
  assign new_n25581 = lo1341 & new_n24963 ;
  assign new_n25582 = ~new_n24852 & ~new_n25126 ;
  assign new_n25583 = new_n24852 & new_n25124 ;
  assign new_n25584 = ~new_n24989 & new_n25583 ;
  assign new_n25585 = ~new_n25582 & ~new_n25584 ;
  assign new_n25586 = ~new_n24961 & ~new_n25585 ;
  assign new_n25587 = ~new_n22464 & new_n24961 ;
  assign new_n25588 = ~new_n25586 & ~new_n25587 ;
  assign new_n25589 = ~new_n24963 & ~new_n25588 ;
  assign new_n25590 = ~new_n25581 & ~new_n25589 ;
  assign new_n25591 = lo1342 & ~new_n23161 ;
  assign new_n25592 = lo0931 & ~new_n3897 ;
  assign new_n25593 = ~new_n3897 & ~new_n25592 ;
  assign new_n25594 = ~new_n14340 & ~new_n25593 ;
  assign new_n25595 = ~lo0931 & new_n3897 ;
  assign new_n25596 = new_n14340 & new_n25595 ;
  assign new_n25597 = ~new_n25594 & ~new_n25596 ;
  assign new_n25598 = ~lo0932 & ~new_n25597 ;
  assign new_n25599 = lo0378 & lo0932 ;
  assign new_n25600 = ~new_n25598 & ~new_n25599 ;
  assign new_n25601 = new_n23161 & ~new_n25600 ;
  assign new_n25602 = ~new_n25591 & ~new_n25601 ;
  assign new_n25603 = lo1343 & new_n23177 ;
  assign new_n25604 = ~lo1343 & new_n24493 ;
  assign new_n25605 = ~new_n24497 & ~new_n25604 ;
  assign new_n25606 = ~new_n24395 & ~new_n25605 ;
  assign new_n25607 = lo1343 & new_n24493 ;
  assign new_n25608 = ~new_n24494 & ~new_n25607 ;
  assign new_n25609 = new_n24395 & ~new_n25608 ;
  assign new_n25610 = ~new_n25606 & ~new_n25609 ;
  assign new_n25611 = ~new_n24936 & ~new_n25610 ;
  assign new_n25612 = new_n24768 & new_n25610 ;
  assign new_n25613 = ~new_n24934 & new_n25612 ;
  assign new_n25614 = ~new_n25611 & ~new_n25613 ;
  assign new_n25615 = ~new_n23175 & ~new_n25614 ;
  assign new_n25616 = ~new_n22662 & new_n23175 ;
  assign new_n25617 = ~new_n25615 & ~new_n25616 ;
  assign new_n25618 = ~new_n23177 & ~new_n25617 ;
  assign new_n25619 = ~new_n25603 & ~new_n25618 ;
  assign new_n25620 = lo1344 & ~new_n17706 ;
  assign new_n25621 = lo0955 & ~new_n14287 ;
  assign new_n25622 = ~lo0955 & new_n2813 ;
  assign new_n25623 = ~new_n25621 & ~new_n25622 ;
  assign new_n25624 = new_n17706 & ~new_n25623 ;
  assign new_n25625 = ~new_n25620 & ~new_n25624 ;
  assign new_n25626 = lo1345 & new_n24963 ;
  assign new_n25627 = new_n24223 & new_n24631 ;
  assign new_n25628 = ~new_n24635 & ~new_n25627 ;
  assign new_n25629 = new_n24213 & ~new_n25628 ;
  assign new_n25630 = ~new_n24223 & new_n24631 ;
  assign new_n25631 = ~new_n24632 & ~new_n25630 ;
  assign new_n25632 = ~new_n24213 & ~new_n25631 ;
  assign new_n25633 = ~new_n25629 & ~new_n25632 ;
  assign new_n25634 = ~new_n24991 & ~new_n25633 ;
  assign new_n25635 = new_n24978 & new_n25633 ;
  assign new_n25636 = ~new_n24989 & new_n25635 ;
  assign new_n25637 = ~new_n25634 & ~new_n25636 ;
  assign new_n25638 = ~new_n24961 & ~new_n25637 ;
  assign new_n25639 = ~new_n22380 & new_n24961 ;
  assign new_n25640 = ~new_n25638 & ~new_n25639 ;
  assign new_n25641 = ~new_n24963 & ~new_n25640 ;
  assign new_n25642 = ~new_n25626 & ~new_n25641 ;
  assign new_n25643 = lo1346 & ~new_n23161 ;
  assign new_n25644 = lo0931 & new_n4168 ;
  assign new_n25645 = new_n4168 & ~new_n25644 ;
  assign new_n25646 = ~new_n14552 & ~new_n25645 ;
  assign new_n25647 = ~lo0931 & ~new_n4168 ;
  assign new_n25648 = new_n14552 & new_n25647 ;
  assign new_n25649 = ~new_n25646 & ~new_n25648 ;
  assign new_n25650 = ~lo0932 & ~new_n25649 ;
  assign new_n25651 = lo0357 & lo0932 ;
  assign new_n25652 = ~new_n25650 & ~new_n25651 ;
  assign new_n25653 = new_n23161 & ~new_n25652 ;
  assign new_n25654 = ~new_n25643 & ~new_n25653 ;
  assign new_n25655 = lo1347 & new_n23177 ;
  assign new_n25656 = ~lo1347 & new_n24439 ;
  assign new_n25657 = ~new_n24443 & ~new_n25656 ;
  assign new_n25658 = new_n24414 & ~new_n25657 ;
  assign new_n25659 = lo1347 & new_n24439 ;
  assign new_n25660 = ~new_n24440 & ~new_n25659 ;
  assign new_n25661 = ~new_n24414 & ~new_n25660 ;
  assign new_n25662 = ~new_n25658 & ~new_n25661 ;
  assign new_n25663 = ~new_n24936 & ~new_n25662 ;
  assign new_n25664 = new_n24768 & new_n25662 ;
  assign new_n25665 = ~new_n24934 & new_n25664 ;
  assign new_n25666 = ~new_n25663 & ~new_n25665 ;
  assign new_n25667 = ~new_n23175 & ~new_n25666 ;
  assign new_n25668 = ~new_n22779 & new_n23175 ;
  assign new_n25669 = ~new_n25667 & ~new_n25668 ;
  assign new_n25670 = ~new_n23177 & ~new_n25669 ;
  assign new_n25671 = ~new_n25655 & ~new_n25670 ;
  assign new_n25672 = lo1348 & ~new_n17706 ;
  assign new_n25673 = lo0955 & ~new_n19223 ;
  assign new_n25674 = ~lo0955 & new_n6899 ;
  assign new_n25675 = ~new_n25673 & ~new_n25674 ;
  assign new_n25676 = new_n17706 & ~new_n25675 ;
  assign new_n25677 = ~new_n25672 & ~new_n25676 ;
  assign new_n25678 = lo1349 & ~new_n17706 ;
  assign new_n25679 = lo0955 & ~new_n14181 ;
  assign new_n25680 = ~lo0955 & new_n3806 ;
  assign new_n25681 = ~new_n25679 & ~new_n25680 ;
  assign new_n25682 = new_n17706 & ~new_n25681 ;
  assign new_n25683 = ~new_n25678 & ~new_n25682 ;
  assign new_n25684 = lo1350 & ~new_n17706 ;
  assign new_n25685 = lo0955 & ~new_n14207 ;
  assign new_n25686 = ~lo0955 & new_n4086 ;
  assign new_n25687 = ~new_n25685 & ~new_n25686 ;
  assign new_n25688 = new_n17706 & ~new_n25687 ;
  assign new_n25689 = ~new_n25684 & ~new_n25688 ;
  assign new_n25690 = lo1351 & ~new_n15033 ;
  assign new_n25691 = ~new_n14525 & new_n15036 ;
  assign new_n25692 = ~new_n4889 & ~new_n15036 ;
  assign new_n25693 = ~new_n25691 & ~new_n25692 ;
  assign new_n25694 = new_n15033 & ~new_n25693 ;
  assign new_n25695 = ~new_n25690 & ~new_n25694 ;
  assign new_n25696 = lo1352 & ~new_n17706 ;
  assign new_n25697 = lo0955 & ~new_n14578 ;
  assign new_n25698 = ~lo0955 & ~new_n4446 ;
  assign new_n25699 = ~new_n25697 & ~new_n25698 ;
  assign new_n25700 = new_n17706 & ~new_n25699 ;
  assign new_n25701 = ~new_n25696 & ~new_n25700 ;
  assign new_n25702 = lo1353 & new_n24963 ;
  assign new_n25703 = ~new_n24803 & ~new_n25126 ;
  assign new_n25704 = new_n24803 & new_n25124 ;
  assign new_n25705 = ~new_n24989 & new_n25704 ;
  assign new_n25706 = ~new_n25703 & ~new_n25705 ;
  assign new_n25707 = ~new_n24961 & ~new_n25706 ;
  assign new_n25708 = ~new_n22548 & new_n24961 ;
  assign new_n25709 = ~new_n25707 & ~new_n25708 ;
  assign new_n25710 = ~new_n24963 & ~new_n25709 ;
  assign new_n25711 = ~new_n25702 & ~new_n25710 ;
  assign new_n25712 = lo1354 & ~new_n23161 ;
  assign new_n25713 = lo0931 & ~new_n3453 ;
  assign new_n25714 = ~new_n3453 & ~new_n25713 ;
  assign new_n25715 = ~new_n14154 & ~new_n25714 ;
  assign new_n25716 = ~lo0931 & new_n3453 ;
  assign new_n25717 = new_n14154 & new_n25716 ;
  assign new_n25718 = ~new_n25715 & ~new_n25717 ;
  assign new_n25719 = ~lo0932 & ~new_n25718 ;
  assign new_n25720 = lo0294 & lo0932 ;
  assign new_n25721 = ~new_n25719 & ~new_n25720 ;
  assign new_n25722 = new_n23161 & ~new_n25721 ;
  assign new_n25723 = ~new_n25712 & ~new_n25722 ;
  assign new_n25724 = lo1355 & new_n23177 ;
  assign new_n25725 = ~lo1355 & new_n24535 ;
  assign new_n25726 = ~new_n24539 & ~new_n25725 ;
  assign new_n25727 = ~new_n24374 & ~new_n25726 ;
  assign new_n25728 = lo1355 & new_n24535 ;
  assign new_n25729 = ~new_n24536 & ~new_n25728 ;
  assign new_n25730 = new_n24374 & ~new_n25729 ;
  assign new_n25731 = ~new_n25727 & ~new_n25730 ;
  assign new_n25732 = ~new_n24936 & ~new_n25731 ;
  assign new_n25733 = new_n24768 & new_n25731 ;
  assign new_n25734 = ~new_n24934 & new_n25733 ;
  assign new_n25735 = ~new_n25732 & ~new_n25734 ;
  assign new_n25736 = ~new_n23175 & ~new_n25735 ;
  assign new_n25737 = ~new_n22788 & new_n23175 ;
  assign new_n25738 = ~new_n25736 & ~new_n25737 ;
  assign new_n25739 = ~new_n23177 & ~new_n25738 ;
  assign new_n25740 = ~new_n25724 & ~new_n25739 ;
  assign new_n25741 = lo1356 & new_n24963 ;
  assign new_n25742 = ~new_n24845 & ~new_n25126 ;
  assign new_n25743 = new_n24845 & new_n25124 ;
  assign new_n25744 = ~new_n24989 & new_n25743 ;
  assign new_n25745 = ~new_n25742 & ~new_n25744 ;
  assign new_n25746 = ~new_n24961 & ~new_n25745 ;
  assign new_n25747 = ~new_n22476 & new_n24961 ;
  assign new_n25748 = ~new_n25746 & ~new_n25747 ;
  assign new_n25749 = ~new_n24963 & ~new_n25748 ;
  assign new_n25750 = ~new_n25741 & ~new_n25749 ;
  assign new_n25751 = lo1357 & ~new_n23161 ;
  assign new_n25752 = lo0931 & ~new_n3538 ;
  assign new_n25753 = ~new_n3538 & ~new_n25752 ;
  assign new_n25754 = ~new_n14313 & ~new_n25753 ;
  assign new_n25755 = ~lo0931 & new_n3538 ;
  assign new_n25756 = new_n14313 & new_n25755 ;
  assign new_n25757 = ~new_n25754 & ~new_n25756 ;
  assign new_n25758 = ~lo0932 & ~new_n25757 ;
  assign new_n25759 = lo0275 & lo0932 ;
  assign new_n25760 = ~new_n25758 & ~new_n25759 ;
  assign new_n25761 = new_n23161 & ~new_n25760 ;
  assign new_n25762 = ~new_n25751 & ~new_n25761 ;
  assign new_n25763 = lo1358 & new_n23177 ;
  assign new_n25764 = ~lo1358 & new_n24499 ;
  assign new_n25765 = ~new_n24503 & ~new_n25764 ;
  assign new_n25766 = ~new_n24392 & ~new_n25765 ;
  assign new_n25767 = lo1358 & new_n24499 ;
  assign new_n25768 = ~new_n24500 & ~new_n25767 ;
  assign new_n25769 = new_n24392 & ~new_n25768 ;
  assign new_n25770 = ~new_n25766 & ~new_n25769 ;
  assign new_n25771 = ~new_n24936 & ~new_n25770 ;
  assign new_n25772 = new_n24768 & new_n25770 ;
  assign new_n25773 = ~new_n24934 & new_n25772 ;
  assign new_n25774 = ~new_n25771 & ~new_n25773 ;
  assign new_n25775 = ~new_n23175 & ~new_n25774 ;
  assign new_n25776 = ~new_n22680 & new_n23175 ;
  assign new_n25777 = ~new_n25775 & ~new_n25776 ;
  assign new_n25778 = ~new_n23177 & ~new_n25777 ;
  assign new_n25779 = ~new_n25763 & ~new_n25778 ;
  assign new_n25780 = lo1359 & ~new_n17706 ;
  assign new_n25781 = lo0955 & ~new_n14260 ;
  assign new_n25782 = ~lo0955 & new_n4807 ;
  assign new_n25783 = ~new_n25781 & ~new_n25782 ;
  assign new_n25784 = new_n17706 & ~new_n25783 ;
  assign new_n25785 = ~new_n25780 & ~new_n25784 ;
  assign new_n25786 = lo1360 & ~new_n17706 ;
  assign new_n25787 = lo0955 & ~new_n10308 ;
  assign new_n25788 = ~lo0955 & new_n2586 ;
  assign new_n25789 = ~new_n25787 & ~new_n25788 ;
  assign new_n25790 = new_n17706 & ~new_n25789 ;
  assign new_n25791 = ~new_n25786 & ~new_n25790 ;
  assign new_n25792 = lo1361 & new_n23177 ;
  assign new_n25793 = ~lo1361 & new_n23187 ;
  assign new_n25794 = lo1361 & ~new_n23187 ;
  assign new_n25795 = ~new_n25793 & ~new_n25794 ;
  assign new_n25796 = ~new_n24936 & ~new_n25795 ;
  assign new_n25797 = new_n24768 & new_n25795 ;
  assign new_n25798 = ~new_n24934 & new_n25797 ;
  assign new_n25799 = ~new_n25796 & ~new_n25798 ;
  assign new_n25800 = ~new_n23175 & ~new_n25799 ;
  assign new_n25801 = ~new_n22112 & new_n23175 ;
  assign new_n25802 = ~new_n25800 & ~new_n25801 ;
  assign new_n25803 = ~new_n23177 & ~new_n25802 ;
  assign new_n25804 = ~new_n25792 & ~new_n25803 ;
  assign new_n25805 = ~new_n22127 & new_n24961 ;
  assign new_n25806 = lo1408 & new_n24026 ;
  assign new_n25807 = ~new_n24027 & ~new_n25806 ;
  assign new_n25808 = new_n24026 & new_n25807 ;
  assign new_n25809 = ~new_n24910 & new_n25808 ;
  assign new_n25810 = ~new_n24754 & ~new_n25807 ;
  assign new_n25811 = ~new_n24928 & new_n25810 ;
  assign new_n25812 = ~new_n25809 & ~new_n25811 ;
  assign new_n25813 = ~new_n21027 & ~new_n25812 ;
  assign new_n25814 = ~new_n24754 & new_n25807 ;
  assign new_n25815 = new_n24928 & ~new_n25814 ;
  assign new_n25816 = ~new_n21027 & ~new_n25808 ;
  assign new_n25817 = ~new_n25815 & new_n25816 ;
  assign new_n25818 = new_n24355 & new_n24559 ;
  assign new_n25819 = ~new_n24563 & ~new_n25818 ;
  assign new_n25820 = new_n24345 & ~new_n25819 ;
  assign new_n25821 = ~new_n24355 & new_n24559 ;
  assign new_n25822 = ~new_n24560 & ~new_n25821 ;
  assign new_n25823 = ~new_n24345 & ~new_n25822 ;
  assign new_n25824 = ~new_n25820 & ~new_n25823 ;
  assign new_n25825 = ~new_n25817 & ~new_n25824 ;
  assign new_n25826 = ~new_n25813 & ~new_n25825 ;
  assign new_n25827 = new_n24960 & ~new_n25826 ;
  assign new_n25828 = ~new_n24365 & new_n24776 ;
  assign new_n25829 = new_n24365 & new_n24979 ;
  assign new_n25830 = ~new_n25828 & ~new_n25829 ;
  assign new_n25831 = lo0941 & ~new_n25830 ;
  assign new_n25832 = lo1362 & ~new_n24960 ;
  assign new_n25833 = ~new_n25831 & ~new_n25832 ;
  assign new_n25834 = ~new_n25827 & new_n25833 ;
  assign new_n25835 = ~new_n24959 & ~new_n24961 ;
  assign new_n25836 = ~new_n25834 & new_n25835 ;
  assign new_n25837 = ~new_n25805 & ~new_n25836 ;
  assign new_n25838 = lo1363 & ~new_n23161 ;
  assign new_n25839 = lo0931 & ~new_n2586 ;
  assign new_n25840 = ~new_n2586 & ~new_n25839 ;
  assign new_n25841 = ~new_n10308 & ~new_n25840 ;
  assign new_n25842 = ~lo0931 & new_n2586 ;
  assign new_n25843 = new_n10308 & new_n25842 ;
  assign new_n25844 = ~new_n25841 & ~new_n25843 ;
  assign new_n25845 = ~lo0932 & ~new_n25844 ;
  assign new_n25846 = lo0759 & lo0932 ;
  assign new_n25847 = ~new_n25845 & ~new_n25846 ;
  assign new_n25848 = new_n23161 & ~new_n25847 ;
  assign new_n25849 = ~new_n25838 & ~new_n25848 ;
  assign new_n25850 = lo1364 & new_n24963 ;
  assign new_n25851 = ~new_n24894 & ~new_n25126 ;
  assign new_n25852 = new_n24894 & new_n25124 ;
  assign new_n25853 = ~new_n24989 & new_n25852 ;
  assign new_n25854 = ~new_n25851 & ~new_n25853 ;
  assign new_n25855 = ~new_n24961 & ~new_n25854 ;
  assign new_n25856 = ~new_n22073 & new_n24961 ;
  assign new_n25857 = ~new_n25855 & ~new_n25856 ;
  assign new_n25858 = ~new_n24963 & ~new_n25857 ;
  assign new_n25859 = ~new_n25850 & ~new_n25858 ;
  assign new_n25860 = lo1365 & ~new_n23161 ;
  assign new_n25861 = lo0931 & ~new_n5549 ;
  assign new_n25862 = ~new_n5549 & ~new_n25861 ;
  assign new_n25863 = ~new_n14036 & ~new_n25862 ;
  assign new_n25864 = ~lo0931 & new_n5549 ;
  assign new_n25865 = new_n14036 & new_n25864 ;
  assign new_n25866 = ~new_n25863 & ~new_n25865 ;
  assign new_n25867 = ~lo0932 & ~new_n25866 ;
  assign new_n25868 = lo0556 & lo0932 ;
  assign new_n25869 = ~new_n25867 & ~new_n25868 ;
  assign new_n25870 = new_n23161 & ~new_n25869 ;
  assign new_n25871 = ~new_n25860 & ~new_n25870 ;
  assign new_n25872 = lo1366 & new_n23177 ;
  assign new_n25873 = ~lo1366 & new_n24463 ;
  assign new_n25874 = ~new_n24467 & ~new_n25873 ;
  assign new_n25875 = ~new_n24410 & ~new_n25874 ;
  assign new_n25876 = lo1366 & new_n24463 ;
  assign new_n25877 = ~new_n24464 & ~new_n25876 ;
  assign new_n25878 = new_n24410 & ~new_n25877 ;
  assign new_n25879 = ~new_n25875 & ~new_n25878 ;
  assign new_n25880 = ~new_n24936 & ~new_n25879 ;
  assign new_n25881 = new_n24768 & new_n25879 ;
  assign new_n25882 = ~new_n24934 & new_n25881 ;
  assign new_n25883 = ~new_n25880 & ~new_n25882 ;
  assign new_n25884 = ~new_n23175 & ~new_n25883 ;
  assign new_n25885 = ~new_n22082 & new_n23175 ;
  assign new_n25886 = ~new_n25884 & ~new_n25885 ;
  assign new_n25887 = ~new_n23177 & ~new_n25886 ;
  assign new_n25888 = ~new_n25872 & ~new_n25887 ;
  assign new_n25889 = lo1367 & ~new_n17706 ;
  assign new_n25890 = lo0955 & ~new_n14446 ;
  assign new_n25891 = ~lo0955 & new_n5265 ;
  assign new_n25892 = ~new_n25890 & ~new_n25891 ;
  assign new_n25893 = new_n17706 & ~new_n25892 ;
  assign new_n25894 = ~new_n25889 & ~new_n25893 ;
  assign new_n25895 = lo1368 & new_n24963 ;
  assign new_n25896 = new_n24333 & new_n24571 ;
  assign new_n25897 = ~new_n24575 & ~new_n25896 ;
  assign new_n25898 = new_n24323 & ~new_n25897 ;
  assign new_n25899 = ~new_n24333 & new_n24571 ;
  assign new_n25900 = ~new_n24572 & ~new_n25899 ;
  assign new_n25901 = ~new_n24323 & ~new_n25900 ;
  assign new_n25902 = ~new_n25898 & ~new_n25901 ;
  assign new_n25903 = ~new_n24991 & ~new_n25902 ;
  assign new_n25904 = new_n24978 & new_n25902 ;
  assign new_n25905 = ~new_n24989 & new_n25904 ;
  assign new_n25906 = ~new_n25903 & ~new_n25905 ;
  assign new_n25907 = ~new_n24961 & ~new_n25906 ;
  assign new_n25908 = ~new_n22260 & new_n24961 ;
  assign new_n25909 = ~new_n25907 & ~new_n25908 ;
  assign new_n25910 = ~new_n24963 & ~new_n25909 ;
  assign new_n25911 = ~new_n25895 & ~new_n25910 ;
  assign new_n25912 = lo1369 & ~new_n23161 ;
  assign new_n25913 = lo0931 & ~new_n6899 ;
  assign new_n25914 = ~new_n6899 & ~new_n25913 ;
  assign new_n25915 = ~new_n19223 & ~new_n25914 ;
  assign new_n25916 = ~lo0931 & new_n6899 ;
  assign new_n25917 = new_n19223 & new_n25916 ;
  assign new_n25918 = ~new_n25915 & ~new_n25917 ;
  assign new_n25919 = ~lo0932 & ~new_n25918 ;
  assign new_n25920 = lo0642 & lo0932 ;
  assign new_n25921 = ~new_n25919 & ~new_n25920 ;
  assign new_n25922 = new_n23161 & ~new_n25921 ;
  assign new_n25923 = ~new_n25912 & ~new_n25922 ;
  assign new_n25924 = lo1370 & new_n23177 ;
  assign new_n25925 = ~lo1370 & new_n23194 ;
  assign new_n25926 = ~new_n23198 & ~new_n25925 ;
  assign new_n25927 = new_n23185 & ~new_n25926 ;
  assign new_n25928 = lo1370 & new_n23194 ;
  assign new_n25929 = ~new_n23195 & ~new_n25928 ;
  assign new_n25930 = ~new_n23185 & ~new_n25929 ;
  assign new_n25931 = ~new_n25927 & ~new_n25930 ;
  assign new_n25932 = ~new_n24936 & ~new_n25931 ;
  assign new_n25933 = new_n24768 & new_n25931 ;
  assign new_n25934 = ~new_n24934 & new_n25933 ;
  assign new_n25935 = ~new_n25932 & ~new_n25934 ;
  assign new_n25936 = ~new_n23175 & ~new_n25935 ;
  assign new_n25937 = ~new_n22599 & new_n23175 ;
  assign new_n25938 = ~new_n25936 & ~new_n25937 ;
  assign new_n25939 = ~new_n23177 & ~new_n25938 ;
  assign new_n25940 = ~new_n25924 & ~new_n25939 ;
  assign new_n25941 = lo1371 & new_n24963 ;
  assign new_n25942 = ~new_n24873 & ~new_n25126 ;
  assign new_n25943 = new_n24873 & new_n25124 ;
  assign new_n25944 = ~new_n24989 & new_n25943 ;
  assign new_n25945 = ~new_n25942 & ~new_n25944 ;
  assign new_n25946 = ~new_n24961 & ~new_n25945 ;
  assign new_n25947 = ~new_n22428 & new_n24961 ;
  assign new_n25948 = ~new_n25946 & ~new_n25947 ;
  assign new_n25949 = ~new_n24963 & ~new_n25948 ;
  assign new_n25950 = ~new_n25941 & ~new_n25949 ;
  assign new_n25951 = lo1372 & ~new_n23161 ;
  assign new_n25952 = lo0931 & ~new_n4981 ;
  assign new_n25953 = ~new_n4981 & ~new_n25952 ;
  assign new_n25954 = ~new_n14419 & ~new_n25953 ;
  assign new_n25955 = ~lo0931 & new_n4981 ;
  assign new_n25956 = new_n14419 & new_n25955 ;
  assign new_n25957 = ~new_n25954 & ~new_n25956 ;
  assign new_n25958 = ~lo0932 & ~new_n25957 ;
  assign new_n25959 = lo0339 & lo0932 ;
  assign new_n25960 = ~new_n25958 & ~new_n25959 ;
  assign new_n25961 = new_n23161 & ~new_n25960 ;
  assign new_n25962 = ~new_n25951 & ~new_n25961 ;
  assign new_n25963 = lo1373 & new_n23177 ;
  assign new_n25964 = ~lo1373 & new_n24475 ;
  assign new_n25965 = ~new_n24479 & ~new_n25964 ;
  assign new_n25966 = ~new_n24404 & ~new_n25965 ;
  assign new_n25967 = lo1373 & new_n24475 ;
  assign new_n25968 = ~new_n24476 & ~new_n25967 ;
  assign new_n25969 = new_n24404 & ~new_n25968 ;
  assign new_n25970 = ~new_n25966 & ~new_n25969 ;
  assign new_n25971 = ~new_n24936 & ~new_n25970 ;
  assign new_n25972 = new_n24768 & new_n25970 ;
  assign new_n25973 = ~new_n24934 & new_n25972 ;
  assign new_n25974 = ~new_n25971 & ~new_n25973 ;
  assign new_n25975 = ~new_n23175 & ~new_n25974 ;
  assign new_n25976 = ~new_n22608 & new_n23175 ;
  assign new_n25977 = ~new_n25975 & ~new_n25976 ;
  assign new_n25978 = ~new_n23177 & ~new_n25977 ;
  assign new_n25979 = ~new_n25963 & ~new_n25978 ;
  assign new_n25980 = lo1374 & new_n24963 ;
  assign new_n25981 = new_n24322 & new_n24577 ;
  assign new_n25982 = ~new_n24581 & ~new_n25981 ;
  assign new_n25983 = new_n24312 & ~new_n25982 ;
  assign new_n25984 = ~new_n24322 & new_n24577 ;
  assign new_n25985 = ~new_n24578 & ~new_n25984 ;
  assign new_n25986 = ~new_n24312 & ~new_n25985 ;
  assign new_n25987 = ~new_n25983 & ~new_n25986 ;
  assign new_n25988 = ~new_n24991 & ~new_n25987 ;
  assign new_n25989 = new_n24978 & new_n25987 ;
  assign new_n25990 = ~new_n24989 & new_n25989 ;
  assign new_n25991 = ~new_n25988 & ~new_n25990 ;
  assign new_n25992 = ~new_n24961 & ~new_n25991 ;
  assign new_n25993 = ~new_n22272 & new_n24961 ;
  assign new_n25994 = ~new_n25992 & ~new_n25993 ;
  assign new_n25995 = ~new_n24963 & ~new_n25994 ;
  assign new_n25996 = ~new_n25980 & ~new_n25995 ;
  assign new_n25997 = lo1375 & ~new_n23161 ;
  assign new_n25998 = lo0931 & ~new_n6667 ;
  assign new_n25999 = ~new_n6667 & ~new_n25998 ;
  assign new_n26000 = ~new_n18863 & ~new_n25999 ;
  assign new_n26001 = ~lo0931 & new_n6667 ;
  assign new_n26002 = new_n18863 & new_n26001 ;
  assign new_n26003 = ~new_n26000 & ~new_n26002 ;
  assign new_n26004 = ~lo0932 & ~new_n26003 ;
  assign new_n26005 = lo0580 & lo0932 ;
  assign new_n26006 = ~new_n26004 & ~new_n26005 ;
  assign new_n26007 = new_n23161 & ~new_n26006 ;
  assign new_n26008 = ~new_n25997 & ~new_n26007 ;
  assign new_n26009 = lo1376 & new_n23177 ;
  assign new_n26010 = ~lo1376 & new_n23200 ;
  assign new_n26011 = ~new_n23204 & ~new_n26010 ;
  assign new_n26012 = new_n23184 & ~new_n26011 ;
  assign new_n26013 = lo1376 & new_n23200 ;
  assign new_n26014 = ~new_n23201 & ~new_n26013 ;
  assign new_n26015 = ~new_n23184 & ~new_n26014 ;
  assign new_n26016 = ~new_n26012 & ~new_n26015 ;
  assign new_n26017 = ~new_n24936 & ~new_n26016 ;
  assign new_n26018 = new_n24768 & new_n26016 ;
  assign new_n26019 = ~new_n24934 & new_n26018 ;
  assign new_n26020 = ~new_n26017 & ~new_n26019 ;
  assign new_n26021 = ~new_n23175 & ~new_n26020 ;
  assign new_n26022 = ~new_n22617 & new_n23175 ;
  assign new_n26023 = ~new_n26021 & ~new_n26022 ;
  assign new_n26024 = ~new_n23177 & ~new_n26023 ;
  assign new_n26025 = ~new_n26009 & ~new_n26024 ;
  assign new_n26026 = lo1377 & new_n24963 ;
  assign new_n26027 = ~new_n24866 & ~new_n25126 ;
  assign new_n26028 = new_n24866 & new_n25124 ;
  assign new_n26029 = ~new_n24989 & new_n26028 ;
  assign new_n26030 = ~new_n26027 & ~new_n26029 ;
  assign new_n26031 = ~new_n24961 & ~new_n26030 ;
  assign new_n26032 = ~new_n22440 & new_n24961 ;
  assign new_n26033 = ~new_n26031 & ~new_n26032 ;
  assign new_n26034 = ~new_n24963 & ~new_n26033 ;
  assign new_n26035 = ~new_n26026 & ~new_n26034 ;
  assign new_n26036 = lo1378 & ~new_n23161 ;
  assign new_n26037 = lo0931 & ~new_n4619 ;
  assign new_n26038 = ~new_n4619 & ~new_n26037 ;
  assign new_n26039 = ~new_n14393 & ~new_n26038 ;
  assign new_n26040 = ~lo0931 & new_n4619 ;
  assign new_n26041 = new_n14393 & new_n26040 ;
  assign new_n26042 = ~new_n26039 & ~new_n26041 ;
  assign new_n26043 = ~lo0932 & ~new_n26042 ;
  assign new_n26044 = lo0318 & lo0932 ;
  assign new_n26045 = ~new_n26043 & ~new_n26044 ;
  assign new_n26046 = new_n23161 & ~new_n26045 ;
  assign new_n26047 = ~new_n26036 & ~new_n26046 ;
  assign new_n26048 = lo1379 & new_n23177 ;
  assign new_n26049 = ~lo1379 & new_n24481 ;
  assign new_n26050 = ~new_n24485 & ~new_n26049 ;
  assign new_n26051 = ~new_n24401 & ~new_n26050 ;
  assign new_n26052 = lo1379 & new_n24481 ;
  assign new_n26053 = ~new_n24482 & ~new_n26052 ;
  assign new_n26054 = new_n24401 & ~new_n26053 ;
  assign new_n26055 = ~new_n26051 & ~new_n26054 ;
  assign new_n26056 = ~new_n24936 & ~new_n26055 ;
  assign new_n26057 = new_n24768 & new_n26055 ;
  assign new_n26058 = ~new_n24934 & new_n26057 ;
  assign new_n26059 = ~new_n26056 & ~new_n26058 ;
  assign new_n26060 = ~new_n23175 & ~new_n26059 ;
  assign new_n26061 = ~new_n22626 & new_n23175 ;
  assign new_n26062 = ~new_n26060 & ~new_n26061 ;
  assign new_n26063 = ~new_n23177 & ~new_n26062 ;
  assign new_n26064 = ~new_n26048 & ~new_n26063 ;
  assign new_n26065 = lo1380 & ~new_n17706 ;
  assign new_n26066 = lo0955 & ~new_n13907 ;
  assign new_n26067 = ~lo0955 & new_n7122 ;
  assign new_n26068 = ~new_n26066 & ~new_n26067 ;
  assign new_n26069 = new_n17706 & ~new_n26068 ;
  assign new_n26070 = ~new_n26065 & ~new_n26069 ;
  assign new_n26071 = lo1381 & ~new_n17706 ;
  assign new_n26072 = lo0955 & ~new_n13977 ;
  assign new_n26073 = ~lo0955 & ~new_n5170 ;
  assign new_n26074 = ~new_n26072 & ~new_n26073 ;
  assign new_n26075 = new_n17706 & ~new_n26074 ;
  assign new_n26076 = ~new_n26071 & ~new_n26075 ;
  assign new_n26077 = lo1382 & new_n23177 ;
  assign new_n26078 = ~lo1382 & ~new_n23188 ;
  assign new_n26079 = ~new_n23192 & ~new_n26078 ;
  assign new_n26080 = new_n23186 & ~new_n26079 ;
  assign new_n26081 = lo1382 & ~new_n23188 ;
  assign new_n26082 = ~new_n23189 & ~new_n26081 ;
  assign new_n26083 = ~new_n23186 & ~new_n26082 ;
  assign new_n26084 = ~new_n26080 & ~new_n26083 ;
  assign new_n26085 = ~new_n24936 & ~new_n26084 ;
  assign new_n26086 = new_n24768 & new_n26084 ;
  assign new_n26087 = ~new_n24934 & new_n26086 ;
  assign new_n26088 = ~new_n26085 & ~new_n26087 ;
  assign new_n26089 = ~new_n23175 & ~new_n26088 ;
  assign new_n26090 = ~new_n22581 & new_n23175 ;
  assign new_n26091 = ~new_n26089 & ~new_n26090 ;
  assign new_n26092 = ~new_n23177 & ~new_n26091 ;
  assign new_n26093 = ~new_n26077 & ~new_n26092 ;
  assign new_n26094 = lo1383 & new_n24963 ;
  assign new_n26095 = new_n24344 & new_n24565 ;
  assign new_n26096 = ~new_n24569 & ~new_n26095 ;
  assign new_n26097 = new_n24334 & ~new_n26096 ;
  assign new_n26098 = ~new_n24344 & new_n24565 ;
  assign new_n26099 = ~new_n24566 & ~new_n26098 ;
  assign new_n26100 = ~new_n24334 & ~new_n26099 ;
  assign new_n26101 = ~new_n26097 & ~new_n26100 ;
  assign new_n26102 = ~new_n24991 & ~new_n26101 ;
  assign new_n26103 = new_n24978 & new_n26101 ;
  assign new_n26104 = ~new_n24989 & new_n26103 ;
  assign new_n26105 = ~new_n26102 & ~new_n26104 ;
  assign new_n26106 = ~new_n24961 & ~new_n26105 ;
  assign new_n26107 = ~new_n22248 & new_n24961 ;
  assign new_n26108 = ~new_n26106 & ~new_n26107 ;
  assign new_n26109 = ~new_n24963 & ~new_n26108 ;
  assign new_n26110 = ~new_n26094 & ~new_n26109 ;
  assign new_n26111 = lo1384 & ~new_n15376 ;
  assign new_n26112 = lo0858 & ~lo1384 ;
  assign new_n26113 = ~lo1384 & ~new_n26112 ;
  assign new_n26114 = new_n7122 & ~new_n26113 ;
  assign new_n26115 = ~lo0858 & lo1384 ;
  assign new_n26116 = ~new_n7122 & new_n26115 ;
  assign new_n26117 = ~new_n26114 & ~new_n26116 ;
  assign new_n26118 = ~lo0859 & ~new_n26117 ;
  assign new_n26119 = lo0859 & ~new_n13907 ;
  assign new_n26120 = ~new_n26118 & ~new_n26119 ;
  assign new_n26121 = new_n15376 & ~new_n26120 ;
  assign new_n26122 = ~new_n26111 & ~new_n26121 ;
  assign new_n26123 = lo1385 & ~new_n23161 ;
  assign new_n26124 = lo0931 & ~new_n7122 ;
  assign new_n26125 = ~new_n7122 & ~new_n26124 ;
  assign new_n26126 = ~new_n13907 & ~new_n26125 ;
  assign new_n26127 = ~lo0931 & new_n7122 ;
  assign new_n26128 = new_n13907 & new_n26127 ;
  assign new_n26129 = ~new_n26126 & ~new_n26128 ;
  assign new_n26130 = ~lo0932 & ~new_n26129 ;
  assign new_n26131 = lo0803 & lo0932 ;
  assign new_n26132 = ~new_n26130 & ~new_n26131 ;
  assign new_n26133 = new_n23161 & ~new_n26132 ;
  assign new_n26134 = ~new_n26123 & ~new_n26133 ;
  assign new_n26135 = lo1386 & new_n23177 ;
  assign new_n26136 = ~lo1386 & new_n24421 ;
  assign new_n26137 = ~new_n24425 & ~new_n26136 ;
  assign new_n26138 = new_n24417 & ~new_n26137 ;
  assign new_n26139 = lo1386 & new_n24421 ;
  assign new_n26140 = ~new_n24422 & ~new_n26139 ;
  assign new_n26141 = ~new_n24417 & ~new_n26140 ;
  assign new_n26142 = ~new_n26138 & ~new_n26141 ;
  assign new_n26143 = ~new_n24936 & ~new_n26142 ;
  assign new_n26144 = new_n24768 & new_n26142 ;
  assign new_n26145 = ~new_n24934 & new_n26144 ;
  assign new_n26146 = ~new_n26143 & ~new_n26145 ;
  assign new_n26147 = ~new_n23175 & ~new_n26146 ;
  assign new_n26148 = ~new_n22725 & new_n23175 ;
  assign new_n26149 = ~new_n26147 & ~new_n26148 ;
  assign new_n26150 = ~new_n23177 & ~new_n26149 ;
  assign new_n26151 = ~new_n26135 & ~new_n26150 ;
  assign new_n26152 = lo1387 & new_n24963 ;
  assign new_n26153 = new_n24256 & new_n24613 ;
  assign new_n26154 = ~new_n24617 & ~new_n26153 ;
  assign new_n26155 = new_n24246 & ~new_n26154 ;
  assign new_n26156 = ~new_n24256 & new_n24613 ;
  assign new_n26157 = ~new_n24614 & ~new_n26156 ;
  assign new_n26158 = ~new_n24246 & ~new_n26157 ;
  assign new_n26159 = ~new_n26155 & ~new_n26158 ;
  assign new_n26160 = ~new_n24991 & ~new_n26159 ;
  assign new_n26161 = new_n24978 & new_n26159 ;
  assign new_n26162 = ~new_n24989 & new_n26161 ;
  assign new_n26163 = ~new_n26160 & ~new_n26162 ;
  assign new_n26164 = ~new_n24961 & ~new_n26163 ;
  assign new_n26165 = ~new_n22344 & new_n24961 ;
  assign new_n26166 = ~new_n26164 & ~new_n26165 ;
  assign new_n26167 = ~new_n24963 & ~new_n26166 ;
  assign new_n26168 = ~new_n26152 & ~new_n26167 ;
  assign new_n26169 = lo1388 & ~new_n23161 ;
  assign new_n26170 = lo0931 & new_n5170 ;
  assign new_n26171 = new_n5170 & ~new_n26170 ;
  assign new_n26172 = ~new_n13977 & ~new_n26171 ;
  assign new_n26173 = ~lo0931 & ~new_n5170 ;
  assign new_n26174 = new_n13977 & new_n26173 ;
  assign new_n26175 = ~new_n26172 & ~new_n26174 ;
  assign new_n26176 = ~lo0932 & ~new_n26175 ;
  assign new_n26177 = lo0825 & lo0932 ;
  assign new_n26178 = ~new_n26176 & ~new_n26177 ;
  assign new_n26179 = new_n23161 & ~new_n26178 ;
  assign new_n26180 = ~new_n26169 & ~new_n26179 ;
  assign new_n26181 = lo1389 & new_n24963 ;
  assign new_n26182 = ~new_n24880 & ~new_n25126 ;
  assign new_n26183 = new_n24880 & new_n25124 ;
  assign new_n26184 = ~new_n24989 & new_n26183 ;
  assign new_n26185 = ~new_n26182 & ~new_n26184 ;
  assign new_n26186 = ~new_n24961 & ~new_n26185 ;
  assign new_n26187 = ~new_n22416 & new_n24961 ;
  assign new_n26188 = ~new_n26186 & ~new_n26187 ;
  assign new_n26189 = ~new_n24963 & ~new_n26188 ;
  assign new_n26190 = ~new_n26181 & ~new_n26189 ;
  assign new_n26191 = lo1390 & ~new_n23161 ;
  assign new_n26192 = lo0931 & ~new_n5265 ;
  assign new_n26193 = ~new_n5265 & ~new_n26192 ;
  assign new_n26194 = ~new_n14446 & ~new_n26193 ;
  assign new_n26195 = ~lo0931 & new_n5265 ;
  assign new_n26196 = new_n14446 & new_n26195 ;
  assign new_n26197 = ~new_n26194 & ~new_n26196 ;
  assign new_n26198 = ~lo0932 & ~new_n26197 ;
  assign new_n26199 = lo0781 & lo0932 ;
  assign new_n26200 = ~new_n26198 & ~new_n26199 ;
  assign new_n26201 = new_n23161 & ~new_n26200 ;
  assign new_n26202 = ~new_n26191 & ~new_n26201 ;
  assign new_n26203 = lo1391 & new_n23177 ;
  assign new_n26204 = ~lo1391 & new_n24469 ;
  assign new_n26205 = ~new_n24473 & ~new_n26204 ;
  assign new_n26206 = ~new_n24407 & ~new_n26205 ;
  assign new_n26207 = lo1391 & new_n24469 ;
  assign new_n26208 = ~new_n24470 & ~new_n26207 ;
  assign new_n26209 = new_n24407 & ~new_n26208 ;
  assign new_n26210 = ~new_n26206 & ~new_n26209 ;
  assign new_n26211 = ~new_n24936 & ~new_n26210 ;
  assign new_n26212 = new_n24768 & new_n26210 ;
  assign new_n26213 = ~new_n24934 & new_n26212 ;
  assign new_n26214 = ~new_n26211 & ~new_n26213 ;
  assign new_n26215 = ~new_n23175 & ~new_n26214 ;
  assign new_n26216 = ~new_n22590 & new_n23175 ;
  assign new_n26217 = ~new_n26215 & ~new_n26216 ;
  assign new_n26218 = ~new_n23177 & ~new_n26217 ;
  assign new_n26219 = ~new_n26203 & ~new_n26218 ;
  assign new_n26220 = lo1392 & ~new_n17706 ;
  assign new_n26221 = lo0955 & ~new_n14234 ;
  assign new_n26222 = ~lo0955 & new_n4530 ;
  assign new_n26223 = ~new_n26221 & ~new_n26222 ;
  assign new_n26224 = new_n17706 & ~new_n26223 ;
  assign new_n26225 = ~new_n26220 & ~new_n26224 ;
  assign new_n26226 = lo1393 & new_n24963 ;
  assign new_n26227 = ~new_n24838 & ~new_n25126 ;
  assign new_n26228 = new_n24838 & new_n25124 ;
  assign new_n26229 = ~new_n24989 & new_n26228 ;
  assign new_n26230 = ~new_n26227 & ~new_n26229 ;
  assign new_n26231 = ~new_n24961 & ~new_n26230 ;
  assign new_n26232 = ~new_n22488 & new_n24961 ;
  assign new_n26233 = ~new_n26231 & ~new_n26232 ;
  assign new_n26234 = ~new_n24963 & ~new_n26233 ;
  assign new_n26235 = ~new_n26226 & ~new_n26234 ;
  assign new_n26236 = lo1394 & ~new_n23161 ;
  assign new_n26237 = lo0931 & ~new_n2813 ;
  assign new_n26238 = ~new_n2813 & ~new_n26237 ;
  assign new_n26239 = ~new_n14287 & ~new_n26238 ;
  assign new_n26240 = ~lo0931 & new_n2813 ;
  assign new_n26241 = new_n14287 & new_n26240 ;
  assign new_n26242 = ~new_n26239 & ~new_n26241 ;
  assign new_n26243 = ~lo0932 & ~new_n26242 ;
  assign new_n26244 = lo0619 & lo0932 ;
  assign new_n26245 = ~new_n26243 & ~new_n26244 ;
  assign new_n26246 = new_n23161 & ~new_n26245 ;
  assign new_n26247 = ~new_n26236 & ~new_n26246 ;
  assign new_n26248 = lo1395 & new_n23177 ;
  assign new_n26249 = ~lo1395 & new_n24505 ;
  assign new_n26250 = ~new_n24509 & ~new_n26249 ;
  assign new_n26251 = ~new_n24389 & ~new_n26250 ;
  assign new_n26252 = lo1395 & new_n24505 ;
  assign new_n26253 = ~new_n24506 & ~new_n26252 ;
  assign new_n26254 = new_n24389 & ~new_n26253 ;
  assign new_n26255 = ~new_n26251 & ~new_n26254 ;
  assign new_n26256 = ~new_n24936 & ~new_n26255 ;
  assign new_n26257 = new_n24768 & new_n26255 ;
  assign new_n26258 = ~new_n24934 & new_n26257 ;
  assign new_n26259 = ~new_n26256 & ~new_n26258 ;
  assign new_n26260 = ~new_n23175 & ~new_n26259 ;
  assign new_n26261 = ~new_n22698 & new_n23175 ;
  assign new_n26262 = ~new_n26260 & ~new_n26261 ;
  assign new_n26263 = ~new_n23177 & ~new_n26262 ;
  assign new_n26264 = ~new_n26248 & ~new_n26263 ;
  assign new_n26265 = lo1396 & new_n23177 ;
  assign new_n26266 = ~lo1396 & new_n24433 ;
  assign new_n26267 = ~new_n24437 & ~new_n26266 ;
  assign new_n26268 = new_n24415 & ~new_n26267 ;
  assign new_n26269 = lo1396 & new_n24433 ;
  assign new_n26270 = ~new_n24434 & ~new_n26269 ;
  assign new_n26271 = ~new_n24415 & ~new_n26270 ;
  assign new_n26272 = ~new_n26268 & ~new_n26271 ;
  assign new_n26273 = ~new_n24936 & ~new_n26272 ;
  assign new_n26274 = new_n24768 & new_n26272 ;
  assign new_n26275 = ~new_n24934 & new_n26274 ;
  assign new_n26276 = ~new_n26273 & ~new_n26275 ;
  assign new_n26277 = ~new_n23175 & ~new_n26276 ;
  assign new_n26278 = ~new_n22761 & new_n23175 ;
  assign new_n26279 = ~new_n26277 & ~new_n26278 ;
  assign new_n26280 = ~new_n23177 & ~new_n26279 ;
  assign new_n26281 = ~new_n26265 & ~new_n26280 ;
  assign new_n26282 = lo1397 & ~new_n23161 ;
  assign new_n26283 = lo0931 & new_n4446 ;
  assign new_n26284 = new_n4446 & ~new_n26283 ;
  assign new_n26285 = ~new_n14578 & ~new_n26284 ;
  assign new_n26286 = ~lo0931 & ~new_n4446 ;
  assign new_n26287 = new_n14578 & new_n26286 ;
  assign new_n26288 = ~new_n26285 & ~new_n26287 ;
  assign new_n26289 = ~lo0932 & ~new_n26288 ;
  assign new_n26290 = lo0720 & lo0932 ;
  assign new_n26291 = ~new_n26289 & ~new_n26290 ;
  assign new_n26292 = new_n23161 & ~new_n26291 ;
  assign new_n26293 = ~new_n26282 & ~new_n26292 ;
  assign new_n26294 = lo1398 & new_n24963 ;
  assign new_n26295 = new_n24234 & new_n24625 ;
  assign new_n26296 = ~new_n24629 & ~new_n26295 ;
  assign new_n26297 = new_n24224 & ~new_n26296 ;
  assign new_n26298 = ~new_n24234 & new_n24625 ;
  assign new_n26299 = ~new_n24626 & ~new_n26298 ;
  assign new_n26300 = ~new_n24224 & ~new_n26299 ;
  assign new_n26301 = ~new_n26297 & ~new_n26300 ;
  assign new_n26302 = ~new_n24991 & ~new_n26301 ;
  assign new_n26303 = new_n24978 & new_n26301 ;
  assign new_n26304 = ~new_n24989 & new_n26303 ;
  assign new_n26305 = ~new_n26302 & ~new_n26304 ;
  assign new_n26306 = ~new_n24961 & ~new_n26305 ;
  assign new_n26307 = ~new_n22368 & new_n24961 ;
  assign new_n26308 = ~new_n26306 & ~new_n26307 ;
  assign new_n26309 = ~new_n24963 & ~new_n26308 ;
  assign new_n26310 = ~new_n26294 & ~new_n26309 ;
  assign new_n26311 = lo1399 & new_n24963 ;
  assign new_n26312 = ~new_n24810 & ~new_n25126 ;
  assign new_n26313 = new_n24810 & new_n25124 ;
  assign new_n26314 = ~new_n24989 & new_n26313 ;
  assign new_n26315 = ~new_n26312 & ~new_n26314 ;
  assign new_n26316 = ~new_n24961 & ~new_n26315 ;
  assign new_n26317 = ~new_n22536 & new_n24961 ;
  assign new_n26318 = ~new_n26316 & ~new_n26317 ;
  assign new_n26319 = ~new_n24963 & ~new_n26318 ;
  assign new_n26320 = ~new_n26311 & ~new_n26319 ;
  assign new_n26321 = lo1400 & ~new_n23161 ;
  assign new_n26322 = lo0931 & ~new_n3806 ;
  assign new_n26323 = ~new_n3806 & ~new_n26322 ;
  assign new_n26324 = ~new_n14181 & ~new_n26323 ;
  assign new_n26325 = ~lo0931 & new_n3806 ;
  assign new_n26326 = new_n14181 & new_n26325 ;
  assign new_n26327 = ~new_n26324 & ~new_n26326 ;
  assign new_n26328 = ~lo0932 & ~new_n26327 ;
  assign new_n26329 = lo0661 & lo0932 ;
  assign new_n26330 = ~new_n26328 & ~new_n26329 ;
  assign new_n26331 = new_n23161 & ~new_n26330 ;
  assign new_n26332 = ~new_n26321 & ~new_n26331 ;
  assign new_n26333 = lo1401 & new_n23177 ;
  assign new_n26334 = ~lo1401 & new_n24529 ;
  assign new_n26335 = ~new_n24533 & ~new_n26334 ;
  assign new_n26336 = ~new_n24377 & ~new_n26335 ;
  assign new_n26337 = lo1401 & new_n24529 ;
  assign new_n26338 = ~new_n24530 & ~new_n26337 ;
  assign new_n26339 = new_n24377 & ~new_n26338 ;
  assign new_n26340 = ~new_n26336 & ~new_n26339 ;
  assign new_n26341 = ~new_n24936 & ~new_n26340 ;
  assign new_n26342 = new_n24768 & new_n26340 ;
  assign new_n26343 = ~new_n24934 & new_n26342 ;
  assign new_n26344 = ~new_n26341 & ~new_n26343 ;
  assign new_n26345 = ~new_n23175 & ~new_n26344 ;
  assign new_n26346 = ~new_n22770 & new_n23175 ;
  assign new_n26347 = ~new_n26345 & ~new_n26346 ;
  assign new_n26348 = ~new_n23177 & ~new_n26347 ;
  assign new_n26349 = ~new_n26333 & ~new_n26348 ;
  assign new_n26350 = lo1402 & new_n24963 ;
  assign new_n26351 = ~new_n24824 & ~new_n25126 ;
  assign new_n26352 = new_n24824 & new_n25124 ;
  assign new_n26353 = ~new_n24989 & new_n26352 ;
  assign new_n26354 = ~new_n26351 & ~new_n26353 ;
  assign new_n26355 = ~new_n24961 & ~new_n26354 ;
  assign new_n26356 = ~new_n22512 & new_n24961 ;
  assign new_n26357 = ~new_n26355 & ~new_n26356 ;
  assign new_n26358 = ~new_n24963 & ~new_n26357 ;
  assign new_n26359 = ~new_n26350 & ~new_n26358 ;
  assign new_n26360 = lo1403 & ~new_n23161 ;
  assign new_n26361 = lo0931 & ~new_n4530 ;
  assign new_n26362 = ~new_n4530 & ~new_n26361 ;
  assign new_n26363 = ~new_n14234 & ~new_n26362 ;
  assign new_n26364 = ~lo0931 & new_n4530 ;
  assign new_n26365 = new_n14234 & new_n26364 ;
  assign new_n26366 = ~new_n26363 & ~new_n26365 ;
  assign new_n26367 = ~lo0932 & ~new_n26366 ;
  assign new_n26368 = lo0843 & lo0932 ;
  assign new_n26369 = ~new_n26367 & ~new_n26368 ;
  assign new_n26370 = new_n23161 & ~new_n26369 ;
  assign new_n26371 = ~new_n26360 & ~new_n26370 ;
  assign new_n26372 = lo1404 & new_n23177 ;
  assign new_n26373 = ~lo1404 & new_n24517 ;
  assign new_n26374 = ~new_n24521 & ~new_n26373 ;
  assign new_n26375 = ~new_n24383 & ~new_n26374 ;
  assign new_n26376 = lo1404 & new_n24517 ;
  assign new_n26377 = ~new_n24518 & ~new_n26376 ;
  assign new_n26378 = new_n24383 & ~new_n26377 ;
  assign new_n26379 = ~new_n26375 & ~new_n26378 ;
  assign new_n26380 = ~new_n24936 & ~new_n26379 ;
  assign new_n26381 = new_n24768 & new_n26379 ;
  assign new_n26382 = ~new_n24934 & new_n26381 ;
  assign new_n26383 = ~new_n26380 & ~new_n26382 ;
  assign new_n26384 = ~new_n23175 & ~new_n26383 ;
  assign new_n26385 = ~new_n22734 & new_n23175 ;
  assign new_n26386 = ~new_n26384 & ~new_n26385 ;
  assign new_n26387 = ~new_n23177 & ~new_n26386 ;
  assign new_n26388 = ~new_n26372 & ~new_n26387 ;
  assign new_n26389 = lo1405 & new_n24963 ;
  assign new_n26390 = ~new_n24796 & ~new_n25126 ;
  assign new_n26391 = new_n24796 & new_n25124 ;
  assign new_n26392 = ~new_n24989 & new_n26391 ;
  assign new_n26393 = ~new_n26390 & ~new_n26392 ;
  assign new_n26394 = ~new_n24961 & ~new_n26393 ;
  assign new_n26395 = ~new_n22560 & new_n24961 ;
  assign new_n26396 = ~new_n26394 & ~new_n26395 ;
  assign new_n26397 = ~new_n24963 & ~new_n26396 ;
  assign new_n26398 = ~new_n26389 & ~new_n26397 ;
  assign new_n26399 = lo1406 & ~new_n23161 ;
  assign new_n26400 = lo0931 & ~new_n2990 ;
  assign new_n26401 = ~new_n2990 & ~new_n26400 ;
  assign new_n26402 = ~new_n14128 & ~new_n26401 ;
  assign new_n26403 = ~lo0931 & new_n2990 ;
  assign new_n26404 = new_n14128 & new_n26403 ;
  assign new_n26405 = ~new_n26402 & ~new_n26404 ;
  assign new_n26406 = ~lo0932 & ~new_n26405 ;
  assign new_n26407 = lo0457 & lo0932 ;
  assign new_n26408 = ~new_n26406 & ~new_n26407 ;
  assign new_n26409 = new_n23161 & ~new_n26408 ;
  assign new_n26410 = ~new_n26399 & ~new_n26409 ;
  assign new_n26411 = lo1407 & new_n23177 ;
  assign new_n26412 = ~lo1407 & new_n24541 ;
  assign new_n26413 = ~new_n24545 & ~new_n26412 ;
  assign new_n26414 = ~new_n24371 & ~new_n26413 ;
  assign new_n26415 = lo1407 & new_n24541 ;
  assign new_n26416 = ~new_n24542 & ~new_n26415 ;
  assign new_n26417 = new_n24371 & ~new_n26416 ;
  assign new_n26418 = ~new_n26414 & ~new_n26417 ;
  assign new_n26419 = ~new_n24936 & ~new_n26418 ;
  assign new_n26420 = new_n24768 & new_n26418 ;
  assign new_n26421 = ~new_n24934 & new_n26420 ;
  assign new_n26422 = ~new_n26419 & ~new_n26421 ;
  assign new_n26423 = ~new_n23175 & ~new_n26422 ;
  assign new_n26424 = ~new_n22806 & new_n23175 ;
  assign new_n26425 = ~new_n26423 & ~new_n26424 ;
  assign new_n26426 = ~new_n23177 & ~new_n26425 ;
  assign new_n26427 = ~new_n26411 & ~new_n26426 ;
  assign new_n26428 = ~new_n22043 & new_n24961 ;
  assign new_n26429 = new_n24960 & ~new_n25831 ;
  assign new_n26430 = ~new_n21027 & ~new_n24026 ;
  assign new_n26431 = new_n26429 & ~new_n26430 ;
  assign new_n26432 = ~new_n24754 & new_n26431 ;
  assign new_n26433 = lo1408 & ~new_n26432 ;
  assign new_n26434 = ~new_n21027 & new_n24026 ;
  assign new_n26435 = new_n26429 & ~new_n26434 ;
  assign new_n26436 = new_n24754 & new_n26435 ;
  assign new_n26437 = ~new_n26433 & ~new_n26436 ;
  assign new_n26438 = new_n25835 & ~new_n26437 ;
  assign new_n26439 = ~new_n26428 & ~new_n26438 ;
  assign new_n26440 = lo1409 & ~new_n23161 ;
  assign new_n26441 = lo0931 & ~new_n2718 ;
  assign new_n26442 = ~new_n2718 & ~new_n26441 ;
  assign new_n26443 = ~new_n14060 & ~new_n26442 ;
  assign new_n26444 = ~lo0931 & new_n2718 ;
  assign new_n26445 = new_n14060 & new_n26444 ;
  assign new_n26446 = ~new_n26443 & ~new_n26445 ;
  assign new_n26447 = ~lo0932 & ~new_n26446 ;
  assign new_n26448 = lo0476 & lo0932 ;
  assign new_n26449 = ~new_n26447 & ~new_n26448 ;
  assign new_n26450 = new_n23161 & ~new_n26449 ;
  assign new_n26451 = ~new_n26440 & ~new_n26450 ;
  assign new_n26452 = ~new_n22024 & new_n23175 ;
  assign new_n26453 = ~new_n24365 & ~new_n24775 ;
  assign new_n26454 = new_n24365 & new_n24775 ;
  assign new_n26455 = lo1410 & ~new_n26454 ;
  assign new_n26456 = ~new_n26453 & ~new_n26455 ;
  assign new_n26457 = lo0941 & ~new_n26456 ;
  assign new_n26458 = ~new_n24775 & ~new_n25817 ;
  assign new_n26459 = ~new_n25813 & ~new_n26458 ;
  assign new_n26460 = ~lo0941 & ~new_n26459 ;
  assign new_n26461 = ~new_n26457 & ~new_n26460 ;
  assign new_n26462 = lo0938 & ~new_n26461 ;
  assign new_n26463 = ~lo0938 & lo1410 ;
  assign new_n26464 = ~new_n26462 & ~new_n26463 ;
  assign new_n26465 = ~new_n23174 & ~new_n23175 ;
  assign new_n26466 = ~new_n26464 & new_n26465 ;
  assign new_n26467 = ~new_n26452 & ~new_n26466 ;
  assign new_n26468 = lo1411 & new_n23177 ;
  assign new_n26469 = ~lo1411 & new_n24427 ;
  assign new_n26470 = ~new_n24431 & ~new_n26469 ;
  assign new_n26471 = new_n24416 & ~new_n26470 ;
  assign new_n26472 = lo1411 & new_n24427 ;
  assign new_n26473 = ~new_n24428 & ~new_n26472 ;
  assign new_n26474 = ~new_n24416 & ~new_n26473 ;
  assign new_n26475 = ~new_n26471 & ~new_n26474 ;
  assign new_n26476 = ~new_n24936 & ~new_n26475 ;
  assign new_n26477 = new_n24768 & new_n26475 ;
  assign new_n26478 = ~new_n24934 & new_n26477 ;
  assign new_n26479 = ~new_n26476 & ~new_n26478 ;
  assign new_n26480 = ~new_n23175 & ~new_n26479 ;
  assign new_n26481 = ~new_n22743 & new_n23175 ;
  assign new_n26482 = ~new_n26480 & ~new_n26481 ;
  assign new_n26483 = ~new_n23177 & ~new_n26482 ;
  assign new_n26484 = ~new_n26468 & ~new_n26483 ;
  assign new_n26485 = lo1412 & ~new_n23161 ;
  assign new_n26486 = lo0931 & new_n4889 ;
  assign new_n26487 = new_n4889 & ~new_n26486 ;
  assign new_n26488 = ~new_n14525 & ~new_n26487 ;
  assign new_n26489 = ~lo0931 & ~new_n4889 ;
  assign new_n26490 = new_n14525 & new_n26489 ;
  assign new_n26491 = ~new_n26488 & ~new_n26490 ;
  assign new_n26492 = ~lo0932 & ~new_n26491 ;
  assign new_n26493 = lo0699 & lo0932 ;
  assign new_n26494 = ~new_n26492 & ~new_n26493 ;
  assign new_n26495 = new_n23161 & ~new_n26494 ;
  assign new_n26496 = ~new_n26485 & ~new_n26495 ;
  assign new_n26497 = lo1413 & new_n24963 ;
  assign new_n26498 = new_n24245 & new_n24619 ;
  assign new_n26499 = ~new_n24623 & ~new_n26498 ;
  assign new_n26500 = new_n24235 & ~new_n26499 ;
  assign new_n26501 = ~new_n24245 & new_n24619 ;
  assign new_n26502 = ~new_n24620 & ~new_n26501 ;
  assign new_n26503 = ~new_n24235 & ~new_n26502 ;
  assign new_n26504 = ~new_n26500 & ~new_n26503 ;
  assign new_n26505 = ~new_n24991 & ~new_n26504 ;
  assign new_n26506 = new_n24978 & new_n26504 ;
  assign new_n26507 = ~new_n24989 & new_n26506 ;
  assign new_n26508 = ~new_n26505 & ~new_n26507 ;
  assign new_n26509 = ~new_n24961 & ~new_n26508 ;
  assign new_n26510 = ~new_n22356 & new_n24961 ;
  assign new_n26511 = ~new_n26509 & ~new_n26510 ;
  assign new_n26512 = ~new_n24963 & ~new_n26511 ;
  assign new_n26513 = ~new_n26497 & ~new_n26512 ;
  assign new_n26514 = lo1414 & new_n24963 ;
  assign new_n26515 = ~new_n24817 & ~new_n25126 ;
  assign new_n26516 = new_n24817 & new_n25124 ;
  assign new_n26517 = ~new_n24989 & new_n26516 ;
  assign new_n26518 = ~new_n26515 & ~new_n26517 ;
  assign new_n26519 = ~new_n24961 & ~new_n26518 ;
  assign new_n26520 = ~new_n22524 & new_n24961 ;
  assign new_n26521 = ~new_n26519 & ~new_n26520 ;
  assign new_n26522 = ~new_n24963 & ~new_n26521 ;
  assign new_n26523 = ~new_n26514 & ~new_n26522 ;
  assign new_n26524 = lo1415 & ~new_n23161 ;
  assign new_n26525 = lo0931 & ~new_n4086 ;
  assign new_n26526 = ~new_n4086 & ~new_n26525 ;
  assign new_n26527 = ~new_n14207 & ~new_n26526 ;
  assign new_n26528 = ~lo0931 & new_n4086 ;
  assign new_n26529 = new_n14207 & new_n26528 ;
  assign new_n26530 = ~new_n26527 & ~new_n26529 ;
  assign new_n26531 = ~lo0932 & ~new_n26530 ;
  assign new_n26532 = lo0680 & lo0932 ;
  assign new_n26533 = ~new_n26531 & ~new_n26532 ;
  assign new_n26534 = new_n23161 & ~new_n26533 ;
  assign new_n26535 = ~new_n26524 & ~new_n26534 ;
  assign new_n26536 = lo1416 & new_n23177 ;
  assign new_n26537 = ~lo1416 & new_n24523 ;
  assign new_n26538 = ~new_n24527 & ~new_n26537 ;
  assign new_n26539 = ~new_n24380 & ~new_n26538 ;
  assign new_n26540 = lo1416 & new_n24523 ;
  assign new_n26541 = ~new_n24524 & ~new_n26540 ;
  assign new_n26542 = new_n24380 & ~new_n26541 ;
  assign new_n26543 = ~new_n26539 & ~new_n26542 ;
  assign new_n26544 = ~new_n24936 & ~new_n26543 ;
  assign new_n26545 = new_n24768 & new_n26543 ;
  assign new_n26546 = ~new_n24934 & new_n26545 ;
  assign new_n26547 = ~new_n26544 & ~new_n26546 ;
  assign new_n26548 = ~new_n23175 & ~new_n26547 ;
  assign new_n26549 = ~new_n22752 & new_n23175 ;
  assign new_n26550 = ~new_n26548 & ~new_n26549 ;
  assign new_n26551 = ~new_n23177 & ~new_n26550 ;
  assign new_n26552 = ~new_n26536 & ~new_n26551 ;
  assign new_n26553 = lo1417 & new_n24963 ;
  assign new_n26554 = ~new_n24831 & ~new_n25126 ;
  assign new_n26555 = new_n24831 & new_n25124 ;
  assign new_n26556 = ~new_n24989 & new_n26555 ;
  assign new_n26557 = ~new_n26554 & ~new_n26556 ;
  assign new_n26558 = ~new_n24961 & ~new_n26557 ;
  assign new_n26559 = ~new_n22500 & new_n24961 ;
  assign new_n26560 = ~new_n26558 & ~new_n26559 ;
  assign new_n26561 = ~new_n24963 & ~new_n26560 ;
  assign new_n26562 = ~new_n26553 & ~new_n26561 ;
  assign new_n26563 = lo1418 & ~new_n23161 ;
  assign new_n26564 = lo0931 & ~new_n4807 ;
  assign new_n26565 = ~new_n4807 & ~new_n26564 ;
  assign new_n26566 = ~new_n14260 & ~new_n26565 ;
  assign new_n26567 = ~lo0931 & new_n4807 ;
  assign new_n26568 = new_n14260 & new_n26567 ;
  assign new_n26569 = ~new_n26566 & ~new_n26568 ;
  assign new_n26570 = ~lo0932 & ~new_n26569 ;
  assign new_n26571 = lo0739 & lo0932 ;
  assign new_n26572 = ~new_n26570 & ~new_n26571 ;
  assign new_n26573 = new_n23161 & ~new_n26572 ;
  assign new_n26574 = ~new_n26563 & ~new_n26573 ;
  assign new_n26575 = lo1419 & new_n23177 ;
  assign new_n26576 = ~lo1419 & new_n24511 ;
  assign new_n26577 = ~new_n24515 & ~new_n26576 ;
  assign new_n26578 = ~new_n24386 & ~new_n26577 ;
  assign new_n26579 = lo1419 & new_n24511 ;
  assign new_n26580 = ~new_n24512 & ~new_n26579 ;
  assign new_n26581 = new_n24386 & ~new_n26580 ;
  assign new_n26582 = ~new_n26578 & ~new_n26581 ;
  assign new_n26583 = ~new_n24936 & ~new_n26582 ;
  assign new_n26584 = new_n24768 & new_n26582 ;
  assign new_n26585 = ~new_n24934 & new_n26584 ;
  assign new_n26586 = ~new_n26583 & ~new_n26585 ;
  assign new_n26587 = ~new_n23175 & ~new_n26586 ;
  assign new_n26588 = ~new_n22716 & new_n23175 ;
  assign new_n26589 = ~new_n26587 & ~new_n26588 ;
  assign new_n26590 = ~new_n23177 & ~new_n26589 ;
  assign new_n26591 = ~new_n26575 & ~new_n26590 ;
  assign new_n26592 = lo1420 & ~new_n21479 ;
  assign new_n26593 = lo1470 & ~new_n14601 ;
  assign new_n26594 = new_n14601 & ~new_n21514 ;
  assign new_n26595 = ~new_n26593 & ~new_n26594 ;
  assign new_n26596 = new_n21479 & ~new_n26595 ;
  assign new_n26597 = ~new_n26592 & ~new_n26596 ;
  assign new_n26598 = lo1421 & ~new_n21479 ;
  assign new_n26599 = lo1471 & ~new_n14601 ;
  assign new_n26600 = new_n14601 & ~new_n21537 ;
  assign new_n26601 = ~new_n26599 & ~new_n26600 ;
  assign new_n26602 = new_n21479 & ~new_n26601 ;
  assign new_n26603 = ~new_n26598 & ~new_n26602 ;
  assign new_n26604 = lo1422 & ~new_n21479 ;
  assign new_n26605 = lo1469 & ~new_n14601 ;
  assign new_n26606 = new_n14601 & ~new_n21491 ;
  assign new_n26607 = ~new_n26605 & ~new_n26606 ;
  assign new_n26608 = new_n21479 & ~new_n26607 ;
  assign new_n26609 = ~new_n26604 & ~new_n26608 ;
  assign new_n26610 = lo1423 & ~new_n21479 ;
  assign new_n26611 = lo1472 & ~new_n14601 ;
  assign new_n26612 = new_n14601 & ~new_n21560 ;
  assign new_n26613 = ~new_n26611 & ~new_n26612 ;
  assign new_n26614 = new_n21479 & ~new_n26613 ;
  assign new_n26615 = ~new_n26610 & ~new_n26614 ;
  assign new_n26616 = lo1424 & ~new_n21479 ;
  assign new_n26617 = lo1473 & ~new_n14601 ;
  assign new_n26618 = new_n14601 & ~new_n21671 ;
  assign new_n26619 = ~new_n26617 & ~new_n26618 ;
  assign new_n26620 = new_n21479 & ~new_n26619 ;
  assign new_n26621 = ~new_n26616 & ~new_n26620 ;
  assign new_n26622 = ~lo0017 & ~new_n14656 ;
  assign new_n26623 = ~lo1425 & new_n14652 ;
  assign new_n26624 = lo1425 & ~new_n14652 ;
  assign new_n26625 = ~new_n26623 & ~new_n26624 ;
  assign new_n26626 = new_n26622 & ~new_n26625 ;
  assign new_n26627 = lo0017 & ~new_n26622 ;
  assign new_n26628 = ~new_n26626 & ~new_n26627 ;
  assign new_n26629 = lo1425 & new_n14652 ;
  assign new_n26630 = lo1426 & ~new_n26629 ;
  assign new_n26631 = ~lo1426 & new_n26629 ;
  assign new_n26632 = ~new_n26630 & ~new_n26631 ;
  assign new_n26633 = new_n26622 & ~new_n26632 ;
  assign new_n26634 = lo1426 & new_n26629 ;
  assign new_n26635 = lo1427 & ~new_n26634 ;
  assign new_n26636 = ~lo1427 & new_n26634 ;
  assign new_n26637 = ~new_n26635 & ~new_n26636 ;
  assign new_n26638 = new_n26622 & ~new_n26637 ;
  assign new_n26639 = lo1427 & new_n26634 ;
  assign new_n26640 = lo1428 & ~new_n26639 ;
  assign new_n26641 = ~lo1428 & new_n26639 ;
  assign new_n26642 = ~new_n26640 & ~new_n26641 ;
  assign new_n26643 = new_n26622 & ~new_n26642 ;
  assign new_n26644 = ~new_n26627 & ~new_n26643 ;
  assign new_n26645 = lo1075 & lo1429 ;
  assign new_n26646 = ~lo1075 & ~lo1429 ;
  assign new_n26647 = ~new_n26645 & ~new_n26646 ;
  assign new_n26648 = lo1074 & ~new_n26647 ;
  assign new_n26649 = ~lo1074 & lo1429 ;
  assign new_n26650 = ~new_n26648 & ~new_n26649 ;
  assign new_n26651 = lo1430 & ~new_n26650 ;
  assign new_n26652 = lo1429 & ~lo1430 ;
  assign new_n26653 = ~new_n26651 & ~new_n26652 ;
  assign new_n26654 = ~lo0017 & ~new_n26653 ;
  assign new_n26655 = lo1075 & lo1430 ;
  assign new_n26656 = ~lo1075 & ~lo1430 ;
  assign new_n26657 = ~new_n26655 & ~new_n26656 ;
  assign new_n26658 = lo1074 & ~new_n26657 ;
  assign new_n26659 = ~lo1074 & lo1430 ;
  assign new_n26660 = ~new_n26658 & ~new_n26659 ;
  assign new_n26661 = ~lo0017 & ~new_n26660 ;
  assign new_n26662 = ~lo0984 & ~new_n16687 ;
  assign new_n26663 = lo1431 & new_n26662 ;
  assign new_n26664 = lo1441 & ~lo1443 ;
  assign new_n26665 = ~lo1441 & ~lo1443 ;
  assign new_n26666 = ~lo1441 & lo1443 ;
  assign new_n26667 = ~new_n26665 & ~new_n26666 ;
  assign new_n26668 = ~new_n26664 & new_n26667 ;
  assign new_n26669 = ~lo1439 & ~new_n26668 ;
  assign new_n26670 = ~lo1439 & new_n26668 ;
  assign new_n26671 = lo1439 & ~new_n26668 ;
  assign new_n26672 = ~new_n26670 & ~new_n26671 ;
  assign new_n26673 = ~new_n26669 & new_n26672 ;
  assign new_n26674 = ~lo1433 & ~new_n26673 ;
  assign new_n26675 = ~lo1433 & new_n26673 ;
  assign new_n26676 = lo1433 & ~new_n26673 ;
  assign new_n26677 = ~new_n26675 & ~new_n26676 ;
  assign new_n26678 = ~new_n26674 & new_n26677 ;
  assign new_n26679 = ~lo1442 & ~new_n26678 ;
  assign new_n26680 = ~lo1442 & new_n26678 ;
  assign new_n26681 = lo1442 & ~new_n26678 ;
  assign new_n26682 = ~new_n26680 & ~new_n26681 ;
  assign new_n26683 = ~new_n26679 & new_n26682 ;
  assign new_n26684 = ~lo1438 & ~new_n26683 ;
  assign new_n26685 = ~lo1438 & new_n26683 ;
  assign new_n26686 = lo1438 & ~new_n26683 ;
  assign new_n26687 = ~new_n26685 & ~new_n26686 ;
  assign new_n26688 = ~new_n26684 & new_n26687 ;
  assign new_n26689 = ~lo1440 & ~new_n26688 ;
  assign new_n26690 = ~lo1440 & new_n26688 ;
  assign new_n26691 = lo1440 & ~new_n26688 ;
  assign new_n26692 = ~new_n26690 & ~new_n26691 ;
  assign new_n26693 = ~new_n26689 & new_n26692 ;
  assign new_n26694 = ~lo1431 & new_n26693 ;
  assign new_n26695 = lo1431 & ~new_n26693 ;
  assign new_n26696 = ~new_n26694 & ~new_n26695 ;
  assign new_n26697 = ~new_n16687 & ~new_n26696 ;
  assign new_n26698 = ~lo1279 & new_n16687 ;
  assign new_n26699 = ~new_n26697 & ~new_n26698 ;
  assign new_n26700 = ~new_n26662 & ~new_n26699 ;
  assign new_n26701 = ~new_n26663 & ~new_n26700 ;
  assign new_n26702 = lo1432 & new_n26662 ;
  assign new_n26703 = ~lo1431 & ~new_n26693 ;
  assign new_n26704 = new_n26696 & ~new_n26703 ;
  assign new_n26705 = ~lo1432 & new_n26704 ;
  assign new_n26706 = lo1432 & ~new_n26704 ;
  assign new_n26707 = ~new_n26705 & ~new_n26706 ;
  assign new_n26708 = ~new_n16687 & ~new_n26707 ;
  assign new_n26709 = ~lo1269 & new_n16687 ;
  assign new_n26710 = ~new_n26708 & ~new_n26709 ;
  assign new_n26711 = ~new_n26662 & ~new_n26710 ;
  assign new_n26712 = ~new_n26702 & ~new_n26711 ;
  assign new_n26713 = lo1433 & new_n26662 ;
  assign new_n26714 = ~new_n16687 & ~new_n26677 ;
  assign new_n26715 = ~lo1275 & new_n16687 ;
  assign new_n26716 = ~new_n26714 & ~new_n26715 ;
  assign new_n26717 = ~new_n26662 & ~new_n26716 ;
  assign new_n26718 = ~new_n26713 & ~new_n26717 ;
  assign new_n26719 = lo0977 & new_n21253 ;
  assign new_n26720 = ~lo0977 & ~new_n21253 ;
  assign new_n26721 = ~new_n15793 & ~new_n26720 ;
  assign new_n26722 = ~new_n26719 & new_n26721 ;
  assign new_n26723 = new_n21249 & new_n26722 ;
  assign new_n26724 = ~lo0050 & lo1434 ;
  assign new_n26725 = ~new_n26723 & new_n26724 ;
  assign new_n26726 = lo0050 & lo1434 ;
  assign new_n26727 = ~lo0897 & new_n26726 ;
  assign new_n26728 = ~new_n26723 & new_n26727 ;
  assign new_n26729 = ~new_n26723 & ~new_n26728 ;
  assign new_n26730 = ~new_n26725 & new_n26729 ;
  assign new_n26731 = ~lo0017 & ~new_n26730 ;
  assign new_n26732 = lo1435 & new_n26662 ;
  assign new_n26733 = ~lo1432 & ~new_n26704 ;
  assign new_n26734 = new_n26707 & ~new_n26733 ;
  assign new_n26735 = ~lo1435 & new_n26734 ;
  assign new_n26736 = lo1435 & ~new_n26734 ;
  assign new_n26737 = ~new_n26735 & ~new_n26736 ;
  assign new_n26738 = ~new_n16687 & ~new_n26737 ;
  assign new_n26739 = ~lo1270 & new_n16687 ;
  assign new_n26740 = ~new_n26738 & ~new_n26739 ;
  assign new_n26741 = ~new_n26662 & ~new_n26740 ;
  assign new_n26742 = ~new_n26732 & ~new_n26741 ;
  assign new_n26743 = lo1436 & new_n26662 ;
  assign new_n26744 = ~lo1435 & ~new_n26734 ;
  assign new_n26745 = new_n26737 & ~new_n26744 ;
  assign new_n26746 = ~lo1437 & ~new_n26745 ;
  assign new_n26747 = ~lo1437 & new_n26745 ;
  assign new_n26748 = lo1437 & ~new_n26745 ;
  assign new_n26749 = ~new_n26747 & ~new_n26748 ;
  assign new_n26750 = ~new_n26746 & new_n26749 ;
  assign new_n26751 = ~lo1436 & new_n26750 ;
  assign new_n26752 = lo1436 & ~new_n26750 ;
  assign new_n26753 = ~new_n26751 & ~new_n26752 ;
  assign new_n26754 = ~new_n16687 & ~new_n26753 ;
  assign new_n26755 = ~lo1420 & new_n16687 ;
  assign new_n26756 = ~new_n26754 & ~new_n26755 ;
  assign new_n26757 = ~new_n26662 & ~new_n26756 ;
  assign new_n26758 = ~new_n26743 & ~new_n26757 ;
  assign new_n26759 = lo1437 & new_n26662 ;
  assign new_n26760 = ~new_n16687 & ~new_n26749 ;
  assign new_n26761 = ~lo1271 & new_n16687 ;
  assign new_n26762 = ~new_n26760 & ~new_n26761 ;
  assign new_n26763 = ~new_n26662 & ~new_n26762 ;
  assign new_n26764 = ~new_n26759 & ~new_n26763 ;
  assign new_n26765 = lo1438 & new_n26662 ;
  assign new_n26766 = ~new_n16687 & ~new_n26687 ;
  assign new_n26767 = ~lo1277 & new_n16687 ;
  assign new_n26768 = ~new_n26766 & ~new_n26767 ;
  assign new_n26769 = ~new_n26662 & ~new_n26768 ;
  assign new_n26770 = ~new_n26765 & ~new_n26769 ;
  assign new_n26771 = lo1439 & new_n26662 ;
  assign new_n26772 = ~new_n16687 & ~new_n26672 ;
  assign new_n26773 = ~lo1274 & new_n16687 ;
  assign new_n26774 = ~new_n26772 & ~new_n26773 ;
  assign new_n26775 = ~new_n26662 & ~new_n26774 ;
  assign new_n26776 = ~new_n26771 & ~new_n26775 ;
  assign new_n26777 = lo1440 & new_n26662 ;
  assign new_n26778 = ~new_n16687 & ~new_n26692 ;
  assign new_n26779 = ~lo1278 & new_n16687 ;
  assign new_n26780 = ~new_n26778 & ~new_n26779 ;
  assign new_n26781 = ~new_n26662 & ~new_n26780 ;
  assign new_n26782 = ~new_n26777 & ~new_n26781 ;
  assign new_n26783 = lo1441 & new_n26662 ;
  assign new_n26784 = ~new_n26664 & ~new_n26666 ;
  assign new_n26785 = ~new_n16687 & ~new_n26784 ;
  assign new_n26786 = ~lo1273 & new_n16687 ;
  assign new_n26787 = ~new_n26785 & ~new_n26786 ;
  assign new_n26788 = ~new_n26662 & ~new_n26787 ;
  assign new_n26789 = ~new_n26783 & ~new_n26788 ;
  assign new_n26790 = lo1442 & new_n26662 ;
  assign new_n26791 = ~new_n16687 & ~new_n26682 ;
  assign new_n26792 = ~lo1276 & new_n16687 ;
  assign new_n26793 = ~new_n26791 & ~new_n26792 ;
  assign new_n26794 = ~new_n26662 & ~new_n26793 ;
  assign new_n26795 = ~new_n26790 & ~new_n26794 ;
  assign new_n26796 = lo1443 & new_n26662 ;
  assign new_n26797 = ~lo1443 & ~new_n16687 ;
  assign new_n26798 = ~lo1272 & new_n16687 ;
  assign new_n26799 = ~new_n26797 & ~new_n26798 ;
  assign new_n26800 = ~new_n26662 & ~new_n26799 ;
  assign new_n26801 = ~new_n26796 & ~new_n26800 ;
  assign new_n26802 = lo1444 & ~new_n21479 ;
  assign new_n26803 = lo0112 & new_n14287 ;
  assign new_n26804 = new_n14287 & ~new_n26803 ;
  assign new_n26805 = ~new_n5880 & ~new_n26804 ;
  assign new_n26806 = ~lo0112 & new_n5880 ;
  assign new_n26807 = ~new_n14287 & new_n26806 ;
  assign new_n26808 = ~new_n26805 & ~new_n26807 ;
  assign new_n26809 = lo0113 & ~new_n26808 ;
  assign new_n26810 = ~new_n21672 & ~new_n26809 ;
  assign new_n26811 = new_n21479 & ~new_n26810 ;
  assign new_n26812 = ~new_n26802 & ~new_n26811 ;
  assign new_n26813 = lo1445 & ~new_n21479 ;
  assign new_n26814 = lo0112 & new_n14313 ;
  assign new_n26815 = new_n14313 & ~new_n26814 ;
  assign new_n26816 = ~new_n6106 & ~new_n26815 ;
  assign new_n26817 = ~lo0112 & new_n6106 ;
  assign new_n26818 = ~new_n14313 & new_n26817 ;
  assign new_n26819 = ~new_n26816 & ~new_n26818 ;
  assign new_n26820 = lo0113 & ~new_n26819 ;
  assign new_n26821 = ~new_n21561 & ~new_n26820 ;
  assign new_n26822 = new_n21479 & ~new_n26821 ;
  assign new_n26823 = ~new_n26813 & ~new_n26822 ;
  assign new_n26824 = lo1446 & ~new_n21479 ;
  assign new_n26825 = lo0112 & new_n14340 ;
  assign new_n26826 = new_n14340 & ~new_n26825 ;
  assign new_n26827 = ~new_n6336 & ~new_n26826 ;
  assign new_n26828 = ~lo0112 & new_n6336 ;
  assign new_n26829 = ~new_n14340 & new_n26828 ;
  assign new_n26830 = ~new_n26827 & ~new_n26829 ;
  assign new_n26831 = lo0113 & ~new_n26830 ;
  assign new_n26832 = ~new_n21492 & ~new_n26831 ;
  assign new_n26833 = new_n21479 & ~new_n26832 ;
  assign new_n26834 = ~new_n26824 & ~new_n26833 ;
  assign new_n26835 = lo1447 & new_n14661 ;
  assign new_n26836 = ~lo0017 & ~lo1434 ;
  assign new_n26837 = new_n15793 & new_n26836 ;
  assign new_n26838 = new_n15790 & new_n26837 ;
  assign new_n26839 = ~lo0017 & ~new_n26838 ;
  assign new_n26840 = ~new_n14661 & ~new_n26839 ;
  assign new_n26841 = ~new_n26835 & ~new_n26840 ;
  assign new_n26842 = ~lo1110 & lo1111 ;
  assign new_n26843 = ~lo1108 & new_n26842 ;
  assign new_n26844 = ~lo0017 & ~new_n26843 ;
  assign new_n26845 = lo1448 & ~new_n21836 ;
  assign new_n26846 = ~lo1448 & new_n21836 ;
  assign new_n26847 = ~new_n26845 & ~new_n26846 ;
  assign new_n26848 = new_n26844 & ~new_n26847 ;
  assign new_n26849 = lo1448 & new_n21836 ;
  assign new_n26850 = lo1449 & ~new_n26849 ;
  assign new_n26851 = ~lo1449 & new_n26849 ;
  assign new_n26852 = ~new_n26850 & ~new_n26851 ;
  assign new_n26853 = new_n26844 & ~new_n26852 ;
  assign new_n26854 = lo0017 & ~new_n26844 ;
  assign new_n26855 = ~new_n26853 & ~new_n26854 ;
  assign new_n26856 = lo1449 & new_n26849 ;
  assign new_n26857 = lo1450 & ~new_n26856 ;
  assign new_n26858 = ~lo1450 & new_n26856 ;
  assign new_n26859 = ~new_n26857 & ~new_n26858 ;
  assign new_n26860 = new_n26844 & ~new_n26859 ;
  assign new_n26861 = lo1450 & new_n26856 ;
  assign new_n26862 = lo1451 & ~new_n26861 ;
  assign new_n26863 = ~lo1451 & new_n26861 ;
  assign new_n26864 = ~new_n26862 & ~new_n26863 ;
  assign new_n26865 = new_n26844 & ~new_n26864 ;
  assign new_n26866 = ~new_n26854 & ~new_n26865 ;
  assign new_n26867 = ~lo0017 & ~lo1074 ;
  assign new_n26868 = lo1142 & lo1454 ;
  assign new_n26869 = lo1452 & ~new_n26868 ;
  assign new_n26870 = ~lo1452 & new_n26868 ;
  assign new_n26871 = ~new_n26869 & ~new_n26870 ;
  assign new_n26872 = new_n26867 & ~new_n26871 ;
  assign new_n26873 = lo1452 & new_n26868 ;
  assign new_n26874 = lo1459 & new_n26873 ;
  assign new_n26875 = lo1456 & new_n26874 ;
  assign new_n26876 = lo1457 & new_n26875 ;
  assign new_n26877 = lo1455 & new_n26876 ;
  assign new_n26878 = lo1458 & new_n26877 ;
  assign new_n26879 = lo1453 & ~new_n26878 ;
  assign new_n26880 = ~lo1453 & new_n26878 ;
  assign new_n26881 = ~new_n26879 & ~new_n26880 ;
  assign new_n26882 = new_n26867 & ~new_n26881 ;
  assign new_n26883 = ~lo1142 & lo1454 ;
  assign new_n26884 = lo1142 & ~lo1454 ;
  assign new_n26885 = ~new_n26883 & ~new_n26884 ;
  assign new_n26886 = new_n26867 & ~new_n26885 ;
  assign new_n26887 = lo1455 & ~new_n26876 ;
  assign new_n26888 = ~lo1455 & new_n26876 ;
  assign new_n26889 = ~new_n26887 & ~new_n26888 ;
  assign new_n26890 = new_n26867 & ~new_n26889 ;
  assign new_n26891 = lo1456 & ~new_n26874 ;
  assign new_n26892 = ~lo1456 & new_n26874 ;
  assign new_n26893 = ~new_n26891 & ~new_n26892 ;
  assign new_n26894 = new_n26867 & ~new_n26893 ;
  assign new_n26895 = lo1457 & ~new_n26875 ;
  assign new_n26896 = ~lo1457 & new_n26875 ;
  assign new_n26897 = ~new_n26895 & ~new_n26896 ;
  assign new_n26898 = new_n26867 & ~new_n26897 ;
  assign new_n26899 = lo1458 & ~new_n26877 ;
  assign new_n26900 = ~lo1458 & new_n26877 ;
  assign new_n26901 = ~new_n26899 & ~new_n26900 ;
  assign new_n26902 = new_n26867 & ~new_n26901 ;
  assign new_n26903 = lo1459 & ~new_n26873 ;
  assign new_n26904 = ~lo1459 & new_n26873 ;
  assign new_n26905 = ~new_n26903 & ~new_n26904 ;
  assign new_n26906 = new_n26867 & ~new_n26905 ;
  assign new_n26907 = ~lo0017 & ~lo1142 ;
  assign new_n26908 = lo1460 & ~lo1462 ;
  assign new_n26909 = ~lo1460 & lo1462 ;
  assign new_n26910 = ~new_n26908 & ~new_n26909 ;
  assign new_n26911 = new_n26907 & ~new_n26910 ;
  assign new_n26912 = lo1460 & lo1462 ;
  assign new_n26913 = lo1467 & new_n26912 ;
  assign new_n26914 = lo1464 & new_n26913 ;
  assign new_n26915 = lo1465 & new_n26914 ;
  assign new_n26916 = lo1463 & new_n26915 ;
  assign new_n26917 = lo1466 & new_n26916 ;
  assign new_n26918 = lo1461 & ~new_n26917 ;
  assign new_n26919 = ~lo1461 & new_n26917 ;
  assign new_n26920 = ~new_n26918 & ~new_n26919 ;
  assign new_n26921 = new_n26907 & ~new_n26920 ;
  assign new_n26922 = ~lo1462 & new_n26907 ;
  assign new_n26923 = lo1463 & ~new_n26915 ;
  assign new_n26924 = ~lo1463 & new_n26915 ;
  assign new_n26925 = ~new_n26923 & ~new_n26924 ;
  assign new_n26926 = new_n26907 & ~new_n26925 ;
  assign new_n26927 = lo1464 & ~new_n26913 ;
  assign new_n26928 = ~lo1464 & new_n26913 ;
  assign new_n26929 = ~new_n26927 & ~new_n26928 ;
  assign new_n26930 = new_n26907 & ~new_n26929 ;
  assign new_n26931 = lo1465 & ~new_n26914 ;
  assign new_n26932 = ~lo1465 & new_n26914 ;
  assign new_n26933 = ~new_n26931 & ~new_n26932 ;
  assign new_n26934 = new_n26907 & ~new_n26933 ;
  assign new_n26935 = lo1466 & ~new_n26916 ;
  assign new_n26936 = ~lo1466 & new_n26916 ;
  assign new_n26937 = ~new_n26935 & ~new_n26936 ;
  assign new_n26938 = new_n26907 & ~new_n26937 ;
  assign new_n26939 = lo1467 & ~new_n26912 ;
  assign new_n26940 = ~lo1467 & new_n26912 ;
  assign new_n26941 = ~new_n26939 & ~new_n26940 ;
  assign new_n26942 = new_n26907 & ~new_n26941 ;
  assign new_n26943 = lo1110 & lo1111 ;
  assign new_n26944 = ~lo1110 & ~lo1111 ;
  assign new_n26945 = ~new_n26943 & ~new_n26944 ;
  assign new_n26946 = ~lo1245 & lo1468 ;
  assign new_n26947 = ~new_n26945 & new_n26946 ;
  assign new_n26948 = lo1110 & ~lo1111 ;
  assign new_n26949 = ~new_n26842 & ~new_n26948 ;
  assign new_n26950 = ~new_n26947 & new_n26949 ;
  assign new_n26951 = ~lo0017 & ~new_n26950 ;
  assign new_n26952 = lo0112 & new_n14005 ;
  assign new_n26953 = new_n14005 & ~new_n26952 ;
  assign new_n26954 = ~new_n7761 & ~new_n26953 ;
  assign new_n26955 = ~lo0112 & new_n7761 ;
  assign new_n26956 = ~new_n14005 & new_n26955 ;
  assign new_n26957 = ~new_n26954 & ~new_n26956 ;
  assign new_n26958 = lo0112 & new_n14578 ;
  assign new_n26959 = new_n14578 & ~new_n26958 ;
  assign new_n26960 = ~new_n8008 & ~new_n26959 ;
  assign new_n26961 = ~lo0112 & new_n8008 ;
  assign new_n26962 = ~new_n14578 & new_n26961 ;
  assign new_n26963 = ~new_n26960 & ~new_n26962 ;
  assign new_n26964 = lo0112 & new_n14552 ;
  assign new_n26965 = new_n14552 & ~new_n26964 ;
  assign new_n26966 = ~new_n7883 & ~new_n26965 ;
  assign new_n26967 = ~lo0112 & new_n7883 ;
  assign new_n26968 = ~new_n14552 & new_n26967 ;
  assign new_n26969 = ~new_n26966 & ~new_n26968 ;
  assign new_n26970 = lo0112 & new_n14499 ;
  assign new_n26971 = new_n14499 & ~new_n26970 ;
  assign new_n26972 = ~new_n7637 & ~new_n26971 ;
  assign new_n26973 = ~lo0112 & new_n7637 ;
  assign new_n26974 = ~new_n14499 & new_n26973 ;
  assign new_n26975 = ~new_n26972 & ~new_n26974 ;
  assign new_n26976 = lo0112 & new_n14472 ;
  assign new_n26977 = new_n14472 & ~new_n26976 ;
  assign new_n26978 = ~new_n7512 & ~new_n26977 ;
  assign new_n26979 = ~lo0112 & new_n7512 ;
  assign new_n26980 = ~new_n14472 & new_n26979 ;
  assign new_n26981 = ~new_n26978 & ~new_n26980 ;
  assign new_n26982 = lo0112 & new_n13936 ;
  assign new_n26983 = new_n13936 & ~new_n26982 ;
  assign new_n26984 = ~new_n8411 & ~new_n26983 ;
  assign new_n26985 = ~lo0112 & new_n8411 ;
  assign new_n26986 = ~new_n13936 & new_n26985 ;
  assign new_n26987 = ~new_n26984 & ~new_n26986 ;
  assign new_n26988 = lo0112 & new_n13977 ;
  assign new_n26989 = new_n13977 & ~new_n26988 ;
  assign new_n26990 = ~new_n8281 & ~new_n26989 ;
  assign new_n26991 = ~lo0112 & new_n8281 ;
  assign new_n26992 = ~new_n13977 & new_n26991 ;
  assign new_n26993 = ~new_n26990 & ~new_n26992 ;
  assign new_n26994 = lo0112 & new_n14525 ;
  assign new_n26995 = new_n14525 & ~new_n26994 ;
  assign new_n26996 = ~new_n8149 & ~new_n26995 ;
  assign new_n26997 = ~lo0112 & new_n8149 ;
  assign new_n26998 = ~new_n14525 & new_n26997 ;
  assign new_n26999 = ~new_n26996 & ~new_n26998 ;
  assign po0000 = lo0000 ;
  assign po0001 = lo0001 ;
  assign po0002 = lo0002 ;
  assign po0003 = lo0003 ;
  assign po0004 = lo0004 ;
  assign po0005 = lo0005 ;
  assign po0006 = lo0006 ;
  assign po0007 = lo0007 ;
  assign po0008 = lo0008 ;
  assign po0009 = lo0009 ;
  assign po0010 = lo0010 ;
  assign po0011 = lo0011 ;
  assign po0012 = lo0012 ;
  assign po0013 = lo0013 ;
  assign po0014 = lo0014 ;
  assign po0015 = lo0015 ;
  assign po0016 = lo1268 ;
  assign po0017 = lo0016 ;
  assign po0018 = new_n1974 ;
  assign po0019 = pi000 ;
  assign po0020 = lo1444 ;
  assign po0021 = lo0917 ;
  assign po0022 = lo1060 ;
  assign po0023 = lo1056 ;
  assign po0024 = lo1057 ;
  assign po0025 = lo1059 ;
  assign po0026 = lo1058 ;
  assign po0027 = lo0019 ;
  assign po0028 = lo0020 ;
  assign po0029 = lo0040 ;
  assign po0030 = new_n1977 ;
  assign po0031 = pi000 ;
  assign po0032 = lo1444 ;
  assign po0033 = lo0917 ;
  assign po0034 = lo1060 ;
  assign po0035 = lo1056 ;
  assign po0036 = lo1057 ;
  assign po0037 = lo1059 ;
  assign po0038 = lo1058 ;
  assign po0039 = lo0019 ;
  assign po0040 = lo0020 ;
  assign po0041 = lo0040 ;
  assign po0042 = new_n1980 ;
  assign po0043 = pi000 ;
  assign po0044 = lo1444 ;
  assign po0045 = lo0917 ;
  assign po0046 = lo1060 ;
  assign po0047 = lo1056 ;
  assign po0048 = lo1057 ;
  assign po0049 = lo1059 ;
  assign po0050 = lo1058 ;
  assign po0051 = lo0019 ;
  assign po0052 = lo0020 ;
  assign po0053 = lo0040 ;
  assign po0054 = new_n1983 ;
  assign po0055 = pi000 ;
  assign po0056 = lo1444 ;
  assign po0057 = lo0917 ;
  assign po0058 = lo1060 ;
  assign po0059 = lo1056 ;
  assign po0060 = lo1057 ;
  assign po0061 = lo1059 ;
  assign po0062 = lo1058 ;
  assign po0063 = lo0019 ;
  assign po0064 = lo0020 ;
  assign po0065 = lo0040 ;
  assign po0066 = new_n1986 ;
  assign po0067 = pi000 ;
  assign po0068 = lo1444 ;
  assign po0069 = lo0917 ;
  assign po0070 = lo1060 ;
  assign po0071 = lo1056 ;
  assign po0072 = lo1057 ;
  assign po0073 = lo1059 ;
  assign po0074 = lo1058 ;
  assign po0075 = lo0019 ;
  assign po0076 = lo0020 ;
  assign po0077 = lo0040 ;
  assign po0078 = new_n1988 ;
  assign po0079 = pi000 ;
  assign po0080 = lo1444 ;
  assign po0081 = lo0917 ;
  assign po0082 = lo1060 ;
  assign po0083 = lo1056 ;
  assign po0084 = lo1057 ;
  assign po0085 = lo1059 ;
  assign po0086 = lo1058 ;
  assign po0087 = lo0019 ;
  assign po0088 = lo0020 ;
  assign po0089 = lo0040 ;
  assign po0090 = new_n1990 ;
  assign po0091 = pi000 ;
  assign po0092 = lo1444 ;
  assign po0093 = lo0917 ;
  assign po0094 = lo1060 ;
  assign po0095 = lo1056 ;
  assign po0096 = lo1057 ;
  assign po0097 = lo1059 ;
  assign po0098 = lo1058 ;
  assign po0099 = lo0019 ;
  assign po0100 = lo0020 ;
  assign po0101 = lo0040 ;
  assign po0102 = new_n1992 ;
  assign po0103 = pi000 ;
  assign po0104 = lo1444 ;
  assign po0105 = lo0917 ;
  assign po0106 = lo1060 ;
  assign po0107 = lo1056 ;
  assign po0108 = lo1057 ;
  assign po0109 = lo1059 ;
  assign po0110 = lo1058 ;
  assign po0111 = lo0019 ;
  assign po0112 = lo0020 ;
  assign po0113 = lo0040 ;
  assign po0114 = new_n1994 ;
  assign po0115 = pi000 ;
  assign po0116 = lo1424 ;
  assign po0117 = lo0917 ;
  assign po0118 = lo1060 ;
  assign po0119 = lo1056 ;
  assign po0120 = lo1057 ;
  assign po0121 = lo1059 ;
  assign po0122 = lo1058 ;
  assign po0123 = lo0019 ;
  assign po0124 = lo0020 ;
  assign po0125 = lo0040 ;
  assign po0126 = new_n1995 ;
  assign po0127 = pi000 ;
  assign po0128 = lo1424 ;
  assign po0129 = lo0917 ;
  assign po0130 = lo1060 ;
  assign po0131 = lo1056 ;
  assign po0132 = lo1057 ;
  assign po0133 = lo1059 ;
  assign po0134 = lo1058 ;
  assign po0135 = lo0019 ;
  assign po0136 = lo0020 ;
  assign po0137 = lo0040 ;
  assign po0138 = new_n1996 ;
  assign po0139 = pi000 ;
  assign po0140 = lo1424 ;
  assign po0141 = lo0917 ;
  assign po0142 = lo1060 ;
  assign po0143 = lo1056 ;
  assign po0144 = lo1057 ;
  assign po0145 = lo1059 ;
  assign po0146 = lo1058 ;
  assign po0147 = lo0019 ;
  assign po0148 = lo0020 ;
  assign po0149 = lo0040 ;
  assign po0150 = new_n1997 ;
  assign po0151 = pi000 ;
  assign po0152 = lo1424 ;
  assign po0153 = lo0917 ;
  assign po0154 = lo1060 ;
  assign po0155 = lo1056 ;
  assign po0156 = lo1057 ;
  assign po0157 = lo1059 ;
  assign po0158 = lo1058 ;
  assign po0159 = lo0019 ;
  assign po0160 = lo0020 ;
  assign po0161 = lo0040 ;
  assign po0162 = new_n1998 ;
  assign po0163 = pi000 ;
  assign po0164 = lo1424 ;
  assign po0165 = lo0917 ;
  assign po0166 = lo1060 ;
  assign po0167 = lo1056 ;
  assign po0168 = lo1057 ;
  assign po0169 = lo1059 ;
  assign po0170 = lo1058 ;
  assign po0171 = lo0019 ;
  assign po0172 = lo0020 ;
  assign po0173 = lo0040 ;
  assign po0174 = new_n1999 ;
  assign po0175 = pi000 ;
  assign po0176 = lo1424 ;
  assign po0177 = lo0917 ;
  assign po0178 = lo1060 ;
  assign po0179 = lo1056 ;
  assign po0180 = lo1057 ;
  assign po0181 = lo1059 ;
  assign po0182 = lo1058 ;
  assign po0183 = lo0019 ;
  assign po0184 = lo0020 ;
  assign po0185 = lo0040 ;
  assign po0186 = new_n2000 ;
  assign po0187 = pi000 ;
  assign po0188 = lo1424 ;
  assign po0189 = lo0917 ;
  assign po0190 = lo1060 ;
  assign po0191 = lo1056 ;
  assign po0192 = lo1057 ;
  assign po0193 = lo1059 ;
  assign po0194 = lo1058 ;
  assign po0195 = lo0019 ;
  assign po0196 = lo0020 ;
  assign po0197 = lo0040 ;
  assign po0198 = new_n2001 ;
  assign po0199 = pi000 ;
  assign po0200 = lo1424 ;
  assign po0201 = lo0917 ;
  assign po0202 = lo1060 ;
  assign po0203 = lo1056 ;
  assign po0204 = lo1057 ;
  assign po0205 = lo1059 ;
  assign po0206 = lo1058 ;
  assign po0207 = lo0019 ;
  assign po0208 = lo0020 ;
  assign po0209 = lo0040 ;
  assign po0210 = new_n2003 ;
  assign po0211 = pi000 ;
  assign po0212 = lo1061 ;
  assign po0213 = lo0917 ;
  assign po0214 = lo1060 ;
  assign po0215 = lo1056 ;
  assign po0216 = lo1057 ;
  assign po0217 = lo1059 ;
  assign po0218 = lo1058 ;
  assign po0219 = lo0019 ;
  assign po0220 = lo0020 ;
  assign po0221 = lo0040 ;
  assign po0222 = new_n2004 ;
  assign po0223 = pi000 ;
  assign po0224 = lo1061 ;
  assign po0225 = lo0917 ;
  assign po0226 = lo1060 ;
  assign po0227 = lo1056 ;
  assign po0228 = lo1057 ;
  assign po0229 = lo1059 ;
  assign po0230 = lo1058 ;
  assign po0231 = lo0019 ;
  assign po0232 = lo0020 ;
  assign po0233 = lo0040 ;
  assign po0234 = new_n2005 ;
  assign po0235 = pi000 ;
  assign po0236 = lo1061 ;
  assign po0237 = lo0917 ;
  assign po0238 = lo1060 ;
  assign po0239 = lo1056 ;
  assign po0240 = lo1057 ;
  assign po0241 = lo1059 ;
  assign po0242 = lo1058 ;
  assign po0243 = lo0019 ;
  assign po0244 = lo0020 ;
  assign po0245 = lo0040 ;
  assign po0246 = new_n2006 ;
  assign po0247 = pi000 ;
  assign po0248 = lo1061 ;
  assign po0249 = lo0917 ;
  assign po0250 = lo1060 ;
  assign po0251 = lo1056 ;
  assign po0252 = lo1057 ;
  assign po0253 = lo1059 ;
  assign po0254 = lo1058 ;
  assign po0255 = lo0019 ;
  assign po0256 = lo0020 ;
  assign po0257 = lo0040 ;
  assign po0258 = new_n2007 ;
  assign po0259 = pi000 ;
  assign po0260 = lo1061 ;
  assign po0261 = lo0917 ;
  assign po0262 = lo1060 ;
  assign po0263 = lo1056 ;
  assign po0264 = lo1057 ;
  assign po0265 = lo1059 ;
  assign po0266 = lo1058 ;
  assign po0267 = lo0019 ;
  assign po0268 = lo0020 ;
  assign po0269 = lo0040 ;
  assign po0270 = new_n2008 ;
  assign po0271 = pi000 ;
  assign po0272 = lo1061 ;
  assign po0273 = lo0917 ;
  assign po0274 = lo1060 ;
  assign po0275 = lo1056 ;
  assign po0276 = lo1057 ;
  assign po0277 = lo1059 ;
  assign po0278 = lo1058 ;
  assign po0279 = lo0019 ;
  assign po0280 = lo0020 ;
  assign po0281 = lo0040 ;
  assign po0282 = new_n2009 ;
  assign po0283 = pi000 ;
  assign po0284 = lo1061 ;
  assign po0285 = lo0917 ;
  assign po0286 = lo1060 ;
  assign po0287 = lo1056 ;
  assign po0288 = lo1057 ;
  assign po0289 = lo1059 ;
  assign po0290 = lo1058 ;
  assign po0291 = lo0019 ;
  assign po0292 = lo0020 ;
  assign po0293 = lo0040 ;
  assign po0294 = new_n2010 ;
  assign po0295 = pi000 ;
  assign po0296 = lo1061 ;
  assign po0297 = lo0917 ;
  assign po0298 = lo1060 ;
  assign po0299 = lo1056 ;
  assign po0300 = lo1057 ;
  assign po0301 = lo1059 ;
  assign po0302 = lo1058 ;
  assign po0303 = lo0019 ;
  assign po0304 = lo0020 ;
  assign po0305 = lo0040 ;
  assign po0306 = new_n2012 ;
  assign po0307 = pi000 ;
  assign po0308 = lo1279 ;
  assign po0309 = lo0917 ;
  assign po0310 = lo1060 ;
  assign po0311 = lo1056 ;
  assign po0312 = lo1057 ;
  assign po0313 = lo1059 ;
  assign po0314 = lo1058 ;
  assign po0315 = lo0019 ;
  assign po0316 = lo0020 ;
  assign po0317 = lo0040 ;
  assign po0318 = new_n2013 ;
  assign po0319 = pi000 ;
  assign po0320 = lo1279 ;
  assign po0321 = lo0917 ;
  assign po0322 = lo1060 ;
  assign po0323 = lo1056 ;
  assign po0324 = lo1057 ;
  assign po0325 = lo1059 ;
  assign po0326 = lo1058 ;
  assign po0327 = lo0019 ;
  assign po0328 = lo0020 ;
  assign po0329 = lo0040 ;
  assign po0330 = new_n2014 ;
  assign po0331 = pi000 ;
  assign po0332 = lo1279 ;
  assign po0333 = lo0917 ;
  assign po0334 = lo1060 ;
  assign po0335 = lo1056 ;
  assign po0336 = lo1057 ;
  assign po0337 = lo1059 ;
  assign po0338 = lo1058 ;
  assign po0339 = lo0019 ;
  assign po0340 = lo0020 ;
  assign po0341 = lo0040 ;
  assign po0342 = new_n2015 ;
  assign po0343 = pi000 ;
  assign po0344 = lo1279 ;
  assign po0345 = lo0917 ;
  assign po0346 = lo1060 ;
  assign po0347 = lo1056 ;
  assign po0348 = lo1057 ;
  assign po0349 = lo1059 ;
  assign po0350 = lo1058 ;
  assign po0351 = lo0019 ;
  assign po0352 = lo0020 ;
  assign po0353 = lo0040 ;
  assign po0354 = new_n2016 ;
  assign po0355 = pi000 ;
  assign po0356 = lo1279 ;
  assign po0357 = lo0917 ;
  assign po0358 = lo1060 ;
  assign po0359 = lo1056 ;
  assign po0360 = lo1057 ;
  assign po0361 = lo1059 ;
  assign po0362 = lo1058 ;
  assign po0363 = lo0019 ;
  assign po0364 = lo0020 ;
  assign po0365 = lo0040 ;
  assign po0366 = new_n2017 ;
  assign po0367 = pi000 ;
  assign po0368 = lo1279 ;
  assign po0369 = lo0917 ;
  assign po0370 = lo1060 ;
  assign po0371 = lo1056 ;
  assign po0372 = lo1057 ;
  assign po0373 = lo1059 ;
  assign po0374 = lo1058 ;
  assign po0375 = lo0019 ;
  assign po0376 = lo0020 ;
  assign po0377 = lo0040 ;
  assign po0378 = new_n2018 ;
  assign po0379 = pi000 ;
  assign po0380 = lo1279 ;
  assign po0381 = lo0917 ;
  assign po0382 = lo1060 ;
  assign po0383 = lo1056 ;
  assign po0384 = lo1057 ;
  assign po0385 = lo1059 ;
  assign po0386 = lo1058 ;
  assign po0387 = lo0019 ;
  assign po0388 = lo0020 ;
  assign po0389 = lo0040 ;
  assign po0390 = new_n2019 ;
  assign po0391 = pi000 ;
  assign po0392 = lo1279 ;
  assign po0393 = lo0917 ;
  assign po0394 = lo1060 ;
  assign po0395 = lo1056 ;
  assign po0396 = lo1057 ;
  assign po0397 = lo1059 ;
  assign po0398 = lo1058 ;
  assign po0399 = lo0019 ;
  assign po0400 = lo0020 ;
  assign po0401 = lo0040 ;
  assign po0402 = new_n2000 ;
  assign po0403 = pi000 ;
  assign po0404 = lo1269 ;
  assign po0405 = lo0917 ;
  assign po0406 = lo1060 ;
  assign po0407 = lo1056 ;
  assign po0408 = lo1057 ;
  assign po0409 = lo1059 ;
  assign po0410 = lo1058 ;
  assign po0411 = lo0019 ;
  assign po0412 = lo0020 ;
  assign po0413 = lo0040 ;
  assign po0414 = new_n1998 ;
  assign po0415 = pi000 ;
  assign po0416 = lo1269 ;
  assign po0417 = lo0917 ;
  assign po0418 = lo1060 ;
  assign po0419 = lo1056 ;
  assign po0420 = lo1057 ;
  assign po0421 = lo1059 ;
  assign po0422 = lo1058 ;
  assign po0423 = lo0019 ;
  assign po0424 = lo0020 ;
  assign po0425 = lo0040 ;
  assign po0426 = new_n1996 ;
  assign po0427 = pi000 ;
  assign po0428 = lo1269 ;
  assign po0429 = lo0917 ;
  assign po0430 = lo1060 ;
  assign po0431 = lo1056 ;
  assign po0432 = lo1057 ;
  assign po0433 = lo1059 ;
  assign po0434 = lo1058 ;
  assign po0435 = lo0019 ;
  assign po0436 = lo0020 ;
  assign po0437 = lo0040 ;
  assign po0438 = new_n1997 ;
  assign po0439 = pi000 ;
  assign po0440 = lo1269 ;
  assign po0441 = lo0917 ;
  assign po0442 = lo1060 ;
  assign po0443 = lo1056 ;
  assign po0444 = lo1057 ;
  assign po0445 = lo1059 ;
  assign po0446 = lo1058 ;
  assign po0447 = lo0019 ;
  assign po0448 = lo0020 ;
  assign po0449 = lo0040 ;
  assign po0450 = new_n1999 ;
  assign po0451 = pi000 ;
  assign po0452 = lo1269 ;
  assign po0453 = lo0917 ;
  assign po0454 = lo1060 ;
  assign po0455 = lo1056 ;
  assign po0456 = lo1057 ;
  assign po0457 = lo1059 ;
  assign po0458 = lo1058 ;
  assign po0459 = lo0019 ;
  assign po0460 = lo0020 ;
  assign po0461 = lo0040 ;
  assign po0462 = new_n1994 ;
  assign po0463 = pi000 ;
  assign po0464 = lo1269 ;
  assign po0465 = lo0917 ;
  assign po0466 = lo1060 ;
  assign po0467 = lo1056 ;
  assign po0468 = lo1057 ;
  assign po0469 = lo1059 ;
  assign po0470 = lo1058 ;
  assign po0471 = lo0019 ;
  assign po0472 = lo0020 ;
  assign po0473 = lo0040 ;
  assign po0474 = new_n1995 ;
  assign po0475 = pi000 ;
  assign po0476 = lo1269 ;
  assign po0477 = lo0917 ;
  assign po0478 = lo1060 ;
  assign po0479 = lo1056 ;
  assign po0480 = lo1057 ;
  assign po0481 = lo1059 ;
  assign po0482 = lo1058 ;
  assign po0483 = lo0019 ;
  assign po0484 = lo0020 ;
  assign po0485 = lo0040 ;
  assign po0486 = new_n2001 ;
  assign po0487 = pi000 ;
  assign po0488 = lo1269 ;
  assign po0489 = lo0917 ;
  assign po0490 = lo1060 ;
  assign po0491 = lo1056 ;
  assign po0492 = lo1057 ;
  assign po0493 = lo1059 ;
  assign po0494 = lo1058 ;
  assign po0495 = lo0019 ;
  assign po0496 = lo0020 ;
  assign po0497 = lo0040 ;
  assign po0498 = new_n2009 ;
  assign po0499 = pi000 ;
  assign po0500 = lo1078 ;
  assign po0501 = lo0917 ;
  assign po0502 = lo1060 ;
  assign po0503 = lo1056 ;
  assign po0504 = lo1057 ;
  assign po0505 = lo1059 ;
  assign po0506 = lo1058 ;
  assign po0507 = lo0019 ;
  assign po0508 = lo0020 ;
  assign po0509 = lo0040 ;
  assign po0510 = new_n2005 ;
  assign po0511 = pi000 ;
  assign po0512 = lo1078 ;
  assign po0513 = lo0917 ;
  assign po0514 = lo1060 ;
  assign po0515 = lo1056 ;
  assign po0516 = lo1057 ;
  assign po0517 = lo1059 ;
  assign po0518 = lo1058 ;
  assign po0519 = lo0019 ;
  assign po0520 = lo0020 ;
  assign po0521 = lo0040 ;
  assign po0522 = new_n2006 ;
  assign po0523 = pi000 ;
  assign po0524 = lo1078 ;
  assign po0525 = lo0917 ;
  assign po0526 = lo1060 ;
  assign po0527 = lo1056 ;
  assign po0528 = lo1057 ;
  assign po0529 = lo1059 ;
  assign po0530 = lo1058 ;
  assign po0531 = lo0019 ;
  assign po0532 = lo0020 ;
  assign po0533 = lo0040 ;
  assign po0534 = new_n2007 ;
  assign po0535 = pi000 ;
  assign po0536 = lo1078 ;
  assign po0537 = lo0917 ;
  assign po0538 = lo1060 ;
  assign po0539 = lo1056 ;
  assign po0540 = lo1057 ;
  assign po0541 = lo1059 ;
  assign po0542 = lo1058 ;
  assign po0543 = lo0019 ;
  assign po0544 = lo0020 ;
  assign po0545 = lo0040 ;
  assign po0546 = new_n2008 ;
  assign po0547 = pi000 ;
  assign po0548 = lo1078 ;
  assign po0549 = lo0917 ;
  assign po0550 = lo1060 ;
  assign po0551 = lo1056 ;
  assign po0552 = lo1057 ;
  assign po0553 = lo1059 ;
  assign po0554 = lo1058 ;
  assign po0555 = lo0019 ;
  assign po0556 = lo0020 ;
  assign po0557 = lo0040 ;
  assign po0558 = new_n2003 ;
  assign po0559 = pi000 ;
  assign po0560 = lo1078 ;
  assign po0561 = lo0917 ;
  assign po0562 = lo1060 ;
  assign po0563 = lo1056 ;
  assign po0564 = lo1057 ;
  assign po0565 = lo1059 ;
  assign po0566 = lo1058 ;
  assign po0567 = lo0019 ;
  assign po0568 = lo0020 ;
  assign po0569 = lo0040 ;
  assign po0570 = new_n2004 ;
  assign po0571 = pi000 ;
  assign po0572 = lo1078 ;
  assign po0573 = lo0917 ;
  assign po0574 = lo1060 ;
  assign po0575 = lo1056 ;
  assign po0576 = lo1057 ;
  assign po0577 = lo1059 ;
  assign po0578 = lo1058 ;
  assign po0579 = lo0019 ;
  assign po0580 = lo0020 ;
  assign po0581 = lo0040 ;
  assign po0582 = new_n2010 ;
  assign po0583 = pi000 ;
  assign po0584 = lo1078 ;
  assign po0585 = lo0917 ;
  assign po0586 = lo1060 ;
  assign po0587 = lo1056 ;
  assign po0588 = lo1057 ;
  assign po0589 = lo1059 ;
  assign po0590 = lo1058 ;
  assign po0591 = lo0019 ;
  assign po0592 = lo0020 ;
  assign po0593 = lo0040 ;
  assign po0594 = new_n2012 ;
  assign po0595 = pi000 ;
  assign po0596 = lo1275 ;
  assign po0597 = lo0917 ;
  assign po0598 = lo1060 ;
  assign po0599 = lo1056 ;
  assign po0600 = lo1057 ;
  assign po0601 = lo1059 ;
  assign po0602 = lo1058 ;
  assign po0603 = lo0019 ;
  assign po0604 = lo0020 ;
  assign po0605 = lo0040 ;
  assign po0606 = new_n2013 ;
  assign po0607 = pi000 ;
  assign po0608 = lo1275 ;
  assign po0609 = lo0917 ;
  assign po0610 = lo1060 ;
  assign po0611 = lo1056 ;
  assign po0612 = lo1057 ;
  assign po0613 = lo1059 ;
  assign po0614 = lo1058 ;
  assign po0615 = lo0019 ;
  assign po0616 = lo0020 ;
  assign po0617 = lo0040 ;
  assign po0618 = new_n2014 ;
  assign po0619 = pi000 ;
  assign po0620 = lo1275 ;
  assign po0621 = lo0917 ;
  assign po0622 = lo1060 ;
  assign po0623 = lo1056 ;
  assign po0624 = lo1057 ;
  assign po0625 = lo1059 ;
  assign po0626 = lo1058 ;
  assign po0627 = lo0019 ;
  assign po0628 = lo0020 ;
  assign po0629 = lo0040 ;
  assign po0630 = new_n2015 ;
  assign po0631 = pi000 ;
  assign po0632 = lo1275 ;
  assign po0633 = lo0917 ;
  assign po0634 = lo1060 ;
  assign po0635 = lo1056 ;
  assign po0636 = lo1057 ;
  assign po0637 = lo1059 ;
  assign po0638 = lo1058 ;
  assign po0639 = lo0019 ;
  assign po0640 = lo0020 ;
  assign po0641 = lo0040 ;
  assign po0642 = new_n2016 ;
  assign po0643 = pi000 ;
  assign po0644 = lo1275 ;
  assign po0645 = lo0917 ;
  assign po0646 = lo1060 ;
  assign po0647 = lo1056 ;
  assign po0648 = lo1057 ;
  assign po0649 = lo1059 ;
  assign po0650 = lo1058 ;
  assign po0651 = lo0019 ;
  assign po0652 = lo0020 ;
  assign po0653 = lo0040 ;
  assign po0654 = new_n2017 ;
  assign po0655 = pi000 ;
  assign po0656 = lo1275 ;
  assign po0657 = lo0917 ;
  assign po0658 = lo1060 ;
  assign po0659 = lo1056 ;
  assign po0660 = lo1057 ;
  assign po0661 = lo1059 ;
  assign po0662 = lo1058 ;
  assign po0663 = lo0019 ;
  assign po0664 = lo0020 ;
  assign po0665 = lo0040 ;
  assign po0666 = new_n2018 ;
  assign po0667 = pi000 ;
  assign po0668 = lo1275 ;
  assign po0669 = lo0917 ;
  assign po0670 = lo1060 ;
  assign po0671 = lo1056 ;
  assign po0672 = lo1057 ;
  assign po0673 = lo1059 ;
  assign po0674 = lo1058 ;
  assign po0675 = lo0019 ;
  assign po0676 = lo0020 ;
  assign po0677 = lo0040 ;
  assign po0678 = new_n2019 ;
  assign po0679 = pi000 ;
  assign po0680 = lo1275 ;
  assign po0681 = lo0917 ;
  assign po0682 = lo1060 ;
  assign po0683 = lo1056 ;
  assign po0684 = lo1057 ;
  assign po0685 = lo1059 ;
  assign po0686 = lo1058 ;
  assign po0687 = lo0019 ;
  assign po0688 = lo0020 ;
  assign po0689 = lo0040 ;
  assign po0690 = new_n1988 ;
  assign po0691 = pi000 ;
  assign po0692 = lo1283 ;
  assign po0693 = lo0917 ;
  assign po0694 = lo1060 ;
  assign po0695 = lo1056 ;
  assign po0696 = lo1057 ;
  assign po0697 = lo1059 ;
  assign po0698 = lo1058 ;
  assign po0699 = lo0019 ;
  assign po0700 = lo0020 ;
  assign po0701 = lo0040 ;
  assign po0702 = new_n1992 ;
  assign po0703 = pi000 ;
  assign po0704 = lo1283 ;
  assign po0705 = lo0917 ;
  assign po0706 = lo1060 ;
  assign po0707 = lo1056 ;
  assign po0708 = lo1057 ;
  assign po0709 = lo1059 ;
  assign po0710 = lo1058 ;
  assign po0711 = lo0019 ;
  assign po0712 = lo0020 ;
  assign po0713 = lo0040 ;
  assign po0714 = new_n1990 ;
  assign po0715 = pi000 ;
  assign po0716 = lo1283 ;
  assign po0717 = lo0917 ;
  assign po0718 = lo1060 ;
  assign po0719 = lo1056 ;
  assign po0720 = lo1057 ;
  assign po0721 = lo1059 ;
  assign po0722 = lo1058 ;
  assign po0723 = lo0019 ;
  assign po0724 = lo0020 ;
  assign po0725 = lo0040 ;
  assign po0726 = new_n1974 ;
  assign po0727 = pi000 ;
  assign po0728 = lo1283 ;
  assign po0729 = lo0917 ;
  assign po0730 = lo1060 ;
  assign po0731 = lo1056 ;
  assign po0732 = lo1057 ;
  assign po0733 = lo1059 ;
  assign po0734 = lo1058 ;
  assign po0735 = lo0019 ;
  assign po0736 = lo0020 ;
  assign po0737 = lo0040 ;
  assign po0738 = new_n1977 ;
  assign po0739 = pi000 ;
  assign po0740 = lo1283 ;
  assign po0741 = lo0917 ;
  assign po0742 = lo1060 ;
  assign po0743 = lo1056 ;
  assign po0744 = lo1057 ;
  assign po0745 = lo1059 ;
  assign po0746 = lo1058 ;
  assign po0747 = lo0019 ;
  assign po0748 = lo0020 ;
  assign po0749 = lo0040 ;
  assign po0750 = new_n1980 ;
  assign po0751 = pi000 ;
  assign po0752 = lo1283 ;
  assign po0753 = lo0917 ;
  assign po0754 = lo1060 ;
  assign po0755 = lo1056 ;
  assign po0756 = lo1057 ;
  assign po0757 = lo1059 ;
  assign po0758 = lo1058 ;
  assign po0759 = lo0019 ;
  assign po0760 = lo0020 ;
  assign po0761 = lo0040 ;
  assign po0762 = new_n1983 ;
  assign po0763 = pi000 ;
  assign po0764 = lo1283 ;
  assign po0765 = lo0917 ;
  assign po0766 = lo1060 ;
  assign po0767 = lo1056 ;
  assign po0768 = lo1057 ;
  assign po0769 = lo1059 ;
  assign po0770 = lo1058 ;
  assign po0771 = lo0019 ;
  assign po0772 = lo0020 ;
  assign po0773 = lo0040 ;
  assign po0774 = new_n1986 ;
  assign po0775 = pi000 ;
  assign po0776 = lo1283 ;
  assign po0777 = lo0917 ;
  assign po0778 = lo1060 ;
  assign po0779 = lo1056 ;
  assign po0780 = lo1057 ;
  assign po0781 = lo1059 ;
  assign po0782 = lo1058 ;
  assign po0783 = lo0019 ;
  assign po0784 = lo0020 ;
  assign po0785 = lo0040 ;
  assign po0786 = new_n1994 ;
  assign po0787 = pi000 ;
  assign po0788 = lo1423 ;
  assign po0789 = lo0917 ;
  assign po0790 = lo1060 ;
  assign po0791 = lo1056 ;
  assign po0792 = lo1057 ;
  assign po0793 = lo1059 ;
  assign po0794 = lo1058 ;
  assign po0795 = lo0019 ;
  assign po0796 = lo0020 ;
  assign po0797 = lo0040 ;
  assign po0798 = new_n1995 ;
  assign po0799 = pi000 ;
  assign po0800 = lo1423 ;
  assign po0801 = lo0917 ;
  assign po0802 = lo1060 ;
  assign po0803 = lo1056 ;
  assign po0804 = lo1057 ;
  assign po0805 = lo1059 ;
  assign po0806 = lo1058 ;
  assign po0807 = lo0019 ;
  assign po0808 = lo0020 ;
  assign po0809 = lo0040 ;
  assign po0810 = new_n1996 ;
  assign po0811 = pi000 ;
  assign po0812 = lo1423 ;
  assign po0813 = lo0917 ;
  assign po0814 = lo1060 ;
  assign po0815 = lo1056 ;
  assign po0816 = lo1057 ;
  assign po0817 = lo1059 ;
  assign po0818 = lo1058 ;
  assign po0819 = lo0019 ;
  assign po0820 = lo0020 ;
  assign po0821 = lo0040 ;
  assign po0822 = new_n1997 ;
  assign po0823 = pi000 ;
  assign po0824 = lo1423 ;
  assign po0825 = lo0917 ;
  assign po0826 = lo1060 ;
  assign po0827 = lo1056 ;
  assign po0828 = lo1057 ;
  assign po0829 = lo1059 ;
  assign po0830 = lo1058 ;
  assign po0831 = lo0019 ;
  assign po0832 = lo0020 ;
  assign po0833 = lo0040 ;
  assign po0834 = new_n1998 ;
  assign po0835 = pi000 ;
  assign po0836 = lo1423 ;
  assign po0837 = lo0917 ;
  assign po0838 = lo1060 ;
  assign po0839 = lo1056 ;
  assign po0840 = lo1057 ;
  assign po0841 = lo1059 ;
  assign po0842 = lo1058 ;
  assign po0843 = lo0019 ;
  assign po0844 = lo0020 ;
  assign po0845 = lo0040 ;
  assign po0846 = new_n1999 ;
  assign po0847 = pi000 ;
  assign po0848 = lo1423 ;
  assign po0849 = lo0917 ;
  assign po0850 = lo1060 ;
  assign po0851 = lo1056 ;
  assign po0852 = lo1057 ;
  assign po0853 = lo1059 ;
  assign po0854 = lo1058 ;
  assign po0855 = lo0019 ;
  assign po0856 = lo0020 ;
  assign po0857 = lo0040 ;
  assign po0858 = new_n2000 ;
  assign po0859 = pi000 ;
  assign po0860 = lo1423 ;
  assign po0861 = lo0917 ;
  assign po0862 = lo1060 ;
  assign po0863 = lo1056 ;
  assign po0864 = lo1057 ;
  assign po0865 = lo1059 ;
  assign po0866 = lo1058 ;
  assign po0867 = lo0019 ;
  assign po0868 = lo0020 ;
  assign po0869 = lo0040 ;
  assign po0870 = new_n2001 ;
  assign po0871 = pi000 ;
  assign po0872 = lo1423 ;
  assign po0873 = lo0917 ;
  assign po0874 = lo1060 ;
  assign po0875 = lo1056 ;
  assign po0876 = lo1057 ;
  assign po0877 = lo1059 ;
  assign po0878 = lo1058 ;
  assign po0879 = lo0019 ;
  assign po0880 = lo0020 ;
  assign po0881 = lo0040 ;
  assign po0882 = new_n2003 ;
  assign po0883 = pi000 ;
  assign po0884 = lo1055 ;
  assign po0885 = lo0917 ;
  assign po0886 = lo1060 ;
  assign po0887 = lo1056 ;
  assign po0888 = lo1057 ;
  assign po0889 = lo1059 ;
  assign po0890 = lo1058 ;
  assign po0891 = lo0019 ;
  assign po0892 = lo0020 ;
  assign po0893 = lo0040 ;
  assign po0894 = new_n2004 ;
  assign po0895 = pi000 ;
  assign po0896 = lo1055 ;
  assign po0897 = lo0917 ;
  assign po0898 = lo1060 ;
  assign po0899 = lo1056 ;
  assign po0900 = lo1057 ;
  assign po0901 = lo1059 ;
  assign po0902 = lo1058 ;
  assign po0903 = lo0019 ;
  assign po0904 = lo0020 ;
  assign po0905 = lo0040 ;
  assign po0906 = new_n2005 ;
  assign po0907 = pi000 ;
  assign po0908 = lo1055 ;
  assign po0909 = lo0917 ;
  assign po0910 = lo1060 ;
  assign po0911 = lo1056 ;
  assign po0912 = lo1057 ;
  assign po0913 = lo1059 ;
  assign po0914 = lo1058 ;
  assign po0915 = lo0019 ;
  assign po0916 = lo0020 ;
  assign po0917 = lo0040 ;
  assign po0918 = new_n2006 ;
  assign po0919 = pi000 ;
  assign po0920 = lo1055 ;
  assign po0921 = lo0917 ;
  assign po0922 = lo1060 ;
  assign po0923 = lo1056 ;
  assign po0924 = lo1057 ;
  assign po0925 = lo1059 ;
  assign po0926 = lo1058 ;
  assign po0927 = lo0019 ;
  assign po0928 = lo0020 ;
  assign po0929 = lo0040 ;
  assign po0930 = new_n2007 ;
  assign po0931 = pi000 ;
  assign po0932 = lo1055 ;
  assign po0933 = lo0917 ;
  assign po0934 = lo1060 ;
  assign po0935 = lo1056 ;
  assign po0936 = lo1057 ;
  assign po0937 = lo1059 ;
  assign po0938 = lo1058 ;
  assign po0939 = lo0019 ;
  assign po0940 = lo0020 ;
  assign po0941 = lo0040 ;
  assign po0942 = new_n2008 ;
  assign po0943 = pi000 ;
  assign po0944 = lo1055 ;
  assign po0945 = lo0917 ;
  assign po0946 = lo1060 ;
  assign po0947 = lo1056 ;
  assign po0948 = lo1057 ;
  assign po0949 = lo1059 ;
  assign po0950 = lo1058 ;
  assign po0951 = lo0019 ;
  assign po0952 = lo0020 ;
  assign po0953 = lo0040 ;
  assign po0954 = new_n2009 ;
  assign po0955 = pi000 ;
  assign po0956 = lo1055 ;
  assign po0957 = lo0917 ;
  assign po0958 = lo1060 ;
  assign po0959 = lo1056 ;
  assign po0960 = lo1057 ;
  assign po0961 = lo1059 ;
  assign po0962 = lo1058 ;
  assign po0963 = lo0019 ;
  assign po0964 = lo0020 ;
  assign po0965 = lo0040 ;
  assign po0966 = new_n2010 ;
  assign po0967 = pi000 ;
  assign po0968 = lo1055 ;
  assign po0969 = lo0917 ;
  assign po0970 = lo1060 ;
  assign po0971 = lo1056 ;
  assign po0972 = lo1057 ;
  assign po0973 = lo1059 ;
  assign po0974 = lo1058 ;
  assign po0975 = lo0019 ;
  assign po0976 = lo0020 ;
  assign po0977 = lo0040 ;
  assign po0978 = new_n1994 ;
  assign po0979 = pi000 ;
  assign po0980 = lo1270 ;
  assign po0981 = lo0917 ;
  assign po0982 = lo1060 ;
  assign po0983 = lo1056 ;
  assign po0984 = lo1057 ;
  assign po0985 = lo1059 ;
  assign po0986 = lo1058 ;
  assign po0987 = lo0019 ;
  assign po0988 = lo0020 ;
  assign po0989 = lo0040 ;
  assign po0990 = new_n1999 ;
  assign po0991 = pi000 ;
  assign po0992 = lo1270 ;
  assign po0993 = lo0917 ;
  assign po0994 = lo1060 ;
  assign po0995 = lo1056 ;
  assign po0996 = lo1057 ;
  assign po0997 = lo1059 ;
  assign po0998 = lo1058 ;
  assign po0999 = lo0019 ;
  assign po1000 = lo0020 ;
  assign po1001 = lo0040 ;
  assign po1002 = new_n1995 ;
  assign po1003 = pi000 ;
  assign po1004 = lo1270 ;
  assign po1005 = lo0917 ;
  assign po1006 = lo1060 ;
  assign po1007 = lo1056 ;
  assign po1008 = lo1057 ;
  assign po1009 = lo1059 ;
  assign po1010 = lo1058 ;
  assign po1011 = lo0019 ;
  assign po1012 = lo0020 ;
  assign po1013 = lo0040 ;
  assign po1014 = new_n2000 ;
  assign po1015 = pi000 ;
  assign po1016 = lo1270 ;
  assign po1017 = lo0917 ;
  assign po1018 = lo1060 ;
  assign po1019 = lo1056 ;
  assign po1020 = lo1057 ;
  assign po1021 = lo1059 ;
  assign po1022 = lo1058 ;
  assign po1023 = lo0019 ;
  assign po1024 = lo0020 ;
  assign po1025 = lo0040 ;
  assign po1026 = new_n1998 ;
  assign po1027 = pi000 ;
  assign po1028 = lo1270 ;
  assign po1029 = lo0917 ;
  assign po1030 = lo1060 ;
  assign po1031 = lo1056 ;
  assign po1032 = lo1057 ;
  assign po1033 = lo1059 ;
  assign po1034 = lo1058 ;
  assign po1035 = lo0019 ;
  assign po1036 = lo0020 ;
  assign po1037 = lo0040 ;
  assign po1038 = new_n1996 ;
  assign po1039 = pi000 ;
  assign po1040 = lo1270 ;
  assign po1041 = lo0917 ;
  assign po1042 = lo1060 ;
  assign po1043 = lo1056 ;
  assign po1044 = lo1057 ;
  assign po1045 = lo1059 ;
  assign po1046 = lo1058 ;
  assign po1047 = lo0019 ;
  assign po1048 = lo0020 ;
  assign po1049 = lo0040 ;
  assign po1050 = new_n1997 ;
  assign po1051 = pi000 ;
  assign po1052 = lo1270 ;
  assign po1053 = lo0917 ;
  assign po1054 = lo1060 ;
  assign po1055 = lo1056 ;
  assign po1056 = lo1057 ;
  assign po1057 = lo1059 ;
  assign po1058 = lo1058 ;
  assign po1059 = lo0019 ;
  assign po1060 = lo0020 ;
  assign po1061 = lo0040 ;
  assign po1062 = new_n2001 ;
  assign po1063 = pi000 ;
  assign po1064 = lo1270 ;
  assign po1065 = lo0917 ;
  assign po1066 = lo1060 ;
  assign po1067 = lo1056 ;
  assign po1068 = lo1057 ;
  assign po1069 = lo1059 ;
  assign po1070 = lo1058 ;
  assign po1071 = lo0019 ;
  assign po1072 = lo0020 ;
  assign po1073 = lo0040 ;
  assign po1074 = new_n2009 ;
  assign po1075 = pi000 ;
  assign po1076 = lo1093 ;
  assign po1077 = lo0917 ;
  assign po1078 = lo1060 ;
  assign po1079 = lo1056 ;
  assign po1080 = lo1057 ;
  assign po1081 = lo1059 ;
  assign po1082 = lo1058 ;
  assign po1083 = lo0019 ;
  assign po1084 = lo0020 ;
  assign po1085 = lo0040 ;
  assign po1086 = new_n2005 ;
  assign po1087 = pi000 ;
  assign po1088 = lo1093 ;
  assign po1089 = lo0917 ;
  assign po1090 = lo1060 ;
  assign po1091 = lo1056 ;
  assign po1092 = lo1057 ;
  assign po1093 = lo1059 ;
  assign po1094 = lo1058 ;
  assign po1095 = lo0019 ;
  assign po1096 = lo0020 ;
  assign po1097 = lo0040 ;
  assign po1098 = new_n2006 ;
  assign po1099 = pi000 ;
  assign po1100 = lo1093 ;
  assign po1101 = lo0917 ;
  assign po1102 = lo1060 ;
  assign po1103 = lo1056 ;
  assign po1104 = lo1057 ;
  assign po1105 = lo1059 ;
  assign po1106 = lo1058 ;
  assign po1107 = lo0019 ;
  assign po1108 = lo0020 ;
  assign po1109 = lo0040 ;
  assign po1110 = new_n2007 ;
  assign po1111 = pi000 ;
  assign po1112 = lo1093 ;
  assign po1113 = lo0917 ;
  assign po1114 = lo1060 ;
  assign po1115 = lo1056 ;
  assign po1116 = lo1057 ;
  assign po1117 = lo1059 ;
  assign po1118 = lo1058 ;
  assign po1119 = lo0019 ;
  assign po1120 = lo0020 ;
  assign po1121 = lo0040 ;
  assign po1122 = new_n2008 ;
  assign po1123 = pi000 ;
  assign po1124 = lo1093 ;
  assign po1125 = lo0917 ;
  assign po1126 = lo1060 ;
  assign po1127 = lo1056 ;
  assign po1128 = lo1057 ;
  assign po1129 = lo1059 ;
  assign po1130 = lo1058 ;
  assign po1131 = lo0019 ;
  assign po1132 = lo0020 ;
  assign po1133 = lo0040 ;
  assign po1134 = new_n2003 ;
  assign po1135 = pi000 ;
  assign po1136 = lo1093 ;
  assign po1137 = lo0917 ;
  assign po1138 = lo1060 ;
  assign po1139 = lo1056 ;
  assign po1140 = lo1057 ;
  assign po1141 = lo1059 ;
  assign po1142 = lo1058 ;
  assign po1143 = lo0019 ;
  assign po1144 = lo0020 ;
  assign po1145 = lo0040 ;
  assign po1146 = new_n2004 ;
  assign po1147 = pi000 ;
  assign po1148 = lo1093 ;
  assign po1149 = lo0917 ;
  assign po1150 = lo1060 ;
  assign po1151 = lo1056 ;
  assign po1152 = lo1057 ;
  assign po1153 = lo1059 ;
  assign po1154 = lo1058 ;
  assign po1155 = lo0019 ;
  assign po1156 = lo0020 ;
  assign po1157 = lo0040 ;
  assign po1158 = new_n2010 ;
  assign po1159 = pi000 ;
  assign po1160 = lo1093 ;
  assign po1161 = lo0917 ;
  assign po1162 = lo1060 ;
  assign po1163 = lo1056 ;
  assign po1164 = lo1057 ;
  assign po1165 = lo1059 ;
  assign po1166 = lo1058 ;
  assign po1167 = lo0019 ;
  assign po1168 = lo0020 ;
  assign po1169 = lo0040 ;
  assign po1170 = new_n1994 ;
  assign po1171 = pi000 ;
  assign po1172 = lo1420 ;
  assign po1173 = lo0917 ;
  assign po1174 = lo1060 ;
  assign po1175 = lo1056 ;
  assign po1176 = lo1057 ;
  assign po1177 = lo1059 ;
  assign po1178 = lo1058 ;
  assign po1179 = lo0019 ;
  assign po1180 = lo0020 ;
  assign po1181 = lo0040 ;
  assign po1182 = new_n1995 ;
  assign po1183 = pi000 ;
  assign po1184 = lo1420 ;
  assign po1185 = lo0917 ;
  assign po1186 = lo1060 ;
  assign po1187 = lo1056 ;
  assign po1188 = lo1057 ;
  assign po1189 = lo1059 ;
  assign po1190 = lo1058 ;
  assign po1191 = lo0019 ;
  assign po1192 = lo0020 ;
  assign po1193 = lo0040 ;
  assign po1194 = new_n1996 ;
  assign po1195 = pi000 ;
  assign po1196 = lo1420 ;
  assign po1197 = lo0917 ;
  assign po1198 = lo1060 ;
  assign po1199 = lo1056 ;
  assign po1200 = lo1057 ;
  assign po1201 = lo1059 ;
  assign po1202 = lo1058 ;
  assign po1203 = lo0019 ;
  assign po1204 = lo0020 ;
  assign po1205 = lo0040 ;
  assign po1206 = new_n1997 ;
  assign po1207 = pi000 ;
  assign po1208 = lo1420 ;
  assign po1209 = lo0917 ;
  assign po1210 = lo1060 ;
  assign po1211 = lo1056 ;
  assign po1212 = lo1057 ;
  assign po1213 = lo1059 ;
  assign po1214 = lo1058 ;
  assign po1215 = lo0019 ;
  assign po1216 = lo0020 ;
  assign po1217 = lo0040 ;
  assign po1218 = new_n1998 ;
  assign po1219 = pi000 ;
  assign po1220 = lo1420 ;
  assign po1221 = lo0917 ;
  assign po1222 = lo1060 ;
  assign po1223 = lo1056 ;
  assign po1224 = lo1057 ;
  assign po1225 = lo1059 ;
  assign po1226 = lo1058 ;
  assign po1227 = lo0019 ;
  assign po1228 = lo0020 ;
  assign po1229 = lo0040 ;
  assign po1230 = new_n1999 ;
  assign po1231 = pi000 ;
  assign po1232 = lo1420 ;
  assign po1233 = lo0917 ;
  assign po1234 = lo1060 ;
  assign po1235 = lo1056 ;
  assign po1236 = lo1057 ;
  assign po1237 = lo1059 ;
  assign po1238 = lo1058 ;
  assign po1239 = lo0019 ;
  assign po1240 = lo0020 ;
  assign po1241 = lo0040 ;
  assign po1242 = new_n2000 ;
  assign po1243 = pi000 ;
  assign po1244 = lo1420 ;
  assign po1245 = lo0917 ;
  assign po1246 = lo1060 ;
  assign po1247 = lo1056 ;
  assign po1248 = lo1057 ;
  assign po1249 = lo1059 ;
  assign po1250 = lo1058 ;
  assign po1251 = lo0019 ;
  assign po1252 = lo0020 ;
  assign po1253 = lo0040 ;
  assign po1254 = new_n2001 ;
  assign po1255 = pi000 ;
  assign po1256 = lo1420 ;
  assign po1257 = lo0917 ;
  assign po1258 = lo1060 ;
  assign po1259 = lo1056 ;
  assign po1260 = lo1057 ;
  assign po1261 = lo1059 ;
  assign po1262 = lo1058 ;
  assign po1263 = lo0019 ;
  assign po1264 = lo0020 ;
  assign po1265 = lo0040 ;
  assign po1266 = new_n2003 ;
  assign po1267 = pi000 ;
  assign po1268 = lo1053 ;
  assign po1269 = lo0917 ;
  assign po1270 = lo1060 ;
  assign po1271 = lo1056 ;
  assign po1272 = lo1057 ;
  assign po1273 = lo1059 ;
  assign po1274 = lo1058 ;
  assign po1275 = lo0019 ;
  assign po1276 = lo0020 ;
  assign po1277 = lo0040 ;
  assign po1278 = new_n2004 ;
  assign po1279 = pi000 ;
  assign po1280 = lo1053 ;
  assign po1281 = lo0917 ;
  assign po1282 = lo1060 ;
  assign po1283 = lo1056 ;
  assign po1284 = lo1057 ;
  assign po1285 = lo1059 ;
  assign po1286 = lo1058 ;
  assign po1287 = lo0019 ;
  assign po1288 = lo0020 ;
  assign po1289 = lo0040 ;
  assign po1290 = new_n2005 ;
  assign po1291 = pi000 ;
  assign po1292 = lo1053 ;
  assign po1293 = lo0917 ;
  assign po1294 = lo1060 ;
  assign po1295 = lo1056 ;
  assign po1296 = lo1057 ;
  assign po1297 = lo1059 ;
  assign po1298 = lo1058 ;
  assign po1299 = lo0019 ;
  assign po1300 = lo0020 ;
  assign po1301 = lo0040 ;
  assign po1302 = new_n2006 ;
  assign po1303 = pi000 ;
  assign po1304 = lo1053 ;
  assign po1305 = lo0917 ;
  assign po1306 = lo1060 ;
  assign po1307 = lo1056 ;
  assign po1308 = lo1057 ;
  assign po1309 = lo1059 ;
  assign po1310 = lo1058 ;
  assign po1311 = lo0019 ;
  assign po1312 = lo0020 ;
  assign po1313 = lo0040 ;
  assign po1314 = new_n2007 ;
  assign po1315 = pi000 ;
  assign po1316 = lo1053 ;
  assign po1317 = lo0917 ;
  assign po1318 = lo1060 ;
  assign po1319 = lo1056 ;
  assign po1320 = lo1057 ;
  assign po1321 = lo1059 ;
  assign po1322 = lo1058 ;
  assign po1323 = lo0019 ;
  assign po1324 = lo0020 ;
  assign po1325 = lo0040 ;
  assign po1326 = new_n2008 ;
  assign po1327 = pi000 ;
  assign po1328 = lo1053 ;
  assign po1329 = lo0917 ;
  assign po1330 = lo1060 ;
  assign po1331 = lo1056 ;
  assign po1332 = lo1057 ;
  assign po1333 = lo1059 ;
  assign po1334 = lo1058 ;
  assign po1335 = lo0019 ;
  assign po1336 = lo0020 ;
  assign po1337 = lo0040 ;
  assign po1338 = new_n2009 ;
  assign po1339 = pi000 ;
  assign po1340 = lo1053 ;
  assign po1341 = lo0917 ;
  assign po1342 = lo1060 ;
  assign po1343 = lo1056 ;
  assign po1344 = lo1057 ;
  assign po1345 = lo1059 ;
  assign po1346 = lo1058 ;
  assign po1347 = lo0019 ;
  assign po1348 = lo0020 ;
  assign po1349 = lo0040 ;
  assign po1350 = new_n2010 ;
  assign po1351 = pi000 ;
  assign po1352 = lo1053 ;
  assign po1353 = lo0917 ;
  assign po1354 = lo1060 ;
  assign po1355 = lo1056 ;
  assign po1356 = lo1057 ;
  assign po1357 = lo1059 ;
  assign po1358 = lo1058 ;
  assign po1359 = lo0019 ;
  assign po1360 = lo0020 ;
  assign po1361 = lo0040 ;
  assign po1362 = new_n1994 ;
  assign po1363 = pi000 ;
  assign po1364 = lo1271 ;
  assign po1365 = lo0917 ;
  assign po1366 = lo1060 ;
  assign po1367 = lo1056 ;
  assign po1368 = lo1057 ;
  assign po1369 = lo1059 ;
  assign po1370 = lo1058 ;
  assign po1371 = lo0019 ;
  assign po1372 = lo0020 ;
  assign po1373 = lo0040 ;
  assign po1374 = new_n1995 ;
  assign po1375 = pi000 ;
  assign po1376 = lo1271 ;
  assign po1377 = lo0917 ;
  assign po1378 = lo1060 ;
  assign po1379 = lo1056 ;
  assign po1380 = lo1057 ;
  assign po1381 = lo1059 ;
  assign po1382 = lo1058 ;
  assign po1383 = lo0019 ;
  assign po1384 = lo0020 ;
  assign po1385 = lo0040 ;
  assign po1386 = new_n1996 ;
  assign po1387 = pi000 ;
  assign po1388 = lo1271 ;
  assign po1389 = lo0917 ;
  assign po1390 = lo1060 ;
  assign po1391 = lo1056 ;
  assign po1392 = lo1057 ;
  assign po1393 = lo1059 ;
  assign po1394 = lo1058 ;
  assign po1395 = lo0019 ;
  assign po1396 = lo0020 ;
  assign po1397 = lo0040 ;
  assign po1398 = new_n1997 ;
  assign po1399 = pi000 ;
  assign po1400 = lo1271 ;
  assign po1401 = lo0917 ;
  assign po1402 = lo1060 ;
  assign po1403 = lo1056 ;
  assign po1404 = lo1057 ;
  assign po1405 = lo1059 ;
  assign po1406 = lo1058 ;
  assign po1407 = lo0019 ;
  assign po1408 = lo0020 ;
  assign po1409 = lo0040 ;
  assign po1410 = new_n1998 ;
  assign po1411 = pi000 ;
  assign po1412 = lo1271 ;
  assign po1413 = lo0917 ;
  assign po1414 = lo1060 ;
  assign po1415 = lo1056 ;
  assign po1416 = lo1057 ;
  assign po1417 = lo1059 ;
  assign po1418 = lo1058 ;
  assign po1419 = lo0019 ;
  assign po1420 = lo0020 ;
  assign po1421 = lo0040 ;
  assign po1422 = new_n1999 ;
  assign po1423 = pi000 ;
  assign po1424 = lo1271 ;
  assign po1425 = lo0917 ;
  assign po1426 = lo1060 ;
  assign po1427 = lo1056 ;
  assign po1428 = lo1057 ;
  assign po1429 = lo1059 ;
  assign po1430 = lo1058 ;
  assign po1431 = lo0019 ;
  assign po1432 = lo0020 ;
  assign po1433 = lo0040 ;
  assign po1434 = new_n2000 ;
  assign po1435 = pi000 ;
  assign po1436 = lo1271 ;
  assign po1437 = lo0917 ;
  assign po1438 = lo1060 ;
  assign po1439 = lo1056 ;
  assign po1440 = lo1057 ;
  assign po1441 = lo1059 ;
  assign po1442 = lo1058 ;
  assign po1443 = lo0019 ;
  assign po1444 = lo0020 ;
  assign po1445 = lo0040 ;
  assign po1446 = new_n2001 ;
  assign po1447 = pi000 ;
  assign po1448 = lo1271 ;
  assign po1449 = lo0917 ;
  assign po1450 = lo1060 ;
  assign po1451 = lo1056 ;
  assign po1452 = lo1057 ;
  assign po1453 = lo1059 ;
  assign po1454 = lo1058 ;
  assign po1455 = lo0019 ;
  assign po1456 = lo0020 ;
  assign po1457 = lo0040 ;
  assign po1458 = new_n2003 ;
  assign po1459 = pi000 ;
  assign po1460 = lo1094 ;
  assign po1461 = lo0917 ;
  assign po1462 = lo1060 ;
  assign po1463 = lo1056 ;
  assign po1464 = lo1057 ;
  assign po1465 = lo1059 ;
  assign po1466 = lo1058 ;
  assign po1467 = lo0019 ;
  assign po1468 = lo0020 ;
  assign po1469 = lo0040 ;
  assign po1470 = new_n2004 ;
  assign po1471 = pi000 ;
  assign po1472 = lo1094 ;
  assign po1473 = lo0917 ;
  assign po1474 = lo1060 ;
  assign po1475 = lo1056 ;
  assign po1476 = lo1057 ;
  assign po1477 = lo1059 ;
  assign po1478 = lo1058 ;
  assign po1479 = lo0019 ;
  assign po1480 = lo0020 ;
  assign po1481 = lo0040 ;
  assign po1482 = new_n2005 ;
  assign po1483 = pi000 ;
  assign po1484 = lo1094 ;
  assign po1485 = lo0917 ;
  assign po1486 = lo1060 ;
  assign po1487 = lo1056 ;
  assign po1488 = lo1057 ;
  assign po1489 = lo1059 ;
  assign po1490 = lo1058 ;
  assign po1491 = lo0019 ;
  assign po1492 = lo0020 ;
  assign po1493 = lo0040 ;
  assign po1494 = new_n2006 ;
  assign po1495 = pi000 ;
  assign po1496 = lo1094 ;
  assign po1497 = lo0917 ;
  assign po1498 = lo1060 ;
  assign po1499 = lo1056 ;
  assign po1500 = lo1057 ;
  assign po1501 = lo1059 ;
  assign po1502 = lo1058 ;
  assign po1503 = lo0019 ;
  assign po1504 = lo0020 ;
  assign po1505 = lo0040 ;
  assign po1506 = new_n2007 ;
  assign po1507 = pi000 ;
  assign po1508 = lo1094 ;
  assign po1509 = lo0917 ;
  assign po1510 = lo1060 ;
  assign po1511 = lo1056 ;
  assign po1512 = lo1057 ;
  assign po1513 = lo1059 ;
  assign po1514 = lo1058 ;
  assign po1515 = lo0019 ;
  assign po1516 = lo0020 ;
  assign po1517 = lo0040 ;
  assign po1518 = new_n2008 ;
  assign po1519 = pi000 ;
  assign po1520 = lo1094 ;
  assign po1521 = lo0917 ;
  assign po1522 = lo1060 ;
  assign po1523 = lo1056 ;
  assign po1524 = lo1057 ;
  assign po1525 = lo1059 ;
  assign po1526 = lo1058 ;
  assign po1527 = lo0019 ;
  assign po1528 = lo0020 ;
  assign po1529 = lo0040 ;
  assign po1530 = new_n2009 ;
  assign po1531 = pi000 ;
  assign po1532 = lo1094 ;
  assign po1533 = lo0917 ;
  assign po1534 = lo1060 ;
  assign po1535 = lo1056 ;
  assign po1536 = lo1057 ;
  assign po1537 = lo1059 ;
  assign po1538 = lo1058 ;
  assign po1539 = lo0019 ;
  assign po1540 = lo0020 ;
  assign po1541 = lo0040 ;
  assign po1542 = new_n2010 ;
  assign po1543 = pi000 ;
  assign po1544 = lo1094 ;
  assign po1545 = lo0917 ;
  assign po1546 = lo1060 ;
  assign po1547 = lo1056 ;
  assign po1548 = lo1057 ;
  assign po1549 = lo1059 ;
  assign po1550 = lo1058 ;
  assign po1551 = lo0019 ;
  assign po1552 = lo0020 ;
  assign po1553 = lo0040 ;
  assign po1554 = new_n2012 ;
  assign po1555 = pi000 ;
  assign po1556 = lo1277 ;
  assign po1557 = lo0917 ;
  assign po1558 = lo1060 ;
  assign po1559 = lo1056 ;
  assign po1560 = lo1057 ;
  assign po1561 = lo1059 ;
  assign po1562 = lo1058 ;
  assign po1563 = lo0019 ;
  assign po1564 = lo0020 ;
  assign po1565 = lo0040 ;
  assign po1566 = new_n2013 ;
  assign po1567 = pi000 ;
  assign po1568 = lo1277 ;
  assign po1569 = lo0917 ;
  assign po1570 = lo1060 ;
  assign po1571 = lo1056 ;
  assign po1572 = lo1057 ;
  assign po1573 = lo1059 ;
  assign po1574 = lo1058 ;
  assign po1575 = lo0019 ;
  assign po1576 = lo0020 ;
  assign po1577 = lo0040 ;
  assign po1578 = new_n2014 ;
  assign po1579 = pi000 ;
  assign po1580 = lo1277 ;
  assign po1581 = lo0917 ;
  assign po1582 = lo1060 ;
  assign po1583 = lo1056 ;
  assign po1584 = lo1057 ;
  assign po1585 = lo1059 ;
  assign po1586 = lo1058 ;
  assign po1587 = lo0019 ;
  assign po1588 = lo0020 ;
  assign po1589 = lo0040 ;
  assign po1590 = new_n2015 ;
  assign po1591 = pi000 ;
  assign po1592 = lo1277 ;
  assign po1593 = lo0917 ;
  assign po1594 = lo1060 ;
  assign po1595 = lo1056 ;
  assign po1596 = lo1057 ;
  assign po1597 = lo1059 ;
  assign po1598 = lo1058 ;
  assign po1599 = lo0019 ;
  assign po1600 = lo0020 ;
  assign po1601 = lo0040 ;
  assign po1602 = new_n2016 ;
  assign po1603 = pi000 ;
  assign po1604 = lo1277 ;
  assign po1605 = lo0917 ;
  assign po1606 = lo1060 ;
  assign po1607 = lo1056 ;
  assign po1608 = lo1057 ;
  assign po1609 = lo1059 ;
  assign po1610 = lo1058 ;
  assign po1611 = lo0019 ;
  assign po1612 = lo0020 ;
  assign po1613 = lo0040 ;
  assign po1614 = new_n2017 ;
  assign po1615 = pi000 ;
  assign po1616 = lo1277 ;
  assign po1617 = lo0917 ;
  assign po1618 = lo1060 ;
  assign po1619 = lo1056 ;
  assign po1620 = lo1057 ;
  assign po1621 = lo1059 ;
  assign po1622 = lo1058 ;
  assign po1623 = lo0019 ;
  assign po1624 = lo0020 ;
  assign po1625 = lo0040 ;
  assign po1626 = new_n2018 ;
  assign po1627 = pi000 ;
  assign po1628 = lo1277 ;
  assign po1629 = lo0917 ;
  assign po1630 = lo1060 ;
  assign po1631 = lo1056 ;
  assign po1632 = lo1057 ;
  assign po1633 = lo1059 ;
  assign po1634 = lo1058 ;
  assign po1635 = lo0019 ;
  assign po1636 = lo0020 ;
  assign po1637 = lo0040 ;
  assign po1638 = new_n2019 ;
  assign po1639 = pi000 ;
  assign po1640 = lo1277 ;
  assign po1641 = lo0917 ;
  assign po1642 = lo1060 ;
  assign po1643 = lo1056 ;
  assign po1644 = lo1057 ;
  assign po1645 = lo1059 ;
  assign po1646 = lo1058 ;
  assign po1647 = lo0019 ;
  assign po1648 = lo0020 ;
  assign po1649 = lo0040 ;
  assign po1650 = new_n1974 ;
  assign po1651 = pi000 ;
  assign po1652 = lo1446 ;
  assign po1653 = lo0917 ;
  assign po1654 = lo1060 ;
  assign po1655 = lo1056 ;
  assign po1656 = lo1057 ;
  assign po1657 = lo1059 ;
  assign po1658 = lo1058 ;
  assign po1659 = lo0019 ;
  assign po1660 = lo0020 ;
  assign po1661 = lo0040 ;
  assign po1662 = new_n1977 ;
  assign po1663 = pi000 ;
  assign po1664 = lo1446 ;
  assign po1665 = lo0917 ;
  assign po1666 = lo1060 ;
  assign po1667 = lo1056 ;
  assign po1668 = lo1057 ;
  assign po1669 = lo1059 ;
  assign po1670 = lo1058 ;
  assign po1671 = lo0019 ;
  assign po1672 = lo0020 ;
  assign po1673 = lo0040 ;
  assign po1674 = new_n1980 ;
  assign po1675 = pi000 ;
  assign po1676 = lo1446 ;
  assign po1677 = lo0917 ;
  assign po1678 = lo1060 ;
  assign po1679 = lo1056 ;
  assign po1680 = lo1057 ;
  assign po1681 = lo1059 ;
  assign po1682 = lo1058 ;
  assign po1683 = lo0019 ;
  assign po1684 = lo0020 ;
  assign po1685 = lo0040 ;
  assign po1686 = new_n1983 ;
  assign po1687 = pi000 ;
  assign po1688 = lo1446 ;
  assign po1689 = lo0917 ;
  assign po1690 = lo1060 ;
  assign po1691 = lo1056 ;
  assign po1692 = lo1057 ;
  assign po1693 = lo1059 ;
  assign po1694 = lo1058 ;
  assign po1695 = lo0019 ;
  assign po1696 = lo0020 ;
  assign po1697 = lo0040 ;
  assign po1698 = new_n1986 ;
  assign po1699 = pi000 ;
  assign po1700 = lo1446 ;
  assign po1701 = lo0917 ;
  assign po1702 = lo1060 ;
  assign po1703 = lo1056 ;
  assign po1704 = lo1057 ;
  assign po1705 = lo1059 ;
  assign po1706 = lo1058 ;
  assign po1707 = lo0019 ;
  assign po1708 = lo0020 ;
  assign po1709 = lo0040 ;
  assign po1710 = new_n1988 ;
  assign po1711 = pi000 ;
  assign po1712 = lo1446 ;
  assign po1713 = lo0917 ;
  assign po1714 = lo1060 ;
  assign po1715 = lo1056 ;
  assign po1716 = lo1057 ;
  assign po1717 = lo1059 ;
  assign po1718 = lo1058 ;
  assign po1719 = lo0019 ;
  assign po1720 = lo0020 ;
  assign po1721 = lo0040 ;
  assign po1722 = new_n1990 ;
  assign po1723 = pi000 ;
  assign po1724 = lo1446 ;
  assign po1725 = lo0917 ;
  assign po1726 = lo1060 ;
  assign po1727 = lo1056 ;
  assign po1728 = lo1057 ;
  assign po1729 = lo1059 ;
  assign po1730 = lo1058 ;
  assign po1731 = lo0019 ;
  assign po1732 = lo0020 ;
  assign po1733 = lo0040 ;
  assign po1734 = new_n1992 ;
  assign po1735 = pi000 ;
  assign po1736 = lo1446 ;
  assign po1737 = lo0917 ;
  assign po1738 = lo1060 ;
  assign po1739 = lo1056 ;
  assign po1740 = lo1057 ;
  assign po1741 = lo1059 ;
  assign po1742 = lo1058 ;
  assign po1743 = lo0019 ;
  assign po1744 = lo0020 ;
  assign po1745 = lo0040 ;
  assign po1746 = new_n2012 ;
  assign po1747 = pi000 ;
  assign po1748 = lo1274 ;
  assign po1749 = lo0917 ;
  assign po1750 = lo1060 ;
  assign po1751 = lo1056 ;
  assign po1752 = lo1057 ;
  assign po1753 = lo1059 ;
  assign po1754 = lo1058 ;
  assign po1755 = lo0019 ;
  assign po1756 = lo0020 ;
  assign po1757 = lo0040 ;
  assign po1758 = new_n2013 ;
  assign po1759 = pi000 ;
  assign po1760 = lo1274 ;
  assign po1761 = lo0917 ;
  assign po1762 = lo1060 ;
  assign po1763 = lo1056 ;
  assign po1764 = lo1057 ;
  assign po1765 = lo1059 ;
  assign po1766 = lo1058 ;
  assign po1767 = lo0019 ;
  assign po1768 = lo0020 ;
  assign po1769 = lo0040 ;
  assign po1770 = new_n2014 ;
  assign po1771 = pi000 ;
  assign po1772 = lo1274 ;
  assign po1773 = lo0917 ;
  assign po1774 = lo1060 ;
  assign po1775 = lo1056 ;
  assign po1776 = lo1057 ;
  assign po1777 = lo1059 ;
  assign po1778 = lo1058 ;
  assign po1779 = lo0019 ;
  assign po1780 = lo0020 ;
  assign po1781 = lo0040 ;
  assign po1782 = new_n2015 ;
  assign po1783 = pi000 ;
  assign po1784 = lo1274 ;
  assign po1785 = lo0917 ;
  assign po1786 = lo1060 ;
  assign po1787 = lo1056 ;
  assign po1788 = lo1057 ;
  assign po1789 = lo1059 ;
  assign po1790 = lo1058 ;
  assign po1791 = lo0019 ;
  assign po1792 = lo0020 ;
  assign po1793 = lo0040 ;
  assign po1794 = new_n2016 ;
  assign po1795 = pi000 ;
  assign po1796 = lo1274 ;
  assign po1797 = lo0917 ;
  assign po1798 = lo1060 ;
  assign po1799 = lo1056 ;
  assign po1800 = lo1057 ;
  assign po1801 = lo1059 ;
  assign po1802 = lo1058 ;
  assign po1803 = lo0019 ;
  assign po1804 = lo0020 ;
  assign po1805 = lo0040 ;
  assign po1806 = new_n2017 ;
  assign po1807 = pi000 ;
  assign po1808 = lo1274 ;
  assign po1809 = lo0917 ;
  assign po1810 = lo1060 ;
  assign po1811 = lo1056 ;
  assign po1812 = lo1057 ;
  assign po1813 = lo1059 ;
  assign po1814 = lo1058 ;
  assign po1815 = lo0019 ;
  assign po1816 = lo0020 ;
  assign po1817 = lo0040 ;
  assign po1818 = new_n2018 ;
  assign po1819 = pi000 ;
  assign po1820 = lo1274 ;
  assign po1821 = lo0917 ;
  assign po1822 = lo1060 ;
  assign po1823 = lo1056 ;
  assign po1824 = lo1057 ;
  assign po1825 = lo1059 ;
  assign po1826 = lo1058 ;
  assign po1827 = lo0019 ;
  assign po1828 = lo0020 ;
  assign po1829 = lo0040 ;
  assign po1830 = new_n2019 ;
  assign po1831 = pi000 ;
  assign po1832 = lo1274 ;
  assign po1833 = lo0917 ;
  assign po1834 = lo1060 ;
  assign po1835 = lo1056 ;
  assign po1836 = lo1057 ;
  assign po1837 = lo1059 ;
  assign po1838 = lo1058 ;
  assign po1839 = lo0019 ;
  assign po1840 = lo0020 ;
  assign po1841 = lo0040 ;
  assign po1842 = new_n1988 ;
  assign po1843 = pi000 ;
  assign po1844 = lo1282 ;
  assign po1845 = lo0917 ;
  assign po1846 = lo1060 ;
  assign po1847 = lo1056 ;
  assign po1848 = lo1057 ;
  assign po1849 = lo1059 ;
  assign po1850 = lo1058 ;
  assign po1851 = lo0019 ;
  assign po1852 = lo0020 ;
  assign po1853 = lo0040 ;
  assign po1854 = new_n1992 ;
  assign po1855 = pi000 ;
  assign po1856 = lo1282 ;
  assign po1857 = lo0917 ;
  assign po1858 = lo1060 ;
  assign po1859 = lo1056 ;
  assign po1860 = lo1057 ;
  assign po1861 = lo1059 ;
  assign po1862 = lo1058 ;
  assign po1863 = lo0019 ;
  assign po1864 = lo0020 ;
  assign po1865 = lo0040 ;
  assign po1866 = new_n1990 ;
  assign po1867 = pi000 ;
  assign po1868 = lo1282 ;
  assign po1869 = lo0917 ;
  assign po1870 = lo1060 ;
  assign po1871 = lo1056 ;
  assign po1872 = lo1057 ;
  assign po1873 = lo1059 ;
  assign po1874 = lo1058 ;
  assign po1875 = lo0019 ;
  assign po1876 = lo0020 ;
  assign po1877 = lo0040 ;
  assign po1878 = new_n1974 ;
  assign po1879 = pi000 ;
  assign po1880 = lo1282 ;
  assign po1881 = lo0917 ;
  assign po1882 = lo1060 ;
  assign po1883 = lo1056 ;
  assign po1884 = lo1057 ;
  assign po1885 = lo1059 ;
  assign po1886 = lo1058 ;
  assign po1887 = lo0019 ;
  assign po1888 = lo0020 ;
  assign po1889 = lo0040 ;
  assign po1890 = new_n1977 ;
  assign po1891 = pi000 ;
  assign po1892 = lo1282 ;
  assign po1893 = lo0917 ;
  assign po1894 = lo1060 ;
  assign po1895 = lo1056 ;
  assign po1896 = lo1057 ;
  assign po1897 = lo1059 ;
  assign po1898 = lo1058 ;
  assign po1899 = lo0019 ;
  assign po1900 = lo0020 ;
  assign po1901 = lo0040 ;
  assign po1902 = new_n1980 ;
  assign po1903 = pi000 ;
  assign po1904 = lo1282 ;
  assign po1905 = lo0917 ;
  assign po1906 = lo1060 ;
  assign po1907 = lo1056 ;
  assign po1908 = lo1057 ;
  assign po1909 = lo1059 ;
  assign po1910 = lo1058 ;
  assign po1911 = lo0019 ;
  assign po1912 = lo0020 ;
  assign po1913 = lo0040 ;
  assign po1914 = new_n1983 ;
  assign po1915 = pi000 ;
  assign po1916 = lo1282 ;
  assign po1917 = lo0917 ;
  assign po1918 = lo1060 ;
  assign po1919 = lo1056 ;
  assign po1920 = lo1057 ;
  assign po1921 = lo1059 ;
  assign po1922 = lo1058 ;
  assign po1923 = lo0019 ;
  assign po1924 = lo0020 ;
  assign po1925 = lo0040 ;
  assign po1926 = new_n1986 ;
  assign po1927 = pi000 ;
  assign po1928 = lo1282 ;
  assign po1929 = lo0917 ;
  assign po1930 = lo1060 ;
  assign po1931 = lo1056 ;
  assign po1932 = lo1057 ;
  assign po1933 = lo1059 ;
  assign po1934 = lo1058 ;
  assign po1935 = lo0019 ;
  assign po1936 = lo0020 ;
  assign po1937 = lo0040 ;
  assign po1938 = new_n1994 ;
  assign po1939 = pi000 ;
  assign po1940 = lo1422 ;
  assign po1941 = lo0917 ;
  assign po1942 = lo1060 ;
  assign po1943 = lo1056 ;
  assign po1944 = lo1057 ;
  assign po1945 = lo1059 ;
  assign po1946 = lo1058 ;
  assign po1947 = lo0019 ;
  assign po1948 = lo0020 ;
  assign po1949 = lo0040 ;
  assign po1950 = new_n1995 ;
  assign po1951 = pi000 ;
  assign po1952 = lo1422 ;
  assign po1953 = lo0917 ;
  assign po1954 = lo1060 ;
  assign po1955 = lo1056 ;
  assign po1956 = lo1057 ;
  assign po1957 = lo1059 ;
  assign po1958 = lo1058 ;
  assign po1959 = lo0019 ;
  assign po1960 = lo0020 ;
  assign po1961 = lo0040 ;
  assign po1962 = new_n1996 ;
  assign po1963 = pi000 ;
  assign po1964 = lo1422 ;
  assign po1965 = lo0917 ;
  assign po1966 = lo1060 ;
  assign po1967 = lo1056 ;
  assign po1968 = lo1057 ;
  assign po1969 = lo1059 ;
  assign po1970 = lo1058 ;
  assign po1971 = lo0019 ;
  assign po1972 = lo0020 ;
  assign po1973 = lo0040 ;
  assign po1974 = new_n1997 ;
  assign po1975 = pi000 ;
  assign po1976 = lo1422 ;
  assign po1977 = lo0917 ;
  assign po1978 = lo1060 ;
  assign po1979 = lo1056 ;
  assign po1980 = lo1057 ;
  assign po1981 = lo1059 ;
  assign po1982 = lo1058 ;
  assign po1983 = lo0019 ;
  assign po1984 = lo0020 ;
  assign po1985 = lo0040 ;
  assign po1986 = new_n1998 ;
  assign po1987 = pi000 ;
  assign po1988 = lo1422 ;
  assign po1989 = lo0917 ;
  assign po1990 = lo1060 ;
  assign po1991 = lo1056 ;
  assign po1992 = lo1057 ;
  assign po1993 = lo1059 ;
  assign po1994 = lo1058 ;
  assign po1995 = lo0019 ;
  assign po1996 = lo0020 ;
  assign po1997 = lo0040 ;
  assign po1998 = new_n1999 ;
  assign po1999 = pi000 ;
  assign po2000 = lo1422 ;
  assign po2001 = lo0917 ;
  assign po2002 = lo1060 ;
  assign po2003 = lo1056 ;
  assign po2004 = lo1057 ;
  assign po2005 = lo1059 ;
  assign po2006 = lo1058 ;
  assign po2007 = lo0019 ;
  assign po2008 = lo0020 ;
  assign po2009 = lo0040 ;
  assign po2010 = new_n2000 ;
  assign po2011 = pi000 ;
  assign po2012 = lo1422 ;
  assign po2013 = lo0917 ;
  assign po2014 = lo1060 ;
  assign po2015 = lo1056 ;
  assign po2016 = lo1057 ;
  assign po2017 = lo1059 ;
  assign po2018 = lo1058 ;
  assign po2019 = lo0019 ;
  assign po2020 = lo0020 ;
  assign po2021 = lo0040 ;
  assign po2022 = new_n2001 ;
  assign po2023 = pi000 ;
  assign po2024 = lo1422 ;
  assign po2025 = lo0917 ;
  assign po2026 = lo1060 ;
  assign po2027 = lo1056 ;
  assign po2028 = lo1057 ;
  assign po2029 = lo1059 ;
  assign po2030 = lo1058 ;
  assign po2031 = lo0019 ;
  assign po2032 = lo0020 ;
  assign po2033 = lo0040 ;
  assign po2034 = new_n2003 ;
  assign po2035 = pi000 ;
  assign po2036 = lo1052 ;
  assign po2037 = lo0917 ;
  assign po2038 = lo1060 ;
  assign po2039 = lo1056 ;
  assign po2040 = lo1057 ;
  assign po2041 = lo1059 ;
  assign po2042 = lo1058 ;
  assign po2043 = lo0019 ;
  assign po2044 = lo0020 ;
  assign po2045 = lo0040 ;
  assign po2046 = new_n2004 ;
  assign po2047 = pi000 ;
  assign po2048 = lo1052 ;
  assign po2049 = lo0917 ;
  assign po2050 = lo1060 ;
  assign po2051 = lo1056 ;
  assign po2052 = lo1057 ;
  assign po2053 = lo1059 ;
  assign po2054 = lo1058 ;
  assign po2055 = lo0019 ;
  assign po2056 = lo0020 ;
  assign po2057 = lo0040 ;
  assign po2058 = new_n2005 ;
  assign po2059 = pi000 ;
  assign po2060 = lo1052 ;
  assign po2061 = lo0917 ;
  assign po2062 = lo1060 ;
  assign po2063 = lo1056 ;
  assign po2064 = lo1057 ;
  assign po2065 = lo1059 ;
  assign po2066 = lo1058 ;
  assign po2067 = lo0019 ;
  assign po2068 = lo0020 ;
  assign po2069 = lo0040 ;
  assign po2070 = new_n2006 ;
  assign po2071 = pi000 ;
  assign po2072 = lo1052 ;
  assign po2073 = lo0917 ;
  assign po2074 = lo1060 ;
  assign po2075 = lo1056 ;
  assign po2076 = lo1057 ;
  assign po2077 = lo1059 ;
  assign po2078 = lo1058 ;
  assign po2079 = lo0019 ;
  assign po2080 = lo0020 ;
  assign po2081 = lo0040 ;
  assign po2082 = new_n2007 ;
  assign po2083 = pi000 ;
  assign po2084 = lo1052 ;
  assign po2085 = lo0917 ;
  assign po2086 = lo1060 ;
  assign po2087 = lo1056 ;
  assign po2088 = lo1057 ;
  assign po2089 = lo1059 ;
  assign po2090 = lo1058 ;
  assign po2091 = lo0019 ;
  assign po2092 = lo0020 ;
  assign po2093 = lo0040 ;
  assign po2094 = new_n2008 ;
  assign po2095 = pi000 ;
  assign po2096 = lo1052 ;
  assign po2097 = lo0917 ;
  assign po2098 = lo1060 ;
  assign po2099 = lo1056 ;
  assign po2100 = lo1057 ;
  assign po2101 = lo1059 ;
  assign po2102 = lo1058 ;
  assign po2103 = lo0019 ;
  assign po2104 = lo0020 ;
  assign po2105 = lo0040 ;
  assign po2106 = new_n2009 ;
  assign po2107 = pi000 ;
  assign po2108 = lo1052 ;
  assign po2109 = lo0917 ;
  assign po2110 = lo1060 ;
  assign po2111 = lo1056 ;
  assign po2112 = lo1057 ;
  assign po2113 = lo1059 ;
  assign po2114 = lo1058 ;
  assign po2115 = lo0019 ;
  assign po2116 = lo0020 ;
  assign po2117 = lo0040 ;
  assign po2118 = new_n2010 ;
  assign po2119 = pi000 ;
  assign po2120 = lo1052 ;
  assign po2121 = lo0917 ;
  assign po2122 = lo1060 ;
  assign po2123 = lo1056 ;
  assign po2124 = lo1057 ;
  assign po2125 = lo1059 ;
  assign po2126 = lo1058 ;
  assign po2127 = lo0019 ;
  assign po2128 = lo0020 ;
  assign po2129 = lo0040 ;
  assign po2130 = new_n1994 ;
  assign po2131 = pi000 ;
  assign po2132 = lo1421 ;
  assign po2133 = lo0917 ;
  assign po2134 = lo1060 ;
  assign po2135 = lo1056 ;
  assign po2136 = lo1057 ;
  assign po2137 = lo1059 ;
  assign po2138 = lo1058 ;
  assign po2139 = lo0019 ;
  assign po2140 = lo0020 ;
  assign po2141 = lo0040 ;
  assign po2142 = new_n1995 ;
  assign po2143 = pi000 ;
  assign po2144 = lo1421 ;
  assign po2145 = lo0917 ;
  assign po2146 = lo1060 ;
  assign po2147 = lo1056 ;
  assign po2148 = lo1057 ;
  assign po2149 = lo1059 ;
  assign po2150 = lo1058 ;
  assign po2151 = lo0019 ;
  assign po2152 = lo0020 ;
  assign po2153 = lo0040 ;
  assign po2154 = new_n1996 ;
  assign po2155 = pi000 ;
  assign po2156 = lo1421 ;
  assign po2157 = lo0917 ;
  assign po2158 = lo1060 ;
  assign po2159 = lo1056 ;
  assign po2160 = lo1057 ;
  assign po2161 = lo1059 ;
  assign po2162 = lo1058 ;
  assign po2163 = lo0019 ;
  assign po2164 = lo0020 ;
  assign po2165 = lo0040 ;
  assign po2166 = new_n1997 ;
  assign po2167 = pi000 ;
  assign po2168 = lo1421 ;
  assign po2169 = lo0917 ;
  assign po2170 = lo1060 ;
  assign po2171 = lo1056 ;
  assign po2172 = lo1057 ;
  assign po2173 = lo1059 ;
  assign po2174 = lo1058 ;
  assign po2175 = lo0019 ;
  assign po2176 = lo0020 ;
  assign po2177 = lo0040 ;
  assign po2178 = new_n1998 ;
  assign po2179 = pi000 ;
  assign po2180 = lo1421 ;
  assign po2181 = lo0917 ;
  assign po2182 = lo1060 ;
  assign po2183 = lo1056 ;
  assign po2184 = lo1057 ;
  assign po2185 = lo1059 ;
  assign po2186 = lo1058 ;
  assign po2187 = lo0019 ;
  assign po2188 = lo0020 ;
  assign po2189 = lo0040 ;
  assign po2190 = new_n1999 ;
  assign po2191 = pi000 ;
  assign po2192 = lo1421 ;
  assign po2193 = lo0917 ;
  assign po2194 = lo1060 ;
  assign po2195 = lo1056 ;
  assign po2196 = lo1057 ;
  assign po2197 = lo1059 ;
  assign po2198 = lo1058 ;
  assign po2199 = lo0019 ;
  assign po2200 = lo0020 ;
  assign po2201 = lo0040 ;
  assign po2202 = new_n2000 ;
  assign po2203 = pi000 ;
  assign po2204 = lo1421 ;
  assign po2205 = lo0917 ;
  assign po2206 = lo1060 ;
  assign po2207 = lo1056 ;
  assign po2208 = lo1057 ;
  assign po2209 = lo1059 ;
  assign po2210 = lo1058 ;
  assign po2211 = lo0019 ;
  assign po2212 = lo0020 ;
  assign po2213 = lo0040 ;
  assign po2214 = new_n2001 ;
  assign po2215 = pi000 ;
  assign po2216 = lo1421 ;
  assign po2217 = lo0917 ;
  assign po2218 = lo1060 ;
  assign po2219 = lo1056 ;
  assign po2220 = lo1057 ;
  assign po2221 = lo1059 ;
  assign po2222 = lo1058 ;
  assign po2223 = lo0019 ;
  assign po2224 = lo0020 ;
  assign po2225 = lo0040 ;
  assign po2226 = new_n2003 ;
  assign po2227 = pi000 ;
  assign po2228 = lo1054 ;
  assign po2229 = lo0917 ;
  assign po2230 = lo1060 ;
  assign po2231 = lo1056 ;
  assign po2232 = lo1057 ;
  assign po2233 = lo1059 ;
  assign po2234 = lo1058 ;
  assign po2235 = lo0019 ;
  assign po2236 = lo0020 ;
  assign po2237 = lo0040 ;
  assign po2238 = new_n2004 ;
  assign po2239 = pi000 ;
  assign po2240 = lo1054 ;
  assign po2241 = lo0917 ;
  assign po2242 = lo1060 ;
  assign po2243 = lo1056 ;
  assign po2244 = lo1057 ;
  assign po2245 = lo1059 ;
  assign po2246 = lo1058 ;
  assign po2247 = lo0019 ;
  assign po2248 = lo0020 ;
  assign po2249 = lo0040 ;
  assign po2250 = new_n2005 ;
  assign po2251 = pi000 ;
  assign po2252 = lo1054 ;
  assign po2253 = lo0917 ;
  assign po2254 = lo1060 ;
  assign po2255 = lo1056 ;
  assign po2256 = lo1057 ;
  assign po2257 = lo1059 ;
  assign po2258 = lo1058 ;
  assign po2259 = lo0019 ;
  assign po2260 = lo0020 ;
  assign po2261 = lo0040 ;
  assign po2262 = new_n2006 ;
  assign po2263 = pi000 ;
  assign po2264 = lo1054 ;
  assign po2265 = lo0917 ;
  assign po2266 = lo1060 ;
  assign po2267 = lo1056 ;
  assign po2268 = lo1057 ;
  assign po2269 = lo1059 ;
  assign po2270 = lo1058 ;
  assign po2271 = lo0019 ;
  assign po2272 = lo0020 ;
  assign po2273 = lo0040 ;
  assign po2274 = new_n2007 ;
  assign po2275 = pi000 ;
  assign po2276 = lo1054 ;
  assign po2277 = lo0917 ;
  assign po2278 = lo1060 ;
  assign po2279 = lo1056 ;
  assign po2280 = lo1057 ;
  assign po2281 = lo1059 ;
  assign po2282 = lo1058 ;
  assign po2283 = lo0019 ;
  assign po2284 = lo0020 ;
  assign po2285 = lo0040 ;
  assign po2286 = new_n2008 ;
  assign po2287 = pi000 ;
  assign po2288 = lo1054 ;
  assign po2289 = lo0917 ;
  assign po2290 = lo1060 ;
  assign po2291 = lo1056 ;
  assign po2292 = lo1057 ;
  assign po2293 = lo1059 ;
  assign po2294 = lo1058 ;
  assign po2295 = lo0019 ;
  assign po2296 = lo0020 ;
  assign po2297 = lo0040 ;
  assign po2298 = new_n2009 ;
  assign po2299 = pi000 ;
  assign po2300 = lo1054 ;
  assign po2301 = lo0917 ;
  assign po2302 = lo1060 ;
  assign po2303 = lo1056 ;
  assign po2304 = lo1057 ;
  assign po2305 = lo1059 ;
  assign po2306 = lo1058 ;
  assign po2307 = lo0019 ;
  assign po2308 = lo0020 ;
  assign po2309 = lo0040 ;
  assign po2310 = new_n2010 ;
  assign po2311 = pi000 ;
  assign po2312 = lo1054 ;
  assign po2313 = lo0917 ;
  assign po2314 = lo1060 ;
  assign po2315 = lo1056 ;
  assign po2316 = lo1057 ;
  assign po2317 = lo1059 ;
  assign po2318 = lo1058 ;
  assign po2319 = lo0019 ;
  assign po2320 = lo0020 ;
  assign po2321 = lo0040 ;
  assign po2322 = new_n2012 ;
  assign po2323 = pi000 ;
  assign po2324 = lo1278 ;
  assign po2325 = lo0917 ;
  assign po2326 = lo1060 ;
  assign po2327 = lo1056 ;
  assign po2328 = lo1057 ;
  assign po2329 = lo1059 ;
  assign po2330 = lo1058 ;
  assign po2331 = lo0019 ;
  assign po2332 = lo0020 ;
  assign po2333 = lo0040 ;
  assign po2334 = new_n2013 ;
  assign po2335 = pi000 ;
  assign po2336 = lo1278 ;
  assign po2337 = lo0917 ;
  assign po2338 = lo1060 ;
  assign po2339 = lo1056 ;
  assign po2340 = lo1057 ;
  assign po2341 = lo1059 ;
  assign po2342 = lo1058 ;
  assign po2343 = lo0019 ;
  assign po2344 = lo0020 ;
  assign po2345 = lo0040 ;
  assign po2346 = new_n2014 ;
  assign po2347 = pi000 ;
  assign po2348 = lo1278 ;
  assign po2349 = lo0917 ;
  assign po2350 = lo1060 ;
  assign po2351 = lo1056 ;
  assign po2352 = lo1057 ;
  assign po2353 = lo1059 ;
  assign po2354 = lo1058 ;
  assign po2355 = lo0019 ;
  assign po2356 = lo0020 ;
  assign po2357 = lo0040 ;
  assign po2358 = new_n2015 ;
  assign po2359 = pi000 ;
  assign po2360 = lo1278 ;
  assign po2361 = lo0917 ;
  assign po2362 = lo1060 ;
  assign po2363 = lo1056 ;
  assign po2364 = lo1057 ;
  assign po2365 = lo1059 ;
  assign po2366 = lo1058 ;
  assign po2367 = lo0019 ;
  assign po2368 = lo0020 ;
  assign po2369 = lo0040 ;
  assign po2370 = new_n2016 ;
  assign po2371 = pi000 ;
  assign po2372 = lo1278 ;
  assign po2373 = lo0917 ;
  assign po2374 = lo1060 ;
  assign po2375 = lo1056 ;
  assign po2376 = lo1057 ;
  assign po2377 = lo1059 ;
  assign po2378 = lo1058 ;
  assign po2379 = lo0019 ;
  assign po2380 = lo0020 ;
  assign po2381 = lo0040 ;
  assign po2382 = new_n2017 ;
  assign po2383 = pi000 ;
  assign po2384 = lo1278 ;
  assign po2385 = lo0917 ;
  assign po2386 = lo1060 ;
  assign po2387 = lo1056 ;
  assign po2388 = lo1057 ;
  assign po2389 = lo1059 ;
  assign po2390 = lo1058 ;
  assign po2391 = lo0019 ;
  assign po2392 = lo0020 ;
  assign po2393 = lo0040 ;
  assign po2394 = new_n2018 ;
  assign po2395 = pi000 ;
  assign po2396 = lo1278 ;
  assign po2397 = lo0917 ;
  assign po2398 = lo1060 ;
  assign po2399 = lo1056 ;
  assign po2400 = lo1057 ;
  assign po2401 = lo1059 ;
  assign po2402 = lo1058 ;
  assign po2403 = lo0019 ;
  assign po2404 = lo0020 ;
  assign po2405 = lo0040 ;
  assign po2406 = new_n2019 ;
  assign po2407 = pi000 ;
  assign po2408 = lo1278 ;
  assign po2409 = lo0917 ;
  assign po2410 = lo1060 ;
  assign po2411 = lo1056 ;
  assign po2412 = lo1057 ;
  assign po2413 = lo1059 ;
  assign po2414 = lo1058 ;
  assign po2415 = lo0019 ;
  assign po2416 = lo0020 ;
  assign po2417 = lo0040 ;
  assign po2418 = new_n1974 ;
  assign po2419 = pi000 ;
  assign po2420 = lo1445 ;
  assign po2421 = lo0917 ;
  assign po2422 = lo1060 ;
  assign po2423 = lo1056 ;
  assign po2424 = lo1057 ;
  assign po2425 = lo1059 ;
  assign po2426 = lo1058 ;
  assign po2427 = lo0019 ;
  assign po2428 = lo0020 ;
  assign po2429 = lo0040 ;
  assign po2430 = new_n1977 ;
  assign po2431 = pi000 ;
  assign po2432 = lo1445 ;
  assign po2433 = lo0917 ;
  assign po2434 = lo1060 ;
  assign po2435 = lo1056 ;
  assign po2436 = lo1057 ;
  assign po2437 = lo1059 ;
  assign po2438 = lo1058 ;
  assign po2439 = lo0019 ;
  assign po2440 = lo0020 ;
  assign po2441 = lo0040 ;
  assign po2442 = new_n1980 ;
  assign po2443 = pi000 ;
  assign po2444 = lo1445 ;
  assign po2445 = lo0917 ;
  assign po2446 = lo1060 ;
  assign po2447 = lo1056 ;
  assign po2448 = lo1057 ;
  assign po2449 = lo1059 ;
  assign po2450 = lo1058 ;
  assign po2451 = lo0019 ;
  assign po2452 = lo0020 ;
  assign po2453 = lo0040 ;
  assign po2454 = new_n1983 ;
  assign po2455 = pi000 ;
  assign po2456 = lo1445 ;
  assign po2457 = lo0917 ;
  assign po2458 = lo1060 ;
  assign po2459 = lo1056 ;
  assign po2460 = lo1057 ;
  assign po2461 = lo1059 ;
  assign po2462 = lo1058 ;
  assign po2463 = lo0019 ;
  assign po2464 = lo0020 ;
  assign po2465 = lo0040 ;
  assign po2466 = new_n1986 ;
  assign po2467 = pi000 ;
  assign po2468 = lo1445 ;
  assign po2469 = lo0917 ;
  assign po2470 = lo1060 ;
  assign po2471 = lo1056 ;
  assign po2472 = lo1057 ;
  assign po2473 = lo1059 ;
  assign po2474 = lo1058 ;
  assign po2475 = lo0019 ;
  assign po2476 = lo0020 ;
  assign po2477 = lo0040 ;
  assign po2478 = new_n1988 ;
  assign po2479 = pi000 ;
  assign po2480 = lo1445 ;
  assign po2481 = lo0917 ;
  assign po2482 = lo1060 ;
  assign po2483 = lo1056 ;
  assign po2484 = lo1057 ;
  assign po2485 = lo1059 ;
  assign po2486 = lo1058 ;
  assign po2487 = lo0019 ;
  assign po2488 = lo0020 ;
  assign po2489 = lo0040 ;
  assign po2490 = new_n1990 ;
  assign po2491 = pi000 ;
  assign po2492 = lo1445 ;
  assign po2493 = lo0917 ;
  assign po2494 = lo1060 ;
  assign po2495 = lo1056 ;
  assign po2496 = lo1057 ;
  assign po2497 = lo1059 ;
  assign po2498 = lo1058 ;
  assign po2499 = lo0019 ;
  assign po2500 = lo0020 ;
  assign po2501 = lo0040 ;
  assign po2502 = new_n1992 ;
  assign po2503 = pi000 ;
  assign po2504 = lo1445 ;
  assign po2505 = lo0917 ;
  assign po2506 = lo1060 ;
  assign po2507 = lo1056 ;
  assign po2508 = lo1057 ;
  assign po2509 = lo1059 ;
  assign po2510 = lo1058 ;
  assign po2511 = lo0019 ;
  assign po2512 = lo0020 ;
  assign po2513 = lo0040 ;
  assign po2514 = new_n2012 ;
  assign po2515 = pi000 ;
  assign po2516 = lo1273 ;
  assign po2517 = lo0917 ;
  assign po2518 = lo1060 ;
  assign po2519 = lo1056 ;
  assign po2520 = lo1057 ;
  assign po2521 = lo1059 ;
  assign po2522 = lo1058 ;
  assign po2523 = lo0019 ;
  assign po2524 = lo0020 ;
  assign po2525 = lo0040 ;
  assign po2526 = new_n2013 ;
  assign po2527 = pi000 ;
  assign po2528 = lo1273 ;
  assign po2529 = lo0917 ;
  assign po2530 = lo1060 ;
  assign po2531 = lo1056 ;
  assign po2532 = lo1057 ;
  assign po2533 = lo1059 ;
  assign po2534 = lo1058 ;
  assign po2535 = lo0019 ;
  assign po2536 = lo0020 ;
  assign po2537 = lo0040 ;
  assign po2538 = new_n2014 ;
  assign po2539 = pi000 ;
  assign po2540 = lo1273 ;
  assign po2541 = lo0917 ;
  assign po2542 = lo1060 ;
  assign po2543 = lo1056 ;
  assign po2544 = lo1057 ;
  assign po2545 = lo1059 ;
  assign po2546 = lo1058 ;
  assign po2547 = lo0019 ;
  assign po2548 = lo0020 ;
  assign po2549 = lo0040 ;
  assign po2550 = new_n2015 ;
  assign po2551 = pi000 ;
  assign po2552 = lo1273 ;
  assign po2553 = lo0917 ;
  assign po2554 = lo1060 ;
  assign po2555 = lo1056 ;
  assign po2556 = lo1057 ;
  assign po2557 = lo1059 ;
  assign po2558 = lo1058 ;
  assign po2559 = lo0019 ;
  assign po2560 = lo0020 ;
  assign po2561 = lo0040 ;
  assign po2562 = new_n2016 ;
  assign po2563 = pi000 ;
  assign po2564 = lo1273 ;
  assign po2565 = lo0917 ;
  assign po2566 = lo1060 ;
  assign po2567 = lo1056 ;
  assign po2568 = lo1057 ;
  assign po2569 = lo1059 ;
  assign po2570 = lo1058 ;
  assign po2571 = lo0019 ;
  assign po2572 = lo0020 ;
  assign po2573 = lo0040 ;
  assign po2574 = new_n2017 ;
  assign po2575 = pi000 ;
  assign po2576 = lo1273 ;
  assign po2577 = lo0917 ;
  assign po2578 = lo1060 ;
  assign po2579 = lo1056 ;
  assign po2580 = lo1057 ;
  assign po2581 = lo1059 ;
  assign po2582 = lo1058 ;
  assign po2583 = lo0019 ;
  assign po2584 = lo0020 ;
  assign po2585 = lo0040 ;
  assign po2586 = new_n2018 ;
  assign po2587 = pi000 ;
  assign po2588 = lo1273 ;
  assign po2589 = lo0917 ;
  assign po2590 = lo1060 ;
  assign po2591 = lo1056 ;
  assign po2592 = lo1057 ;
  assign po2593 = lo1059 ;
  assign po2594 = lo1058 ;
  assign po2595 = lo0019 ;
  assign po2596 = lo0020 ;
  assign po2597 = lo0040 ;
  assign po2598 = new_n2019 ;
  assign po2599 = pi000 ;
  assign po2600 = lo1273 ;
  assign po2601 = lo0917 ;
  assign po2602 = lo1060 ;
  assign po2603 = lo1056 ;
  assign po2604 = lo1057 ;
  assign po2605 = lo1059 ;
  assign po2606 = lo1058 ;
  assign po2607 = lo0019 ;
  assign po2608 = lo0020 ;
  assign po2609 = lo0040 ;
  assign po2610 = new_n1988 ;
  assign po2611 = pi000 ;
  assign po2612 = lo1281 ;
  assign po2613 = lo0917 ;
  assign po2614 = lo1060 ;
  assign po2615 = lo1056 ;
  assign po2616 = lo1057 ;
  assign po2617 = lo1059 ;
  assign po2618 = lo1058 ;
  assign po2619 = lo0019 ;
  assign po2620 = lo0020 ;
  assign po2621 = lo0040 ;
  assign po2622 = new_n1992 ;
  assign po2623 = pi000 ;
  assign po2624 = lo1281 ;
  assign po2625 = lo0917 ;
  assign po2626 = lo1060 ;
  assign po2627 = lo1056 ;
  assign po2628 = lo1057 ;
  assign po2629 = lo1059 ;
  assign po2630 = lo1058 ;
  assign po2631 = lo0019 ;
  assign po2632 = lo0020 ;
  assign po2633 = lo0040 ;
  assign po2634 = new_n1990 ;
  assign po2635 = pi000 ;
  assign po2636 = lo1281 ;
  assign po2637 = lo0917 ;
  assign po2638 = lo1060 ;
  assign po2639 = lo1056 ;
  assign po2640 = lo1057 ;
  assign po2641 = lo1059 ;
  assign po2642 = lo1058 ;
  assign po2643 = lo0019 ;
  assign po2644 = lo0020 ;
  assign po2645 = lo0040 ;
  assign po2646 = new_n1974 ;
  assign po2647 = pi000 ;
  assign po2648 = lo1281 ;
  assign po2649 = lo0917 ;
  assign po2650 = lo1060 ;
  assign po2651 = lo1056 ;
  assign po2652 = lo1057 ;
  assign po2653 = lo1059 ;
  assign po2654 = lo1058 ;
  assign po2655 = lo0019 ;
  assign po2656 = lo0020 ;
  assign po2657 = lo0040 ;
  assign po2658 = new_n1977 ;
  assign po2659 = pi000 ;
  assign po2660 = lo1281 ;
  assign po2661 = lo0917 ;
  assign po2662 = lo1060 ;
  assign po2663 = lo1056 ;
  assign po2664 = lo1057 ;
  assign po2665 = lo1059 ;
  assign po2666 = lo1058 ;
  assign po2667 = lo0019 ;
  assign po2668 = lo0020 ;
  assign po2669 = lo0040 ;
  assign po2670 = new_n1980 ;
  assign po2671 = pi000 ;
  assign po2672 = lo1281 ;
  assign po2673 = lo0917 ;
  assign po2674 = lo1060 ;
  assign po2675 = lo1056 ;
  assign po2676 = lo1057 ;
  assign po2677 = lo1059 ;
  assign po2678 = lo1058 ;
  assign po2679 = lo0019 ;
  assign po2680 = lo0020 ;
  assign po2681 = lo0040 ;
  assign po2682 = new_n1983 ;
  assign po2683 = pi000 ;
  assign po2684 = lo1281 ;
  assign po2685 = lo0917 ;
  assign po2686 = lo1060 ;
  assign po2687 = lo1056 ;
  assign po2688 = lo1057 ;
  assign po2689 = lo1059 ;
  assign po2690 = lo1058 ;
  assign po2691 = lo0019 ;
  assign po2692 = lo0020 ;
  assign po2693 = lo0040 ;
  assign po2694 = new_n1986 ;
  assign po2695 = pi000 ;
  assign po2696 = lo1281 ;
  assign po2697 = lo0917 ;
  assign po2698 = lo1060 ;
  assign po2699 = lo1056 ;
  assign po2700 = lo1057 ;
  assign po2701 = lo1059 ;
  assign po2702 = lo1058 ;
  assign po2703 = lo0019 ;
  assign po2704 = lo0020 ;
  assign po2705 = lo0040 ;
  assign po2706 = new_n2012 ;
  assign po2707 = pi000 ;
  assign po2708 = lo1276 ;
  assign po2709 = lo0917 ;
  assign po2710 = lo1060 ;
  assign po2711 = lo1056 ;
  assign po2712 = lo1057 ;
  assign po2713 = lo1059 ;
  assign po2714 = lo1058 ;
  assign po2715 = lo0019 ;
  assign po2716 = lo0020 ;
  assign po2717 = lo0040 ;
  assign po2718 = new_n2013 ;
  assign po2719 = pi000 ;
  assign po2720 = lo1276 ;
  assign po2721 = lo0917 ;
  assign po2722 = lo1060 ;
  assign po2723 = lo1056 ;
  assign po2724 = lo1057 ;
  assign po2725 = lo1059 ;
  assign po2726 = lo1058 ;
  assign po2727 = lo0019 ;
  assign po2728 = lo0020 ;
  assign po2729 = lo0040 ;
  assign po2730 = new_n2014 ;
  assign po2731 = pi000 ;
  assign po2732 = lo1276 ;
  assign po2733 = lo0917 ;
  assign po2734 = lo1060 ;
  assign po2735 = lo1056 ;
  assign po2736 = lo1057 ;
  assign po2737 = lo1059 ;
  assign po2738 = lo1058 ;
  assign po2739 = lo0019 ;
  assign po2740 = lo0020 ;
  assign po2741 = lo0040 ;
  assign po2742 = new_n2015 ;
  assign po2743 = pi000 ;
  assign po2744 = lo1276 ;
  assign po2745 = lo0917 ;
  assign po2746 = lo1060 ;
  assign po2747 = lo1056 ;
  assign po2748 = lo1057 ;
  assign po2749 = lo1059 ;
  assign po2750 = lo1058 ;
  assign po2751 = lo0019 ;
  assign po2752 = lo0020 ;
  assign po2753 = lo0040 ;
  assign po2754 = new_n2016 ;
  assign po2755 = pi000 ;
  assign po2756 = lo1276 ;
  assign po2757 = lo0917 ;
  assign po2758 = lo1060 ;
  assign po2759 = lo1056 ;
  assign po2760 = lo1057 ;
  assign po2761 = lo1059 ;
  assign po2762 = lo1058 ;
  assign po2763 = lo0019 ;
  assign po2764 = lo0020 ;
  assign po2765 = lo0040 ;
  assign po2766 = new_n2017 ;
  assign po2767 = pi000 ;
  assign po2768 = lo1276 ;
  assign po2769 = lo0917 ;
  assign po2770 = lo1060 ;
  assign po2771 = lo1056 ;
  assign po2772 = lo1057 ;
  assign po2773 = lo1059 ;
  assign po2774 = lo1058 ;
  assign po2775 = lo0019 ;
  assign po2776 = lo0020 ;
  assign po2777 = lo0040 ;
  assign po2778 = new_n2018 ;
  assign po2779 = pi000 ;
  assign po2780 = lo1276 ;
  assign po2781 = lo0917 ;
  assign po2782 = lo1060 ;
  assign po2783 = lo1056 ;
  assign po2784 = lo1057 ;
  assign po2785 = lo1059 ;
  assign po2786 = lo1058 ;
  assign po2787 = lo0019 ;
  assign po2788 = lo0020 ;
  assign po2789 = lo0040 ;
  assign po2790 = new_n2019 ;
  assign po2791 = pi000 ;
  assign po2792 = lo1276 ;
  assign po2793 = lo0917 ;
  assign po2794 = lo1060 ;
  assign po2795 = lo1056 ;
  assign po2796 = lo1057 ;
  assign po2797 = lo1059 ;
  assign po2798 = lo1058 ;
  assign po2799 = lo0019 ;
  assign po2800 = lo0020 ;
  assign po2801 = lo0040 ;
  assign po2802 = new_n1988 ;
  assign po2803 = pi000 ;
  assign po2804 = lo1284 ;
  assign po2805 = lo0917 ;
  assign po2806 = lo1060 ;
  assign po2807 = lo1056 ;
  assign po2808 = lo1057 ;
  assign po2809 = lo1059 ;
  assign po2810 = lo1058 ;
  assign po2811 = lo0019 ;
  assign po2812 = lo0020 ;
  assign po2813 = lo0040 ;
  assign po2814 = new_n1992 ;
  assign po2815 = pi000 ;
  assign po2816 = lo1284 ;
  assign po2817 = lo0917 ;
  assign po2818 = lo1060 ;
  assign po2819 = lo1056 ;
  assign po2820 = lo1057 ;
  assign po2821 = lo1059 ;
  assign po2822 = lo1058 ;
  assign po2823 = lo0019 ;
  assign po2824 = lo0020 ;
  assign po2825 = lo0040 ;
  assign po2826 = new_n1990 ;
  assign po2827 = pi000 ;
  assign po2828 = lo1284 ;
  assign po2829 = lo0917 ;
  assign po2830 = lo1060 ;
  assign po2831 = lo1056 ;
  assign po2832 = lo1057 ;
  assign po2833 = lo1059 ;
  assign po2834 = lo1058 ;
  assign po2835 = lo0019 ;
  assign po2836 = lo0020 ;
  assign po2837 = lo0040 ;
  assign po2838 = new_n1974 ;
  assign po2839 = pi000 ;
  assign po2840 = lo1284 ;
  assign po2841 = lo0917 ;
  assign po2842 = lo1060 ;
  assign po2843 = lo1056 ;
  assign po2844 = lo1057 ;
  assign po2845 = lo1059 ;
  assign po2846 = lo1058 ;
  assign po2847 = lo0019 ;
  assign po2848 = lo0020 ;
  assign po2849 = lo0040 ;
  assign po2850 = new_n1977 ;
  assign po2851 = pi000 ;
  assign po2852 = lo1284 ;
  assign po2853 = lo0917 ;
  assign po2854 = lo1060 ;
  assign po2855 = lo1056 ;
  assign po2856 = lo1057 ;
  assign po2857 = lo1059 ;
  assign po2858 = lo1058 ;
  assign po2859 = lo0019 ;
  assign po2860 = lo0020 ;
  assign po2861 = lo0040 ;
  assign po2862 = new_n1980 ;
  assign po2863 = pi000 ;
  assign po2864 = lo1284 ;
  assign po2865 = lo0917 ;
  assign po2866 = lo1060 ;
  assign po2867 = lo1056 ;
  assign po2868 = lo1057 ;
  assign po2869 = lo1059 ;
  assign po2870 = lo1058 ;
  assign po2871 = lo0019 ;
  assign po2872 = lo0020 ;
  assign po2873 = lo0040 ;
  assign po2874 = new_n1983 ;
  assign po2875 = pi000 ;
  assign po2876 = lo1284 ;
  assign po2877 = lo0917 ;
  assign po2878 = lo1060 ;
  assign po2879 = lo1056 ;
  assign po2880 = lo1057 ;
  assign po2881 = lo1059 ;
  assign po2882 = lo1058 ;
  assign po2883 = lo0019 ;
  assign po2884 = lo0020 ;
  assign po2885 = lo0040 ;
  assign po2886 = new_n1986 ;
  assign po2887 = pi000 ;
  assign po2888 = lo1284 ;
  assign po2889 = lo0917 ;
  assign po2890 = lo1060 ;
  assign po2891 = lo1056 ;
  assign po2892 = lo1057 ;
  assign po2893 = lo1059 ;
  assign po2894 = lo1058 ;
  assign po2895 = lo0019 ;
  assign po2896 = lo0020 ;
  assign po2897 = lo0040 ;
  assign po2898 = new_n2012 ;
  assign po2899 = pi000 ;
  assign po2900 = lo1272 ;
  assign po2901 = lo0917 ;
  assign po2902 = lo1060 ;
  assign po2903 = lo1056 ;
  assign po2904 = lo1057 ;
  assign po2905 = lo1059 ;
  assign po2906 = lo1058 ;
  assign po2907 = lo0019 ;
  assign po2908 = lo0020 ;
  assign po2909 = lo0040 ;
  assign po2910 = new_n2013 ;
  assign po2911 = pi000 ;
  assign po2912 = lo1272 ;
  assign po2913 = lo0917 ;
  assign po2914 = lo1060 ;
  assign po2915 = lo1056 ;
  assign po2916 = lo1057 ;
  assign po2917 = lo1059 ;
  assign po2918 = lo1058 ;
  assign po2919 = lo0019 ;
  assign po2920 = lo0020 ;
  assign po2921 = lo0040 ;
  assign po2922 = new_n2014 ;
  assign po2923 = pi000 ;
  assign po2924 = lo1272 ;
  assign po2925 = lo0917 ;
  assign po2926 = lo1060 ;
  assign po2927 = lo1056 ;
  assign po2928 = lo1057 ;
  assign po2929 = lo1059 ;
  assign po2930 = lo1058 ;
  assign po2931 = lo0019 ;
  assign po2932 = lo0020 ;
  assign po2933 = lo0040 ;
  assign po2934 = new_n2015 ;
  assign po2935 = pi000 ;
  assign po2936 = lo1272 ;
  assign po2937 = lo0917 ;
  assign po2938 = lo1060 ;
  assign po2939 = lo1056 ;
  assign po2940 = lo1057 ;
  assign po2941 = lo1059 ;
  assign po2942 = lo1058 ;
  assign po2943 = lo0019 ;
  assign po2944 = lo0020 ;
  assign po2945 = lo0040 ;
  assign po2946 = new_n2016 ;
  assign po2947 = pi000 ;
  assign po2948 = lo1272 ;
  assign po2949 = lo0917 ;
  assign po2950 = lo1060 ;
  assign po2951 = lo1056 ;
  assign po2952 = lo1057 ;
  assign po2953 = lo1059 ;
  assign po2954 = lo1058 ;
  assign po2955 = lo0019 ;
  assign po2956 = lo0020 ;
  assign po2957 = lo0040 ;
  assign po2958 = new_n2017 ;
  assign po2959 = pi000 ;
  assign po2960 = lo1272 ;
  assign po2961 = lo0917 ;
  assign po2962 = lo1060 ;
  assign po2963 = lo1056 ;
  assign po2964 = lo1057 ;
  assign po2965 = lo1059 ;
  assign po2966 = lo1058 ;
  assign po2967 = lo0019 ;
  assign po2968 = lo0020 ;
  assign po2969 = lo0040 ;
  assign po2970 = new_n2018 ;
  assign po2971 = pi000 ;
  assign po2972 = lo1272 ;
  assign po2973 = lo0917 ;
  assign po2974 = lo1060 ;
  assign po2975 = lo1056 ;
  assign po2976 = lo1057 ;
  assign po2977 = lo1059 ;
  assign po2978 = lo1058 ;
  assign po2979 = lo0019 ;
  assign po2980 = lo0020 ;
  assign po2981 = lo0040 ;
  assign po2982 = new_n2019 ;
  assign po2983 = pi000 ;
  assign po2984 = lo1272 ;
  assign po2985 = lo0917 ;
  assign po2986 = lo1060 ;
  assign po2987 = lo1056 ;
  assign po2988 = lo1057 ;
  assign po2989 = lo1059 ;
  assign po2990 = lo1058 ;
  assign po2991 = lo0019 ;
  assign po2992 = lo0020 ;
  assign po2993 = lo0040 ;
  assign po2994 = new_n1988 ;
  assign po2995 = pi000 ;
  assign po2996 = lo1280 ;
  assign po2997 = lo0917 ;
  assign po2998 = lo1060 ;
  assign po2999 = lo1056 ;
  assign po3000 = lo1057 ;
  assign po3001 = lo1059 ;
  assign po3002 = lo1058 ;
  assign po3003 = lo0019 ;
  assign po3004 = lo0020 ;
  assign po3005 = lo0040 ;
  assign po3006 = new_n1992 ;
  assign po3007 = pi000 ;
  assign po3008 = lo1280 ;
  assign po3009 = lo0917 ;
  assign po3010 = lo1060 ;
  assign po3011 = lo1056 ;
  assign po3012 = lo1057 ;
  assign po3013 = lo1059 ;
  assign po3014 = lo1058 ;
  assign po3015 = lo0019 ;
  assign po3016 = lo0020 ;
  assign po3017 = lo0040 ;
  assign po3018 = new_n1990 ;
  assign po3019 = pi000 ;
  assign po3020 = lo1280 ;
  assign po3021 = lo0917 ;
  assign po3022 = lo1060 ;
  assign po3023 = lo1056 ;
  assign po3024 = lo1057 ;
  assign po3025 = lo1059 ;
  assign po3026 = lo1058 ;
  assign po3027 = lo0019 ;
  assign po3028 = lo0020 ;
  assign po3029 = lo0040 ;
  assign po3030 = new_n1974 ;
  assign po3031 = pi000 ;
  assign po3032 = lo1280 ;
  assign po3033 = lo0917 ;
  assign po3034 = lo1060 ;
  assign po3035 = lo1056 ;
  assign po3036 = lo1057 ;
  assign po3037 = lo1059 ;
  assign po3038 = lo1058 ;
  assign po3039 = lo0019 ;
  assign po3040 = lo0020 ;
  assign po3041 = lo0040 ;
  assign po3042 = new_n1977 ;
  assign po3043 = pi000 ;
  assign po3044 = lo1280 ;
  assign po3045 = lo0917 ;
  assign po3046 = lo1060 ;
  assign po3047 = lo1056 ;
  assign po3048 = lo1057 ;
  assign po3049 = lo1059 ;
  assign po3050 = lo1058 ;
  assign po3051 = lo0019 ;
  assign po3052 = lo0020 ;
  assign po3053 = lo0040 ;
  assign po3054 = new_n1980 ;
  assign po3055 = pi000 ;
  assign po3056 = lo1280 ;
  assign po3057 = lo0917 ;
  assign po3058 = lo1060 ;
  assign po3059 = lo1056 ;
  assign po3060 = lo1057 ;
  assign po3061 = lo1059 ;
  assign po3062 = lo1058 ;
  assign po3063 = lo0019 ;
  assign po3064 = lo0020 ;
  assign po3065 = lo0040 ;
  assign po3066 = new_n1983 ;
  assign po3067 = pi000 ;
  assign po3068 = lo1280 ;
  assign po3069 = lo0917 ;
  assign po3070 = lo1060 ;
  assign po3071 = lo1056 ;
  assign po3072 = lo1057 ;
  assign po3073 = lo1059 ;
  assign po3074 = lo1058 ;
  assign po3075 = lo0019 ;
  assign po3076 = lo0020 ;
  assign po3077 = lo0040 ;
  assign po3078 = new_n1986 ;
  assign po3079 = pi000 ;
  assign po3080 = lo1280 ;
  assign po3081 = lo0917 ;
  assign po3082 = lo1060 ;
  assign po3083 = lo1056 ;
  assign po3084 = lo1057 ;
  assign po3085 = lo1059 ;
  assign po3086 = lo1058 ;
  assign po3087 = lo0019 ;
  assign po3088 = lo0020 ;
  assign po3089 = lo0040 ;
  assign po3090 = ~new_n2025 ;
  assign po3091 = ~new_n2028 ;
  assign po3092 = ~new_n2031 ;
  assign po3093 = ~new_n2034 ;
  assign po3094 = ~new_n2037 ;
  assign po3095 = ~new_n2040 ;
  assign po3096 = ~new_n2043 ;
  assign po3097 = ~new_n2046 ;
  assign po3098 = ~new_n2049 ;
  assign po3099 = ~new_n2052 ;
  assign po3100 = ~new_n2055 ;
  assign po3101 = ~new_n2058 ;
  assign po3102 = ~new_n2061 ;
  assign po3103 = ~new_n2064 ;
  assign po3104 = ~new_n2067 ;
  assign po3105 = new_n2075 ;
  assign po3106 = new_n2079 ;
  assign po3107 = new_n2083 ;
  assign po3108 = new_n2087 ;
  assign po3109 = new_n2091 ;
  assign po3110 = new_n2095 ;
  assign po3111 = new_n2099 ;
  assign po3112 = new_n2103 ;
  assign po3113 = new_n2107 ;
  assign po3114 = new_n2111 ;
  assign po3115 = new_n2115 ;
  assign po3116 = new_n2119 ;
  assign po3117 = new_n2123 ;
  assign po3118 = new_n2127 ;
  assign po3119 = new_n2131 ;
  assign po3120 = new_n2135 ;
  assign po3121 = ~new_n2142 ;
  assign po3122 = ~new_n2145 ;
  assign po3123 = ~new_n2148 ;
  assign po3124 = ~new_n2151 ;
  assign po3125 = ~new_n2154 ;
  assign po3126 = ~new_n2157 ;
  assign po3127 = ~new_n2160 ;
  assign po3128 = ~new_n2163 ;
  assign po3129 = ~new_n2166 ;
  assign po3130 = ~new_n2169 ;
  assign po3131 = ~new_n2172 ;
  assign po3132 = ~new_n2175 ;
  assign po3133 = ~new_n2178 ;
  assign po3134 = ~new_n2181 ;
  assign po3135 = ~new_n2184 ;
  assign po3136 = new_n2186 ;
  assign po3137 = ~new_n2064 ;
  assign po3138 = ~new_n2067 ;
  assign po3139 = new_n2075 ;
  assign po3140 = new_n2079 ;
  assign po3141 = new_n2083 ;
  assign po3142 = new_n2087 ;
  assign po3143 = new_n2091 ;
  assign po3144 = new_n2095 ;
  assign po3145 = new_n2099 ;
  assign po3146 = new_n2103 ;
  assign po3147 = new_n2107 ;
  assign po3148 = new_n2111 ;
  assign po3149 = new_n2115 ;
  assign po3150 = new_n2119 ;
  assign po3151 = new_n2123 ;
  assign po3152 = new_n2127 ;
  assign po3153 = new_n2131 ;
  assign po3154 = new_n2135 ;
  assign po3155 = ~new_n2025 ;
  assign po3156 = ~new_n2028 ;
  assign po3157 = ~new_n2031 ;
  assign po3158 = ~new_n2034 ;
  assign po3159 = ~new_n2037 ;
  assign po3160 = ~new_n2040 ;
  assign po3161 = ~new_n2043 ;
  assign po3162 = ~new_n2046 ;
  assign po3163 = ~new_n2049 ;
  assign po3164 = ~new_n2052 ;
  assign po3165 = ~new_n2055 ;
  assign po3166 = ~new_n2058 ;
  assign po3167 = ~new_n2061 ;
  assign po3168 = ~new_n2142 ;
  assign po3169 = ~new_n2145 ;
  assign po3170 = ~new_n2148 ;
  assign po3171 = ~new_n2151 ;
  assign po3172 = ~new_n2154 ;
  assign po3173 = ~new_n2157 ;
  assign po3174 = ~new_n2160 ;
  assign po3175 = ~new_n2163 ;
  assign po3176 = ~new_n2166 ;
  assign po3177 = ~new_n2169 ;
  assign po3178 = ~new_n2172 ;
  assign po3179 = ~new_n2175 ;
  assign po3180 = ~new_n2178 ;
  assign po3181 = ~new_n2181 ;
  assign po3182 = ~new_n2184 ;
  assign po3183 = new_n2186 ;
  assign po3184 = pi273 ;
  assign po3185 = pi274 ;
  assign po3186 = pi275 ;
  assign po3187 = pi276 ;
  assign po3188 = pi277 ;
  assign po3189 = pi278 ;
  assign po3190 = pi279 ;
  assign po3191 = pi280 ;
  assign po3192 = pi281 ;
  assign po3193 = pi282 ;
  assign po3194 = pi283 ;
  assign po3195 = pi284 ;
  assign po3196 = pi285 ;
  assign po3197 = pi286 ;
  assign po3198 = pi287 ;
  assign po3199 = pi288 ;
  assign po3200 = pi289 ;
  assign po3201 = pi290 ;
  assign po3202 = pi291 ;
  assign po3203 = pi292 ;
  assign po3204 = pi293 ;
  assign po3205 = pi294 ;
  assign po3206 = pi295 ;
  assign po3207 = pi296 ;
  assign po3208 = pi297 ;
  assign po3209 = pi298 ;
  assign po3210 = pi299 ;
  assign po3211 = pi300 ;
  assign po3212 = pi301 ;
  assign po3213 = pi302 ;
  assign po3214 = pi303 ;
  assign po3215 = pi304 ;
  assign po3216 = pi305 ;
  assign po3217 = pi306 ;
  assign po3218 = pi307 ;
  assign po3219 = pi308 ;
  assign po3220 = pi309 ;
  assign po3221 = pi310 ;
  assign po3222 = pi311 ;
  assign po3223 = pi312 ;
  assign po3224 = pi313 ;
  assign po3225 = pi314 ;
  assign po3226 = pi315 ;
  assign po3227 = pi316 ;
  assign po3228 = pi317 ;
  assign po3229 = pi318 ;
  assign po3230 = pi319 ;
  assign po3231 = pi320 ;
  assign po3232 = pi321 ;
  assign po3233 = pi322 ;
  assign po3234 = pi323 ;
  assign po3235 = pi324 ;
  assign po3236 = pi325 ;
  assign po3237 = pi326 ;
  assign po3238 = pi327 ;
  assign po3239 = pi328 ;
  assign po3240 = pi329 ;
  assign po3241 = pi330 ;
  assign po3242 = pi331 ;
  assign po3243 = pi332 ;
  assign po3244 = pi333 ;
  assign po3245 = pi334 ;
  assign po3246 = pi335 ;
  assign po3247 = pi336 ;
  assign po3248 = pi337 ;
  assign po3249 = pi338 ;
  assign po3250 = pi339 ;
  assign po3251 = pi340 ;
  assign po3252 = pi341 ;
  assign po3253 = pi342 ;
  assign po3254 = pi343 ;
  assign po3255 = pi344 ;
  assign po3256 = pi345 ;
  assign po3257 = pi346 ;
  assign po3258 = pi347 ;
  assign po3259 = pi348 ;
  assign po3260 = pi349 ;
  assign po3261 = pi350 ;
  assign po3262 = pi351 ;
  assign po3263 = pi352 ;
  assign po3264 = pi353 ;
  assign po3265 = pi354 ;
  assign po3266 = pi355 ;
  assign po3267 = pi356 ;
  assign po3268 = pi357 ;
  assign po3269 = pi358 ;
  assign po3270 = pi359 ;
  assign po3271 = pi360 ;
  assign po3272 = pi361 ;
  assign po3273 = pi362 ;
  assign po3274 = pi363 ;
  assign po3275 = pi364 ;
  assign po3276 = pi365 ;
  assign po3277 = pi366 ;
  assign po3278 = pi367 ;
  assign po3279 = pi368 ;
  assign po3280 = pi369 ;
  assign po3281 = pi370 ;
  assign po3282 = pi371 ;
  assign po3283 = pi372 ;
  assign po3284 = pi373 ;
  assign po3285 = pi374 ;
  assign po3286 = pi375 ;
  assign po3287 = pi376 ;
  assign po3288 = pi377 ;
  assign po3289 = pi378 ;
  assign po3290 = pi379 ;
  assign po3291 = pi380 ;
  assign po3292 = pi381 ;
  assign po3293 = pi382 ;
  assign po3294 = pi383 ;
  assign po3295 = pi384 ;
  assign po3296 = pi385 ;
  assign po3297 = pi386 ;
  assign po3298 = pi387 ;
  assign po3299 = pi388 ;
  assign po3300 = pi389 ;
  assign po3301 = pi390 ;
  assign po3302 = pi391 ;
  assign po3303 = pi392 ;
  assign po3304 = pi393 ;
  assign po3305 = pi394 ;
  assign po3306 = pi395 ;
  assign po3307 = pi396 ;
  assign po3308 = pi397 ;
  assign po3309 = pi398 ;
  assign po3310 = pi399 ;
  assign po3311 = pi400 ;
  assign po3312 = pi401 ;
  assign po3313 = pi402 ;
  assign po3314 = pi403 ;
  assign po3315 = pi404 ;
  assign po3316 = pi405 ;
  assign po3317 = pi406 ;
  assign po3318 = pi407 ;
  assign po3319 = pi408 ;
  assign po3320 = pi409 ;
  assign po3321 = pi410 ;
  assign po3322 = pi411 ;
  assign po3323 = pi412 ;
  assign po3324 = pi413 ;
  assign po3325 = pi414 ;
  assign po3326 = pi415 ;
  assign po3327 = pi416 ;
  assign li0000 = ~new_n2191 ;
  assign li0001 = ~new_n2194 ;
  assign li0002 = ~new_n2197 ;
  assign li0003 = ~new_n2201 ;
  assign li0004 = ~new_n2204 ;
  assign li0005 = ~new_n2207 ;
  assign li0006 = ~new_n2210 ;
  assign li0007 = ~new_n2213 ;
  assign li0008 = ~new_n2216 ;
  assign li0009 = ~new_n2219 ;
  assign li0010 = ~new_n2222 ;
  assign li0011 = ~new_n2226 ;
  assign li0012 = ~new_n2229 ;
  assign li0013 = ~new_n2232 ;
  assign li0014 = ~new_n2235 ;
  assign li0015 = ~new_n2238 ;
  assign li0016 = new_n2246 ;
  assign li0017 = lo0894 ;
  assign li0018 = ~new_n13929 ;
  assign li0019 = ~new_n13970 ;
  assign li0020 = ~new_n13998 ;
  assign li0021 = ~new_n14029 ;
  assign li0022 = ~new_n14053 ;
  assign li0023 = ~new_n14094 ;
  assign li0024 = ~new_n14121 ;
  assign li0025 = ~new_n14147 ;
  assign li0026 = ~new_n14174 ;
  assign li0027 = ~new_n14200 ;
  assign li0028 = ~new_n14227 ;
  assign li0029 = ~new_n14253 ;
  assign li0030 = ~new_n14280 ;
  assign li0031 = ~new_n14306 ;
  assign li0032 = ~new_n14333 ;
  assign li0033 = ~new_n14359 ;
  assign li0034 = ~new_n14386 ;
  assign li0035 = ~new_n14412 ;
  assign li0036 = ~new_n14439 ;
  assign li0037 = ~new_n14465 ;
  assign li0038 = ~new_n14492 ;
  assign li0039 = ~new_n14518 ;
  assign li0040 = ~new_n14545 ;
  assign li0041 = ~new_n14571 ;
  assign li0042 = ~new_n14598 ;
  assign li0043 = ~new_n14629 ;
  assign li0044 = ~new_n14634 ;
  assign li0045 = ~new_n14641 ;
  assign li0046 = ~new_n14651 ;
  assign li0047 = new_n14657 ;
  assign li0048 = ~new_n14660 ;
  assign li0049 = ~new_n14665 ;
  assign li0050 = new_n14667 ;
  assign li0051 = ~new_n14675 ;
  assign li0052 = ~new_n14683 ;
  assign li0053 = ~new_n14686 ;
  assign li0054 = ~new_n14689 ;
  assign li0055 = ~new_n14692 ;
  assign li0056 = ~new_n14695 ;
  assign li0057 = ~new_n14698 ;
  assign li0058 = ~new_n14702 ;
  assign li0059 = ~new_n14705 ;
  assign li0060 = ~new_n14708 ;
  assign li0061 = ~new_n14711 ;
  assign li0062 = ~new_n14714 ;
  assign li0063 = ~new_n14717 ;
  assign li0064 = ~new_n14720 ;
  assign li0065 = ~new_n14723 ;
  assign li0066 = ~new_n14726 ;
  assign li0067 = ~new_n14734 ;
  assign li0068 = ~new_n14770 ;
  assign li0069 = ~new_n14783 ;
  assign li0070 = ~new_n14801 ;
  assign li0071 = ~new_n14804 ;
  assign li0072 = ~new_n14808 ;
  assign li0073 = ~new_n14817 ;
  assign li0074 = ~new_n14858 ;
  assign li0075 = ~new_n14877 ;
  assign li0076 = ~new_n14894 ;
  assign li0077 = ~new_n14911 ;
  assign li0078 = ~new_n14932 ;
  assign li0079 = ~new_n14951 ;
  assign li0080 = ~new_n14968 ;
  assign li0081 = ~new_n14985 ;
  assign li0082 = ~new_n15005 ;
  assign li0083 = ~new_n15024 ;
  assign li0084 = ~new_n15041 ;
  assign li0085 = ~new_n15058 ;
  assign li0086 = ~new_n15079 ;
  assign li0087 = ~new_n15098 ;
  assign li0088 = ~new_n15115 ;
  assign li0089 = ~new_n15132 ;
  assign li0090 = ~new_n15135 ;
  assign li0091 = ~new_n15140 ;
  assign li0092 = ~new_n15143 ;
  assign li0093 = ~new_n15146 ;
  assign li0094 = ~new_n15172 ;
  assign li0095 = ~new_n15175 ;
  assign li0096 = ~new_n15198 ;
  assign li0097 = ~new_n15221 ;
  assign li0098 = ~new_n15264 ;
  assign li0099 = ~new_n15290 ;
  assign li0100 = ~new_n15315 ;
  assign li0101 = ~new_n15318 ;
  assign li0102 = ~new_n15332 ;
  assign li0103 = ~new_n15340 ;
  assign li0104 = ~new_n15343 ;
  assign li0105 = ~new_n15350 ;
  assign li0106 = ~new_n15355 ;
  assign li0107 = ~new_n15359 ;
  assign li0108 = ~new_n15363 ;
  assign li0109 = ~new_n15371 ;
  assign li0110 = ~new_n15392 ;
  assign li0111 = ~new_n15460 ;
  assign li0112 = ~new_n15493 ;
  assign li0113 = ~new_n15542 ;
  assign li0114 = ~new_n15569 ;
  assign li0115 = ~new_n15572 ;
  assign li0116 = new_n15575 ;
  assign li0117 = ~new_n2261 ;
  assign li0118 = ~new_n13925 ;
  assign li0119 = ~new_n13860 ;
  assign li0120 = ~new_n15610 ;
  assign li0121 = ~new_n15615 ;
  assign li0122 = ~new_n15618 ;
  assign li0123 = ~new_n15624 ;
  assign li0124 = ~new_n15627 ;
  assign li0125 = ~new_n15630 ;
  assign li0126 = ~new_n15633 ;
  assign li0127 = ~new_n15636 ;
  assign li0128 = ~new_n15639 ;
  assign li0129 = ~new_n15653 ;
  assign li0130 = ~new_n15656 ;
  assign li0131 = ~new_n15698 ;
  assign li0132 = ~new_n15725 ;
  assign li0133 = ~new_n15728 ;
  assign li0134 = ~new_n15751 ;
  assign li0135 = ~new_n15773 ;
  assign li0136 = ~new_n15776 ;
  assign li0137 = ~new_n15809 ;
  assign li0138 = ~new_n15834 ;
  assign li0139 = ~new_n15837 ;
  assign li0140 = ~new_n15860 ;
  assign li0141 = ~new_n15882 ;
  assign li0142 = ~new_n15885 ;
  assign li0143 = ~new_n15908 ;
  assign li0144 = ~new_n15930 ;
  assign li0145 = ~new_n15933 ;
  assign li0146 = ~new_n15975 ;
  assign li0147 = ~new_n16000 ;
  assign li0148 = ~new_n16003 ;
  assign li0149 = ~new_n16006 ;
  assign li0150 = ~new_n16009 ;
  assign li0151 = ~new_n16012 ;
  assign li0152 = ~new_n16054 ;
  assign li0153 = ~new_n16081 ;
  assign li0154 = ~new_n16084 ;
  assign li0155 = ~new_n16107 ;
  assign li0156 = ~new_n16129 ;
  assign li0157 = ~new_n16132 ;
  assign li0158 = ~new_n16155 ;
  assign li0159 = ~new_n16177 ;
  assign li0160 = ~new_n16180 ;
  assign li0161 = ~new_n16183 ;
  assign li0162 = ~new_n16186 ;
  assign li0163 = ~new_n16189 ;
  assign li0164 = ~new_n16231 ;
  assign li0165 = ~new_n16256 ;
  assign li0166 = ~new_n16259 ;
  assign li0167 = ~new_n16301 ;
  assign li0168 = ~new_n16328 ;
  assign li0169 = ~new_n16331 ;
  assign li0170 = ~new_n16373 ;
  assign li0171 = ~new_n16400 ;
  assign li0172 = ~new_n16403 ;
  assign li0173 = ~new_n16445 ;
  assign li0174 = ~new_n16472 ;
  assign li0175 = ~new_n16498 ;
  assign li0176 = ~new_n16502 ;
  assign li0177 = ~new_n16506 ;
  assign li0178 = ~new_n16513 ;
  assign li0179 = ~new_n16529 ;
  assign li0180 = ~new_n16663 ;
  assign li0181 = ~new_n16686 ;
  assign li0182 = ~new_n16690 ;
  assign li0183 = ~new_n16706 ;
  assign li0184 = ~new_n16709 ;
  assign li0185 = ~new_n16725 ;
  assign li0186 = ~new_n16728 ;
  assign li0187 = ~new_n16744 ;
  assign li0188 = ~new_n16747 ;
  assign li0189 = ~new_n16750 ;
  assign li0190 = ~new_n16753 ;
  assign li0191 = ~new_n16756 ;
  assign li0192 = ~new_n16759 ;
  assign li0193 = ~new_n16762 ;
  assign li0194 = ~new_n16765 ;
  assign li0195 = ~new_n16768 ;
  assign li0196 = ~new_n16771 ;
  assign li0197 = ~new_n16774 ;
  assign li0198 = ~new_n16777 ;
  assign li0199 = ~new_n16780 ;
  assign li0200 = ~new_n16783 ;
  assign li0201 = ~new_n16789 ;
  assign li0202 = ~new_n16795 ;
  assign li0203 = ~new_n16801 ;
  assign li0204 = ~new_n16807 ;
  assign li0205 = ~new_n16813 ;
  assign li0206 = ~new_n16819 ;
  assign li0207 = ~new_n16825 ;
  assign li0208 = ~new_n16831 ;
  assign li0209 = ~new_n16837 ;
  assign li0210 = ~new_n16843 ;
  assign li0211 = ~new_n16849 ;
  assign li0212 = ~new_n16855 ;
  assign li0213 = ~new_n16861 ;
  assign li0214 = ~new_n16867 ;
  assign li0215 = ~new_n16873 ;
  assign li0216 = ~new_n16879 ;
  assign li0217 = ~new_n16882 ;
  assign li0218 = ~new_n16885 ;
  assign li0219 = ~new_n16888 ;
  assign li0220 = ~new_n16891 ;
  assign li0221 = ~new_n16894 ;
  assign li0222 = ~new_n16904 ;
  assign li0223 = ~new_n16906 ;
  assign li0224 = ~new_n16909 ;
  assign li0225 = ~new_n16915 ;
  assign li0226 = ~new_n16924 ;
  assign li0227 = ~new_n16930 ;
  assign li0228 = ~new_n16935 ;
  assign li0229 = ~new_n16938 ;
  assign li0230 = ~new_n16944 ;
  assign li0231 = ~new_n16950 ;
  assign li0232 = ~new_n16956 ;
  assign li0233 = ~new_n16962 ;
  assign li0234 = ~new_n16968 ;
  assign li0235 = ~new_n16974 ;
  assign li0236 = ~new_n16980 ;
  assign li0237 = ~new_n16986 ;
  assign li0238 = ~new_n16992 ;
  assign li0239 = ~new_n16998 ;
  assign li0240 = ~new_n17004 ;
  assign li0241 = ~new_n17010 ;
  assign li0242 = ~new_n17016 ;
  assign li0243 = ~new_n17022 ;
  assign li0244 = ~new_n17028 ;
  assign li0245 = ~new_n17034 ;
  assign li0246 = ~new_n17040 ;
  assign li0247 = ~new_n17043 ;
  assign li0248 = ~new_n17054 ;
  assign li0249 = ~new_n17057 ;
  assign li0250 = ~new_n17060 ;
  assign li0251 = ~new_n17063 ;
  assign li0252 = ~new_n17066 ;
  assign li0253 = ~new_n17073 ;
  assign li0254 = ~new_n17078 ;
  assign li0255 = ~new_n17082 ;
  assign li0256 = ~new_n17108 ;
  assign li0257 = ~new_n17111 ;
  assign li0258 = ~new_n17117 ;
  assign li0259 = ~new_n17123 ;
  assign li0260 = ~new_n17129 ;
  assign li0261 = ~new_n17135 ;
  assign li0262 = ~new_n17141 ;
  assign li0263 = ~new_n17147 ;
  assign li0264 = ~new_n17153 ;
  assign li0265 = ~new_n17159 ;
  assign li0266 = ~new_n17165 ;
  assign li0267 = ~new_n17171 ;
  assign li0268 = ~new_n17177 ;
  assign li0269 = ~new_n17183 ;
  assign li0270 = ~new_n17189 ;
  assign li0271 = ~new_n17195 ;
  assign li0272 = ~new_n17201 ;
  assign li0273 = ~new_n17207 ;
  assign li0274 = ~new_n17210 ;
  assign li0275 = ~new_n17216 ;
  assign li0276 = ~new_n17222 ;
  assign li0277 = ~new_n17226 ;
  assign li0278 = ~new_n17232 ;
  assign li0279 = ~new_n17238 ;
  assign li0280 = ~new_n17244 ;
  assign li0281 = ~new_n17250 ;
  assign li0282 = ~new_n17256 ;
  assign li0283 = ~new_n17262 ;
  assign li0284 = ~new_n17268 ;
  assign li0285 = ~new_n17274 ;
  assign li0286 = ~new_n17280 ;
  assign li0287 = ~new_n17286 ;
  assign li0288 = ~new_n17292 ;
  assign li0289 = ~new_n17298 ;
  assign li0290 = ~new_n17304 ;
  assign li0291 = ~new_n17310 ;
  assign li0292 = ~new_n17316 ;
  assign li0293 = ~new_n17322 ;
  assign li0294 = ~new_n17328 ;
  assign li0295 = ~new_n17334 ;
  assign li0296 = ~new_n17337 ;
  assign li0297 = ~new_n17343 ;
  assign li0298 = ~new_n17351 ;
  assign li0299 = ~new_n17364 ;
  assign li0300 = ~new_n17368 ;
  assign li0301 = ~new_n17374 ;
  assign li0302 = ~new_n17380 ;
  assign li0303 = ~new_n17386 ;
  assign li0304 = ~new_n17392 ;
  assign li0305 = ~new_n17398 ;
  assign li0306 = ~new_n17404 ;
  assign li0307 = ~new_n17410 ;
  assign li0308 = ~new_n17416 ;
  assign li0309 = ~new_n17422 ;
  assign li0310 = ~new_n17428 ;
  assign li0311 = ~new_n17434 ;
  assign li0312 = ~new_n17440 ;
  assign li0313 = ~new_n17446 ;
  assign li0314 = ~new_n17452 ;
  assign li0315 = ~new_n17458 ;
  assign li0316 = ~new_n17464 ;
  assign li0317 = ~new_n17467 ;
  assign li0318 = ~new_n17473 ;
  assign li0319 = ~new_n17479 ;
  assign li0320 = ~new_n17482 ;
  assign li0321 = ~new_n17485 ;
  assign li0322 = ~new_n17491 ;
  assign li0323 = ~new_n17497 ;
  assign li0324 = ~new_n17503 ;
  assign li0325 = ~new_n17509 ;
  assign li0326 = ~new_n17515 ;
  assign li0327 = ~new_n17521 ;
  assign li0328 = ~new_n17527 ;
  assign li0329 = ~new_n17533 ;
  assign li0330 = ~new_n17539 ;
  assign li0331 = ~new_n17545 ;
  assign li0332 = ~new_n17551 ;
  assign li0333 = ~new_n17557 ;
  assign li0334 = ~new_n17563 ;
  assign li0335 = ~new_n17569 ;
  assign li0336 = ~new_n17575 ;
  assign li0337 = ~new_n17581 ;
  assign li0338 = ~new_n17584 ;
  assign li0339 = ~new_n17590 ;
  assign li0340 = ~new_n17596 ;
  assign li0341 = ~new_n17599 ;
  assign li0342 = ~new_n17605 ;
  assign li0343 = ~new_n17611 ;
  assign li0344 = ~new_n17617 ;
  assign li0345 = ~new_n17623 ;
  assign li0346 = ~new_n17629 ;
  assign li0347 = ~new_n17635 ;
  assign li0348 = ~new_n17641 ;
  assign li0349 = ~new_n17647 ;
  assign li0350 = ~new_n17653 ;
  assign li0351 = ~new_n17659 ;
  assign li0352 = ~new_n17665 ;
  assign li0353 = ~new_n17671 ;
  assign li0354 = ~new_n17677 ;
  assign li0355 = ~new_n17683 ;
  assign li0356 = ~new_n17689 ;
  assign li0357 = ~new_n17695 ;
  assign li0358 = ~new_n17701 ;
  assign li0359 = ~new_n17704 ;
  assign li0360 = ~new_n17712 ;
  assign li0361 = ~new_n17718 ;
  assign li0362 = ~new_n17724 ;
  assign li0363 = ~new_n17730 ;
  assign li0364 = ~new_n17736 ;
  assign li0365 = ~new_n17742 ;
  assign li0366 = ~new_n17748 ;
  assign li0367 = ~new_n17754 ;
  assign li0368 = ~new_n17760 ;
  assign li0369 = ~new_n17766 ;
  assign li0370 = ~new_n17772 ;
  assign li0371 = ~new_n17778 ;
  assign li0372 = ~new_n17784 ;
  assign li0373 = ~new_n17790 ;
  assign li0374 = ~new_n17796 ;
  assign li0375 = ~new_n17802 ;
  assign li0376 = ~new_n17808 ;
  assign li0377 = ~new_n17811 ;
  assign li0378 = ~new_n17817 ;
  assign li0379 = ~new_n17823 ;
  assign li0380 = ~new_n17826 ;
  assign li0381 = ~new_n17829 ;
  assign li0382 = ~new_n17835 ;
  assign li0383 = ~new_n17841 ;
  assign li0384 = ~new_n17847 ;
  assign li0385 = ~new_n17853 ;
  assign li0386 = ~new_n17859 ;
  assign li0387 = ~new_n17865 ;
  assign li0388 = ~new_n17871 ;
  assign li0389 = ~new_n17877 ;
  assign li0390 = ~new_n17883 ;
  assign li0391 = ~new_n17889 ;
  assign li0392 = ~new_n17895 ;
  assign li0393 = ~new_n17901 ;
  assign li0394 = ~new_n17907 ;
  assign li0395 = ~new_n17913 ;
  assign li0396 = ~new_n17919 ;
  assign li0397 = ~new_n17925 ;
  assign li0398 = ~new_n17928 ;
  assign li0399 = ~new_n17937 ;
  assign li0400 = ~new_n17943 ;
  assign li0401 = ~new_n17949 ;
  assign li0402 = ~new_n17955 ;
  assign li0403 = ~new_n17961 ;
  assign li0404 = ~new_n17967 ;
  assign li0405 = ~new_n17973 ;
  assign li0406 = ~new_n17979 ;
  assign li0407 = ~new_n17985 ;
  assign li0408 = ~new_n17991 ;
  assign li0409 = ~new_n17997 ;
  assign li0410 = ~new_n18003 ;
  assign li0411 = ~new_n18009 ;
  assign li0412 = ~new_n18015 ;
  assign li0413 = ~new_n18021 ;
  assign li0414 = ~new_n18027 ;
  assign li0415 = ~new_n18033 ;
  assign li0416 = ~new_n18039 ;
  assign li0417 = ~new_n18045 ;
  assign li0418 = ~new_n18051 ;
  assign li0419 = ~new_n18057 ;
  assign li0420 = ~new_n18063 ;
  assign li0421 = ~new_n18069 ;
  assign li0422 = ~new_n18075 ;
  assign li0423 = ~new_n18081 ;
  assign li0424 = ~new_n18087 ;
  assign li0425 = ~new_n18093 ;
  assign li0426 = ~new_n18099 ;
  assign li0427 = ~new_n18105 ;
  assign li0428 = ~new_n18111 ;
  assign li0429 = ~new_n18117 ;
  assign li0430 = ~new_n18123 ;
  assign li0431 = ~new_n18129 ;
  assign li0432 = ~new_n18135 ;
  assign li0433 = ~new_n18141 ;
  assign li0434 = ~new_n18147 ;
  assign li0435 = ~new_n18150 ;
  assign li0436 = ~new_n18153 ;
  assign li0437 = ~new_n18159 ;
  assign li0438 = ~new_n18165 ;
  assign li0439 = ~new_n18168 ;
  assign li0440 = ~new_n18174 ;
  assign li0441 = ~new_n18180 ;
  assign li0442 = ~new_n18186 ;
  assign li0443 = ~new_n18192 ;
  assign li0444 = ~new_n18198 ;
  assign li0445 = ~new_n18204 ;
  assign li0446 = ~new_n18210 ;
  assign li0447 = ~new_n18216 ;
  assign li0448 = ~new_n18222 ;
  assign li0449 = ~new_n18228 ;
  assign li0450 = ~new_n18234 ;
  assign li0451 = ~new_n18240 ;
  assign li0452 = ~new_n18246 ;
  assign li0453 = ~new_n18252 ;
  assign li0454 = ~new_n18258 ;
  assign li0455 = ~new_n18264 ;
  assign li0456 = ~new_n18267 ;
  assign li0457 = ~new_n18273 ;
  assign li0458 = ~new_n18279 ;
  assign li0459 = ~new_n18282 ;
  assign li0460 = ~new_n18288 ;
  assign li0461 = ~new_n18294 ;
  assign li0462 = ~new_n18300 ;
  assign li0463 = ~new_n18306 ;
  assign li0464 = ~new_n18312 ;
  assign li0465 = ~new_n18318 ;
  assign li0466 = ~new_n18324 ;
  assign li0467 = ~new_n18330 ;
  assign li0468 = ~new_n18336 ;
  assign li0469 = ~new_n18342 ;
  assign li0470 = ~new_n18348 ;
  assign li0471 = ~new_n18354 ;
  assign li0472 = ~new_n18360 ;
  assign li0473 = ~new_n18366 ;
  assign li0474 = ~new_n18372 ;
  assign li0475 = ~new_n18378 ;
  assign li0476 = ~new_n18384 ;
  assign li0477 = ~new_n18390 ;
  assign li0478 = ~new_n18393 ;
  assign li0479 = ~new_n18399 ;
  assign li0480 = ~new_n18405 ;
  assign li0481 = ~new_n18411 ;
  assign li0482 = ~new_n18417 ;
  assign li0483 = ~new_n18423 ;
  assign li0484 = ~new_n18429 ;
  assign li0485 = ~new_n18435 ;
  assign li0486 = ~new_n18441 ;
  assign li0487 = ~new_n18447 ;
  assign li0488 = ~new_n18453 ;
  assign li0489 = ~new_n18459 ;
  assign li0490 = ~new_n18465 ;
  assign li0491 = ~new_n18471 ;
  assign li0492 = ~new_n18477 ;
  assign li0493 = ~new_n18483 ;
  assign li0494 = ~new_n18489 ;
  assign li0495 = ~new_n18495 ;
  assign li0496 = ~new_n18501 ;
  assign li0497 = ~new_n18504 ;
  assign li0498 = ~new_n18510 ;
  assign li0499 = ~new_n18516 ;
  assign li0500 = ~new_n18522 ;
  assign li0501 = ~new_n18528 ;
  assign li0502 = ~new_n18534 ;
  assign li0503 = ~new_n18540 ;
  assign li0504 = ~new_n18546 ;
  assign li0505 = ~new_n18552 ;
  assign li0506 = ~new_n18558 ;
  assign li0507 = ~new_n18564 ;
  assign li0508 = ~new_n18570 ;
  assign li0509 = ~new_n18576 ;
  assign li0510 = ~new_n18582 ;
  assign li0511 = ~new_n18588 ;
  assign li0512 = ~new_n18594 ;
  assign li0513 = ~new_n18600 ;
  assign li0514 = ~new_n18603 ;
  assign li0515 = ~new_n18609 ;
  assign li0516 = ~new_n18618 ;
  assign li0517 = ~new_n18621 ;
  assign li0518 = ~new_n18627 ;
  assign li0519 = ~new_n18633 ;
  assign li0520 = ~new_n18639 ;
  assign li0521 = ~new_n18645 ;
  assign li0522 = ~new_n18651 ;
  assign li0523 = ~new_n18657 ;
  assign li0524 = ~new_n18663 ;
  assign li0525 = ~new_n18669 ;
  assign li0526 = ~new_n18675 ;
  assign li0527 = ~new_n18681 ;
  assign li0528 = ~new_n18687 ;
  assign li0529 = ~new_n18693 ;
  assign li0530 = ~new_n18699 ;
  assign li0531 = ~new_n18705 ;
  assign li0532 = ~new_n18711 ;
  assign li0533 = ~new_n18717 ;
  assign li0534 = ~new_n18720 ;
  assign li0535 = ~new_n18726 ;
  assign li0536 = ~new_n18732 ;
  assign li0537 = ~new_n18735 ;
  assign li0538 = ~new_n18738 ;
  assign li0539 = ~new_n18744 ;
  assign li0540 = ~new_n18750 ;
  assign li0541 = ~new_n18756 ;
  assign li0542 = ~new_n18762 ;
  assign li0543 = ~new_n18768 ;
  assign li0544 = ~new_n18774 ;
  assign li0545 = ~new_n18780 ;
  assign li0546 = ~new_n18786 ;
  assign li0547 = ~new_n18792 ;
  assign li0548 = ~new_n18798 ;
  assign li0549 = ~new_n18804 ;
  assign li0550 = ~new_n18810 ;
  assign li0551 = ~new_n18816 ;
  assign li0552 = ~new_n18822 ;
  assign li0553 = ~new_n18828 ;
  assign li0554 = ~new_n18834 ;
  assign li0555 = ~new_n18837 ;
  assign li0556 = ~new_n18843 ;
  assign li0557 = ~new_n18849 ;
  assign li0558 = ~new_n18852 ;
  assign li0559 = ~new_n18855 ;
  assign li0560 = ~new_n18867 ;
  assign li0561 = ~new_n18873 ;
  assign li0562 = ~new_n18879 ;
  assign li0563 = ~new_n18885 ;
  assign li0564 = ~new_n18891 ;
  assign li0565 = ~new_n18897 ;
  assign li0566 = ~new_n18903 ;
  assign li0567 = ~new_n18909 ;
  assign li0568 = ~new_n18915 ;
  assign li0569 = ~new_n18921 ;
  assign li0570 = ~new_n18927 ;
  assign li0571 = ~new_n18933 ;
  assign li0572 = ~new_n18939 ;
  assign li0573 = ~new_n18945 ;
  assign li0574 = ~new_n18951 ;
  assign li0575 = ~new_n18957 ;
  assign li0576 = ~new_n18960 ;
  assign li0577 = ~new_n18963 ;
  assign li0578 = ~new_n18966 ;
  assign li0579 = ~new_n18969 ;
  assign li0580 = ~new_n18978 ;
  assign li0581 = ~new_n18981 ;
  assign li0582 = ~new_n18987 ;
  assign li0583 = ~new_n18993 ;
  assign li0584 = ~new_n18999 ;
  assign li0585 = ~new_n19005 ;
  assign li0586 = ~new_n19011 ;
  assign li0587 = ~new_n19017 ;
  assign li0588 = ~new_n19023 ;
  assign li0589 = ~new_n19029 ;
  assign li0590 = ~new_n19035 ;
  assign li0591 = ~new_n19041 ;
  assign li0592 = ~new_n19047 ;
  assign li0593 = ~new_n19053 ;
  assign li0594 = ~new_n19059 ;
  assign li0595 = ~new_n19065 ;
  assign li0596 = ~new_n19071 ;
  assign li0597 = ~new_n19077 ;
  assign li0598 = ~new_n19083 ;
  assign li0599 = ~new_n19086 ;
  assign li0600 = ~new_n19095 ;
  assign li0601 = ~new_n19098 ;
  assign li0602 = ~new_n19104 ;
  assign li0603 = ~new_n19110 ;
  assign li0604 = ~new_n19116 ;
  assign li0605 = ~new_n19122 ;
  assign li0606 = ~new_n19128 ;
  assign li0607 = ~new_n19134 ;
  assign li0608 = ~new_n19140 ;
  assign li0609 = ~new_n19146 ;
  assign li0610 = ~new_n19152 ;
  assign li0611 = ~new_n19158 ;
  assign li0612 = ~new_n19164 ;
  assign li0613 = ~new_n19170 ;
  assign li0614 = ~new_n19176 ;
  assign li0615 = ~new_n19182 ;
  assign li0616 = ~new_n19188 ;
  assign li0617 = ~new_n19194 ;
  assign li0618 = ~new_n19200 ;
  assign li0619 = ~new_n19206 ;
  assign li0620 = ~new_n19212 ;
  assign li0621 = ~new_n19215 ;
  assign li0622 = ~new_n19227 ;
  assign li0623 = ~new_n19233 ;
  assign li0624 = ~new_n19239 ;
  assign li0625 = ~new_n19245 ;
  assign li0626 = ~new_n19251 ;
  assign li0627 = ~new_n19257 ;
  assign li0628 = ~new_n19263 ;
  assign li0629 = ~new_n19269 ;
  assign li0630 = ~new_n19275 ;
  assign li0631 = ~new_n19281 ;
  assign li0632 = ~new_n19287 ;
  assign li0633 = ~new_n19293 ;
  assign li0634 = ~new_n19299 ;
  assign li0635 = ~new_n19305 ;
  assign li0636 = ~new_n19311 ;
  assign li0637 = ~new_n19317 ;
  assign li0638 = ~new_n19320 ;
  assign li0639 = ~new_n19323 ;
  assign li0640 = ~new_n19326 ;
  assign li0641 = ~new_n19329 ;
  assign li0642 = ~new_n19338 ;
  assign li0643 = ~new_n19341 ;
  assign li0644 = ~new_n19347 ;
  assign li0645 = ~new_n19353 ;
  assign li0646 = ~new_n19359 ;
  assign li0647 = ~new_n19365 ;
  assign li0648 = ~new_n19371 ;
  assign li0649 = ~new_n19377 ;
  assign li0650 = ~new_n19383 ;
  assign li0651 = ~new_n19389 ;
  assign li0652 = ~new_n19395 ;
  assign li0653 = ~new_n19401 ;
  assign li0654 = ~new_n19407 ;
  assign li0655 = ~new_n19413 ;
  assign li0656 = ~new_n19419 ;
  assign li0657 = ~new_n19425 ;
  assign li0658 = ~new_n19431 ;
  assign li0659 = ~new_n19437 ;
  assign li0660 = ~new_n19443 ;
  assign li0661 = ~new_n19449 ;
  assign li0662 = ~new_n19455 ;
  assign li0663 = ~new_n19458 ;
  assign li0664 = ~new_n19464 ;
  assign li0665 = ~new_n19470 ;
  assign li0666 = ~new_n19476 ;
  assign li0667 = ~new_n19482 ;
  assign li0668 = ~new_n19488 ;
  assign li0669 = ~new_n19494 ;
  assign li0670 = ~new_n19500 ;
  assign li0671 = ~new_n19506 ;
  assign li0672 = ~new_n19512 ;
  assign li0673 = ~new_n19518 ;
  assign li0674 = ~new_n19524 ;
  assign li0675 = ~new_n19530 ;
  assign li0676 = ~new_n19536 ;
  assign li0677 = ~new_n19542 ;
  assign li0678 = ~new_n19548 ;
  assign li0679 = ~new_n19554 ;
  assign li0680 = ~new_n19560 ;
  assign li0681 = ~new_n19566 ;
  assign li0682 = ~new_n19569 ;
  assign li0683 = ~new_n19575 ;
  assign li0684 = ~new_n19581 ;
  assign li0685 = ~new_n19587 ;
  assign li0686 = ~new_n19593 ;
  assign li0687 = ~new_n19599 ;
  assign li0688 = ~new_n19605 ;
  assign li0689 = ~new_n19611 ;
  assign li0690 = ~new_n19617 ;
  assign li0691 = ~new_n19623 ;
  assign li0692 = ~new_n19629 ;
  assign li0693 = ~new_n19635 ;
  assign li0694 = ~new_n19641 ;
  assign li0695 = ~new_n19647 ;
  assign li0696 = ~new_n19653 ;
  assign li0697 = ~new_n19659 ;
  assign li0698 = ~new_n19662 ;
  assign li0699 = ~new_n19668 ;
  assign li0700 = ~new_n19674 ;
  assign li0701 = ~new_n19677 ;
  assign li0702 = ~new_n19683 ;
  assign li0703 = ~new_n19689 ;
  assign li0704 = ~new_n19695 ;
  assign li0705 = ~new_n19701 ;
  assign li0706 = ~new_n19707 ;
  assign li0707 = ~new_n19713 ;
  assign li0708 = ~new_n19719 ;
  assign li0709 = ~new_n19725 ;
  assign li0710 = ~new_n19731 ;
  assign li0711 = ~new_n19737 ;
  assign li0712 = ~new_n19743 ;
  assign li0713 = ~new_n19749 ;
  assign li0714 = ~new_n19755 ;
  assign li0715 = ~new_n19761 ;
  assign li0716 = ~new_n19767 ;
  assign li0717 = ~new_n19773 ;
  assign li0718 = ~new_n19779 ;
  assign li0719 = ~new_n19782 ;
  assign li0720 = ~new_n19788 ;
  assign li0721 = ~new_n19791 ;
  assign li0722 = ~new_n19797 ;
  assign li0723 = ~new_n19803 ;
  assign li0724 = ~new_n19809 ;
  assign li0725 = ~new_n19815 ;
  assign li0726 = ~new_n19821 ;
  assign li0727 = ~new_n19827 ;
  assign li0728 = ~new_n19833 ;
  assign li0729 = ~new_n19839 ;
  assign li0730 = ~new_n19845 ;
  assign li0731 = ~new_n19851 ;
  assign li0732 = ~new_n19857 ;
  assign li0733 = ~new_n19863 ;
  assign li0734 = ~new_n19869 ;
  assign li0735 = ~new_n19875 ;
  assign li0736 = ~new_n19881 ;
  assign li0737 = ~new_n19887 ;
  assign li0738 = ~new_n19893 ;
  assign li0739 = ~new_n19899 ;
  assign li0740 = ~new_n19905 ;
  assign li0741 = ~new_n19908 ;
  assign li0742 = ~new_n19914 ;
  assign li0743 = ~new_n19920 ;
  assign li0744 = ~new_n19926 ;
  assign li0745 = ~new_n19932 ;
  assign li0746 = ~new_n19938 ;
  assign li0747 = ~new_n19944 ;
  assign li0748 = ~new_n19950 ;
  assign li0749 = ~new_n19956 ;
  assign li0750 = ~new_n19962 ;
  assign li0751 = ~new_n19968 ;
  assign li0752 = ~new_n19974 ;
  assign li0753 = ~new_n19980 ;
  assign li0754 = ~new_n19986 ;
  assign li0755 = ~new_n19992 ;
  assign li0756 = ~new_n19998 ;
  assign li0757 = ~new_n20004 ;
  assign li0758 = ~new_n20007 ;
  assign li0759 = ~new_n20010 ;
  assign li0760 = ~new_n20013 ;
  assign li0761 = ~new_n20019 ;
  assign li0762 = ~new_n20022 ;
  assign li0763 = ~new_n20025 ;
  assign li0764 = ~new_n20031 ;
  assign li0765 = ~new_n20037 ;
  assign li0766 = ~new_n20043 ;
  assign li0767 = ~new_n20049 ;
  assign li0768 = ~new_n20055 ;
  assign li0769 = ~new_n20061 ;
  assign li0770 = ~new_n20067 ;
  assign li0771 = ~new_n20073 ;
  assign li0772 = ~new_n20079 ;
  assign li0773 = ~new_n20085 ;
  assign li0774 = ~new_n20091 ;
  assign li0775 = ~new_n20097 ;
  assign li0776 = ~new_n20103 ;
  assign li0777 = ~new_n20109 ;
  assign li0778 = ~new_n20115 ;
  assign li0779 = ~new_n20121 ;
  assign li0780 = ~new_n20124 ;
  assign li0781 = ~new_n20130 ;
  assign li0782 = ~new_n20136 ;
  assign li0783 = ~new_n20139 ;
  assign li0784 = ~new_n20145 ;
  assign li0785 = ~new_n20151 ;
  assign li0786 = ~new_n20157 ;
  assign li0787 = ~new_n20163 ;
  assign li0788 = ~new_n20169 ;
  assign li0789 = ~new_n20175 ;
  assign li0790 = ~new_n20181 ;
  assign li0791 = ~new_n20187 ;
  assign li0792 = ~new_n20193 ;
  assign li0793 = ~new_n20199 ;
  assign li0794 = ~new_n20205 ;
  assign li0795 = ~new_n20211 ;
  assign li0796 = ~new_n20217 ;
  assign li0797 = ~new_n20223 ;
  assign li0798 = ~new_n20229 ;
  assign li0799 = ~new_n20235 ;
  assign li0800 = ~new_n20238 ;
  assign li0801 = ~new_n20241 ;
  assign li0802 = ~new_n20244 ;
  assign li0803 = ~new_n20250 ;
  assign li0804 = ~new_n20253 ;
  assign li0805 = ~new_n20259 ;
  assign li0806 = ~new_n20265 ;
  assign li0807 = ~new_n20271 ;
  assign li0808 = ~new_n20277 ;
  assign li0809 = ~new_n20283 ;
  assign li0810 = ~new_n20289 ;
  assign li0811 = ~new_n20295 ;
  assign li0812 = ~new_n20301 ;
  assign li0813 = ~new_n20307 ;
  assign li0814 = ~new_n20313 ;
  assign li0815 = ~new_n20319 ;
  assign li0816 = ~new_n20325 ;
  assign li0817 = ~new_n20331 ;
  assign li0818 = ~new_n20337 ;
  assign li0819 = ~new_n20343 ;
  assign li0820 = ~new_n20349 ;
  assign li0821 = ~new_n20355 ;
  assign li0822 = ~new_n20357 ;
  assign li0823 = ~new_n20360 ;
  assign li0824 = ~new_n20366 ;
  assign li0825 = ~new_n20372 ;
  assign li0826 = ~new_n20384 ;
  assign li0827 = ~new_n20390 ;
  assign li0828 = ~new_n20396 ;
  assign li0829 = ~new_n20402 ;
  assign li0830 = ~new_n20408 ;
  assign li0831 = ~new_n20414 ;
  assign li0832 = ~new_n20420 ;
  assign li0833 = ~new_n20426 ;
  assign li0834 = ~new_n20432 ;
  assign li0835 = ~new_n20438 ;
  assign li0836 = ~new_n20444 ;
  assign li0837 = ~new_n20450 ;
  assign li0838 = ~new_n20456 ;
  assign li0839 = ~new_n20462 ;
  assign li0840 = ~new_n20468 ;
  assign li0841 = ~new_n20474 ;
  assign li0842 = ~new_n20480 ;
  assign li0843 = ~new_n20486 ;
  assign li0844 = ~new_n20492 ;
  assign li0845 = ~new_n20495 ;
  assign li0846 = ~new_n20502 ;
  assign li0847 = ~new_n20516 ;
  assign li0848 = ~new_n20525 ;
  assign li0849 = ~new_n20543 ;
  assign li0850 = ~new_n20558 ;
  assign li0851 = ~new_n20562 ;
  assign li0852 = ~new_n20568 ;
  assign li0853 = ~new_n20573 ;
  assign li0854 = ~new_n20578 ;
  assign li0855 = ~new_n20583 ;
  assign li0856 = ~new_n20594 ;
  assign li0857 = ~new_n20598 ;
  assign li0858 = ~new_n20601 ;
  assign li0859 = ~new_n20606 ;
  assign li0860 = ~new_n20609 ;
  assign li0861 = ~new_n20612 ;
  assign li0862 = ~new_n20615 ;
  assign li0863 = ~new_n20618 ;
  assign li0864 = ~new_n20621 ;
  assign li0865 = ~new_n20624 ;
  assign li0866 = ~new_n20627 ;
  assign li0867 = ~new_n20630 ;
  assign li0868 = ~new_n20633 ;
  assign li0869 = ~new_n20636 ;
  assign li0870 = ~new_n20639 ;
  assign li0871 = ~new_n20642 ;
  assign li0872 = ~new_n20669 ;
  assign li0873 = ~new_n20697 ;
  assign li0874 = ~new_n20716 ;
  assign li0875 = ~new_n20732 ;
  assign li0876 = ~new_n20749 ;
  assign li0877 = ~new_n20752 ;
  assign li0878 = ~new_n20755 ;
  assign li0879 = ~new_n20758 ;
  assign li0880 = ~new_n20761 ;
  assign li0881 = ~new_n20766 ;
  assign li0882 = ~new_n20773 ;
  assign li0883 = ~new_n20776 ;
  assign li0884 = ~new_n20779 ;
  assign li0885 = ~new_n20792 ;
  assign li0886 = new_n20802 ;
  assign li0887 = new_n20806 ;
  assign li0888 = new_n20811 ;
  assign li0889 = new_n20812 ;
  assign li0890 = new_n20814 ;
  assign li0891 = new_n20815 ;
  assign li0892 = ~new_n20824 ;
  assign li0893 = ~new_n20833 ;
  assign li0894 = ~pi014 ;
  assign li0895 = ~new_n20861 ;
  assign li0896 = ~new_n20885 ;
  assign li0897 = new_n20887 ;
  assign li0898 = new_n14666 ;
  assign li0899 = new_n14670 ;
  assign li0900 = new_n20890 ;
  assign li0901 = lo0900 ;
  assign li0902 = ~new_n20893 ;
  assign li0903 = ~new_n20896 ;
  assign li0904 = ~new_n20899 ;
  assign li0905 = ~new_n20902 ;
  assign li0906 = ~new_n20905 ;
  assign li0907 = ~new_n20908 ;
  assign li0908 = ~new_n20912 ;
  assign li0909 = ~new_n20915 ;
  assign li0910 = ~new_n20918 ;
  assign li0911 = ~new_n20921 ;
  assign li0912 = ~new_n20924 ;
  assign li0913 = ~new_n20927 ;
  assign li0914 = ~new_n20930 ;
  assign li0915 = ~new_n20933 ;
  assign li0916 = ~new_n20937 ;
  assign li0917 = ~new_n20954 ;
  assign li0918 = ~new_n20959 ;
  assign li0919 = ~new_n20962 ;
  assign li0920 = ~new_n20966 ;
  assign li0921 = ~new_n20969 ;
  assign li0922 = ~new_n20972 ;
  assign li0923 = ~new_n20977 ;
  assign li0924 = ~new_n20982 ;
  assign li0925 = ~new_n20986 ;
  assign li0926 = ~new_n20990 ;
  assign li0927 = ~new_n20993 ;
  assign li0928 = ~new_n20996 ;
  assign li0929 = ~new_n20999 ;
  assign li0930 = ~new_n21002 ;
  assign li0931 = ~new_n21006 ;
  assign li0932 = ~new_n21020 ;
  assign li0933 = new_n21022 ;
  assign li0934 = new_n21024 ;
  assign li0935 = new_n21026 ;
  assign li0936 = new_n21028 ;
  assign li0937 = new_n21030 ;
  assign li0938 = ~new_n21047 ;
  assign li0939 = new_n21050 ;
  assign li0940 = new_n21051 ;
  assign li0941 = new_n21052 ;
  assign li0942 = ~new_n21058 ;
  assign li0943 = ~new_n21063 ;
  assign li0944 = ~new_n21068 ;
  assign li0945 = ~new_n21071 ;
  assign li0946 = ~new_n21076 ;
  assign li0947 = ~new_n21079 ;
  assign li0948 = ~new_n21084 ;
  assign li0949 = ~new_n21087 ;
  assign li0950 = ~new_n21091 ;
  assign li0951 = ~new_n21101 ;
  assign li0952 = ~new_n21104 ;
  assign li0953 = ~new_n21107 ;
  assign li0954 = ~new_n21113 ;
  assign li0955 = ~new_n21122 ;
  assign li0956 = ~new_n21125 ;
  assign li0957 = ~new_n21133 ;
  assign li0958 = ~new_n21184 ;
  assign li0959 = ~new_n21187 ;
  assign li0960 = ~new_n21190 ;
  assign li0961 = ~new_n21193 ;
  assign li0962 = ~new_n21200 ;
  assign li0963 = ~new_n21204 ;
  assign li0964 = ~new_n21207 ;
  assign li0965 = ~new_n21210 ;
  assign li0966 = ~new_n21213 ;
  assign li0967 = ~new_n21216 ;
  assign li0968 = ~new_n21219 ;
  assign li0969 = ~new_n21222 ;
  assign li0970 = ~new_n21225 ;
  assign li0971 = ~new_n21228 ;
  assign li0972 = ~new_n21231 ;
  assign li0973 = ~new_n21234 ;
  assign li0974 = ~new_n21237 ;
  assign li0975 = ~new_n21240 ;
  assign li0976 = ~new_n21243 ;
  assign li0977 = ~new_n21247 ;
  assign li0978 = ~new_n21255 ;
  assign li0979 = ~new_n21258 ;
  assign li0980 = new_n21260 ;
  assign li0981 = ~new_n21263 ;
  assign li0982 = ~new_n21266 ;
  assign li0983 = ~new_n21269 ;
  assign li0984 = ~new_n21272 ;
  assign li0985 = ~new_n21275 ;
  assign li0986 = ~new_n21278 ;
  assign li0987 = ~new_n21281 ;
  assign li0988 = ~new_n21284 ;
  assign li0989 = ~new_n21287 ;
  assign li0990 = ~new_n21290 ;
  assign li0991 = ~new_n21293 ;
  assign li0992 = ~new_n21296 ;
  assign li0993 = ~new_n21299 ;
  assign li0994 = ~new_n21302 ;
  assign li0995 = ~new_n21305 ;
  assign li0996 = ~new_n21308 ;
  assign li0997 = ~new_n21311 ;
  assign li0998 = ~new_n21314 ;
  assign li0999 = ~new_n21317 ;
  assign li1000 = ~new_n21320 ;
  assign li1001 = ~new_n21323 ;
  assign li1002 = ~new_n21326 ;
  assign li1003 = ~new_n21329 ;
  assign li1004 = ~new_n21332 ;
  assign li1005 = ~new_n21335 ;
  assign li1006 = ~new_n21338 ;
  assign li1007 = ~new_n21341 ;
  assign li1008 = ~new_n21344 ;
  assign li1009 = ~new_n21347 ;
  assign li1010 = ~new_n21350 ;
  assign li1011 = ~new_n21353 ;
  assign li1012 = ~new_n21356 ;
  assign li1013 = ~new_n21359 ;
  assign li1014 = ~new_n21362 ;
  assign li1015 = ~new_n21365 ;
  assign li1016 = ~new_n21368 ;
  assign li1017 = ~new_n21371 ;
  assign li1018 = ~new_n21374 ;
  assign li1019 = ~new_n21377 ;
  assign li1020 = ~new_n21380 ;
  assign li1021 = ~new_n21383 ;
  assign li1022 = ~new_n21386 ;
  assign li1023 = ~new_n21389 ;
  assign li1024 = ~new_n21392 ;
  assign li1025 = ~new_n21395 ;
  assign li1026 = ~new_n21398 ;
  assign li1027 = ~new_n21401 ;
  assign li1028 = ~new_n21404 ;
  assign li1029 = ~new_n21407 ;
  assign li1030 = ~new_n21410 ;
  assign li1031 = ~new_n21413 ;
  assign li1032 = ~new_n21416 ;
  assign li1033 = ~new_n21419 ;
  assign li1034 = ~new_n21422 ;
  assign li1035 = ~new_n21425 ;
  assign li1036 = ~new_n21428 ;
  assign li1037 = ~new_n21431 ;
  assign li1038 = ~new_n21434 ;
  assign li1039 = ~new_n21437 ;
  assign li1040 = ~new_n21440 ;
  assign li1041 = ~new_n21443 ;
  assign li1042 = ~new_n21446 ;
  assign li1043 = ~new_n21449 ;
  assign li1044 = ~new_n21452 ;
  assign li1045 = ~new_n21455 ;
  assign li1046 = ~new_n21458 ;
  assign li1047 = ~new_n21461 ;
  assign li1048 = ~new_n21464 ;
  assign li1049 = ~new_n21467 ;
  assign li1050 = ~new_n21470 ;
  assign li1051 = ~new_n21478 ;
  assign li1052 = ~new_n21506 ;
  assign li1053 = ~new_n21529 ;
  assign li1054 = ~new_n21552 ;
  assign li1055 = ~new_n21575 ;
  assign li1056 = ~new_n21592 ;
  assign li1057 = ~new_n21610 ;
  assign li1058 = ~new_n21628 ;
  assign li1059 = ~new_n21645 ;
  assign li1060 = ~new_n21663 ;
  assign li1061 = ~new_n21686 ;
  assign li1062 = ~new_n21690 ;
  assign li1063 = ~new_n21693 ;
  assign li1064 = ~new_n21696 ;
  assign li1065 = ~new_n21699 ;
  assign li1066 = ~new_n21713 ;
  assign li1067 = ~new_n21716 ;
  assign li1068 = ~new_n21724 ;
  assign li1069 = ~new_n21745 ;
  assign li1070 = ~new_n21749 ;
  assign li1071 = ~new_n21754 ;
  assign li1072 = ~new_n21758 ;
  assign li1073 = ~new_n21762 ;
  assign li1074 = new_n21793 ;
  assign li1075 = lo1074 ;
  assign li1076 = ~new_n21835 ;
  assign li1077 = ~new_n21839 ;
  assign li1078 = ~new_n21862 ;
  assign li1079 = ~new_n21865 ;
  assign li1080 = ~new_n21868 ;
  assign li1081 = ~new_n21871 ;
  assign li1082 = ~new_n21874 ;
  assign li1083 = ~new_n21877 ;
  assign li1084 = ~new_n21880 ;
  assign li1085 = ~new_n21883 ;
  assign li1086 = ~new_n21886 ;
  assign li1087 = ~new_n21889 ;
  assign li1088 = ~new_n21892 ;
  assign li1089 = ~new_n21895 ;
  assign li1090 = ~new_n21898 ;
  assign li1091 = ~new_n21901 ;
  assign li1092 = new_n21248 ;
  assign li1093 = ~new_n21924 ;
  assign li1094 = ~new_n21947 ;
  assign li1095 = ~new_n21950 ;
  assign li1096 = ~new_n21953 ;
  assign li1097 = ~new_n21956 ;
  assign li1098 = ~new_n21959 ;
  assign li1099 = ~new_n21962 ;
  assign li1100 = ~new_n21965 ;
  assign li1101 = ~new_n21975 ;
  assign li1102 = ~new_n21996 ;
  assign li1103 = ~new_n21999 ;
  assign li1104 = ~new_n22002 ;
  assign li1105 = ~new_n22005 ;
  assign li1106 = ~new_n22008 ;
  assign li1107 = ~new_n22011 ;
  assign li1108 = ~new_n22013 ;
  assign li1109 = new_n22014 ;
  assign li1110 = pi016 ;
  assign li1111 = lo1110 ;
  assign li1112 = ~new_n22026 ;
  assign li1113 = ~new_n22032 ;
  assign li1114 = ~new_n22045 ;
  assign li1115 = ~new_n22049 ;
  assign li1116 = ~new_n22054 ;
  assign li1117 = ~new_n22057 ;
  assign li1118 = ~new_n22060 ;
  assign li1119 = ~new_n22063 ;
  assign li1120 = ~new_n22066 ;
  assign li1121 = ~new_n22075 ;
  assign li1122 = ~new_n22084 ;
  assign li1123 = ~new_n22093 ;
  assign li1124 = ~new_n22096 ;
  assign li1125 = ~new_n22105 ;
  assign li1126 = ~new_n22114 ;
  assign li1127 = ~new_n22117 ;
  assign li1128 = ~new_n22129 ;
  assign li1129 = ~new_n22139 ;
  assign li1130 = ~new_n22142 ;
  assign li1131 = ~new_n22146 ;
  assign li1132 = ~new_n22149 ;
  assign li1133 = ~new_n22153 ;
  assign li1134 = ~new_n22164 ;
  assign li1135 = ~new_n22167 ;
  assign li1136 = ~new_n22188 ;
  assign li1137 = ~new_n22191 ;
  assign li1138 = ~new_n22194 ;
  assign li1139 = ~new_n22197 ;
  assign li1140 = ~new_n22200 ;
  assign li1141 = ~new_n22203 ;
  assign li1142 = new_n22234 ;
  assign li1143 = ~lo1236 ;
  assign li1144 = lo1143 ;
  assign li1145 = ~new_n22238 ;
  assign li1146 = ~new_n22241 ;
  assign li1147 = ~new_n22250 ;
  assign li1148 = ~new_n22253 ;
  assign li1149 = ~new_n22262 ;
  assign li1150 = ~new_n22265 ;
  assign li1151 = ~new_n22274 ;
  assign li1152 = ~new_n22277 ;
  assign li1153 = ~new_n22286 ;
  assign li1154 = ~new_n22289 ;
  assign li1155 = ~new_n22298 ;
  assign li1156 = ~new_n22301 ;
  assign li1157 = ~new_n22310 ;
  assign li1158 = ~new_n22313 ;
  assign li1159 = ~new_n22322 ;
  assign li1160 = ~new_n22325 ;
  assign li1161 = ~new_n22334 ;
  assign li1162 = ~new_n22337 ;
  assign li1163 = ~new_n22346 ;
  assign li1164 = ~new_n22349 ;
  assign li1165 = ~new_n22358 ;
  assign li1166 = ~new_n22361 ;
  assign li1167 = ~new_n22370 ;
  assign li1168 = ~new_n22373 ;
  assign li1169 = ~new_n22382 ;
  assign li1170 = ~new_n22385 ;
  assign li1171 = ~new_n22394 ;
  assign li1172 = ~new_n22397 ;
  assign li1173 = ~new_n22406 ;
  assign li1174 = ~new_n22409 ;
  assign li1175 = ~new_n22418 ;
  assign li1176 = ~new_n22421 ;
  assign li1177 = ~new_n22430 ;
  assign li1178 = ~new_n22433 ;
  assign li1179 = ~new_n22442 ;
  assign li1180 = ~new_n22445 ;
  assign li1181 = ~new_n22454 ;
  assign li1182 = ~new_n22457 ;
  assign li1183 = ~new_n22466 ;
  assign li1184 = ~new_n22469 ;
  assign li1185 = ~new_n22478 ;
  assign li1186 = ~new_n22481 ;
  assign li1187 = ~new_n22490 ;
  assign li1188 = ~new_n22493 ;
  assign li1189 = ~new_n22502 ;
  assign li1190 = ~new_n22505 ;
  assign li1191 = ~new_n22514 ;
  assign li1192 = ~new_n22517 ;
  assign li1193 = ~new_n22526 ;
  assign li1194 = ~new_n22529 ;
  assign li1195 = ~new_n22538 ;
  assign li1196 = ~new_n22541 ;
  assign li1197 = ~new_n22550 ;
  assign li1198 = ~new_n22553 ;
  assign li1199 = ~new_n22562 ;
  assign li1200 = ~new_n22565 ;
  assign li1201 = ~new_n22574 ;
  assign li1202 = ~new_n22583 ;
  assign li1203 = ~new_n22592 ;
  assign li1204 = ~new_n22601 ;
  assign li1205 = ~new_n22610 ;
  assign li1206 = ~new_n22619 ;
  assign li1207 = ~new_n22628 ;
  assign li1208 = ~new_n22637 ;
  assign li1209 = ~new_n22646 ;
  assign li1210 = ~new_n22655 ;
  assign li1211 = ~new_n22664 ;
  assign li1212 = ~new_n22673 ;
  assign li1213 = ~new_n22682 ;
  assign li1214 = ~new_n22691 ;
  assign li1215 = ~new_n22700 ;
  assign li1216 = ~new_n22709 ;
  assign li1217 = ~new_n22718 ;
  assign li1218 = ~new_n22727 ;
  assign li1219 = ~new_n22736 ;
  assign li1220 = ~new_n22745 ;
  assign li1221 = ~new_n22754 ;
  assign li1222 = ~new_n22763 ;
  assign li1223 = ~new_n22772 ;
  assign li1224 = ~new_n22781 ;
  assign li1225 = ~new_n22790 ;
  assign li1226 = ~new_n22799 ;
  assign li1227 = ~new_n22808 ;
  assign li1228 = ~new_n22817 ;
  assign li1229 = ~new_n22826 ;
  assign li1230 = ~new_n22847 ;
  assign li1231 = ~new_n22850 ;
  assign li1232 = ~new_n22853 ;
  assign li1233 = ~new_n22856 ;
  assign li1234 = ~new_n22859 ;
  assign li1235 = ~new_n22862 ;
  assign li1236 = ~new_n22866 ;
  assign li1237 = ~new_n22869 ;
  assign li1238 = ~new_n22890 ;
  assign li1239 = ~new_n22893 ;
  assign li1240 = ~new_n22896 ;
  assign li1241 = ~new_n22899 ;
  assign li1242 = ~new_n22902 ;
  assign li1243 = ~new_n22905 ;
  assign li1244 = ~new_n22911 ;
  assign li1245 = lo1255 ;
  assign li1246 = ~new_n22914 ;
  assign li1247 = ~new_n22935 ;
  assign li1248 = ~new_n22938 ;
  assign li1249 = ~new_n22941 ;
  assign li1250 = ~new_n22944 ;
  assign li1251 = ~new_n22947 ;
  assign li1252 = ~new_n22950 ;
  assign li1253 = ~new_n22956 ;
  assign li1254 = ~new_n22960 ;
  assign li1255 = new_n22961 ;
  assign li1256 = ~new_n22980 ;
  assign li1257 = ~new_n22983 ;
  assign li1258 = ~new_n22986 ;
  assign li1259 = ~new_n22989 ;
  assign li1260 = ~new_n22992 ;
  assign li1261 = ~new_n22995 ;
  assign li1262 = ~new_n22998 ;
  assign li1263 = ~new_n23001 ;
  assign li1264 = ~new_n23004 ;
  assign li1265 = ~new_n23007 ;
  assign li1266 = ~new_n23010 ;
  assign li1267 = ~new_n23013 ;
  assign li1268 = ~new_n23023 ;
  assign li1269 = ~new_n23029 ;
  assign li1270 = ~new_n23035 ;
  assign li1271 = ~new_n23041 ;
  assign li1272 = ~new_n23048 ;
  assign li1273 = ~new_n23054 ;
  assign li1274 = ~new_n23060 ;
  assign li1275 = ~new_n23066 ;
  assign li1276 = ~new_n23072 ;
  assign li1277 = ~new_n23078 ;
  assign li1278 = ~new_n23084 ;
  assign li1279 = ~new_n23090 ;
  assign li1280 = ~new_n23101 ;
  assign li1281 = ~new_n23112 ;
  assign li1282 = ~new_n23123 ;
  assign li1283 = ~new_n23134 ;
  assign li1284 = ~new_n23145 ;
  assign li1285 = new_n23158 ;
  assign li1286 = ~new_n23173 ;
  assign li1287 = ~new_n24945 ;
  assign li1288 = ~new_n24951 ;
  assign li1289 = ~new_n25000 ;
  assign li1290 = ~new_n25028 ;
  assign li1291 = new_n25054 ;
  assign li1292 = new_n25058 ;
  assign li1293 = new_n25063 ;
  assign li1294 = new_n25068 ;
  assign li1295 = ~new_n25074 ;
  assign li1296 = ~new_n25091 ;
  assign li1297 = ~new_n25103 ;
  assign li1298 = ~new_n25120 ;
  assign li1299 = ~new_n25135 ;
  assign li1300 = ~new_n25141 ;
  assign li1301 = ~new_n25153 ;
  assign li1302 = ~new_n25170 ;
  assign li1303 = ~new_n25176 ;
  assign li1304 = ~new_n25182 ;
  assign li1305 = ~new_n25188 ;
  assign li1306 = ~new_n25194 ;
  assign li1307 = ~new_n25200 ;
  assign li1308 = ~new_n25206 ;
  assign li1309 = ~new_n25212 ;
  assign li1310 = ~new_n25229 ;
  assign li1311 = ~new_n25246 ;
  assign li1312 = ~new_n25258 ;
  assign li1313 = ~new_n25268 ;
  assign li1314 = ~new_n25274 ;
  assign li1315 = ~new_n25286 ;
  assign li1316 = ~new_n25303 ;
  assign li1317 = ~new_n25309 ;
  assign li1318 = ~new_n25315 ;
  assign li1319 = ~new_n25321 ;
  assign li1320 = ~new_n25327 ;
  assign li1321 = ~new_n25344 ;
  assign li1322 = ~new_n25350 ;
  assign li1323 = ~new_n25367 ;
  assign li1324 = ~new_n25379 ;
  assign li1325 = ~new_n25396 ;
  assign li1326 = ~new_n25408 ;
  assign li1327 = ~new_n25425 ;
  assign li1328 = ~new_n25431 ;
  assign li1329 = ~new_n25437 ;
  assign li1330 = ~new_n25447 ;
  assign li1331 = ~new_n25459 ;
  assign li1332 = ~new_n25476 ;
  assign li1333 = ~new_n25482 ;
  assign li1334 = ~new_n25488 ;
  assign li1335 = ~new_n25505 ;
  assign li1336 = ~new_n25517 ;
  assign li1337 = ~new_n25534 ;
  assign li1338 = ~new_n25551 ;
  assign li1339 = ~new_n25563 ;
  assign li1340 = ~new_n25580 ;
  assign li1341 = ~new_n25590 ;
  assign li1342 = ~new_n25602 ;
  assign li1343 = ~new_n25619 ;
  assign li1344 = ~new_n25625 ;
  assign li1345 = ~new_n25642 ;
  assign li1346 = ~new_n25654 ;
  assign li1347 = ~new_n25671 ;
  assign li1348 = ~new_n25677 ;
  assign li1349 = ~new_n25683 ;
  assign li1350 = ~new_n25689 ;
  assign li1351 = ~new_n25695 ;
  assign li1352 = ~new_n25701 ;
  assign li1353 = ~new_n25711 ;
  assign li1354 = ~new_n25723 ;
  assign li1355 = ~new_n25740 ;
  assign li1356 = ~new_n25750 ;
  assign li1357 = ~new_n25762 ;
  assign li1358 = ~new_n25779 ;
  assign li1359 = ~new_n25785 ;
  assign li1360 = ~new_n25791 ;
  assign li1361 = ~new_n25804 ;
  assign li1362 = ~new_n25837 ;
  assign li1363 = ~new_n25849 ;
  assign li1364 = ~new_n25859 ;
  assign li1365 = ~new_n25871 ;
  assign li1366 = ~new_n25888 ;
  assign li1367 = ~new_n25894 ;
  assign li1368 = ~new_n25911 ;
  assign li1369 = ~new_n25923 ;
  assign li1370 = ~new_n25940 ;
  assign li1371 = ~new_n25950 ;
  assign li1372 = ~new_n25962 ;
  assign li1373 = ~new_n25979 ;
  assign li1374 = ~new_n25996 ;
  assign li1375 = ~new_n26008 ;
  assign li1376 = ~new_n26025 ;
  assign li1377 = ~new_n26035 ;
  assign li1378 = ~new_n26047 ;
  assign li1379 = ~new_n26064 ;
  assign li1380 = ~new_n26070 ;
  assign li1381 = ~new_n26076 ;
  assign li1382 = ~new_n26093 ;
  assign li1383 = ~new_n26110 ;
  assign li1384 = ~new_n26122 ;
  assign li1385 = ~new_n26134 ;
  assign li1386 = ~new_n26151 ;
  assign li1387 = ~new_n26168 ;
  assign li1388 = ~new_n26180 ;
  assign li1389 = ~new_n26190 ;
  assign li1390 = ~new_n26202 ;
  assign li1391 = ~new_n26219 ;
  assign li1392 = ~new_n26225 ;
  assign li1393 = ~new_n26235 ;
  assign li1394 = ~new_n26247 ;
  assign li1395 = ~new_n26264 ;
  assign li1396 = ~new_n26281 ;
  assign li1397 = ~new_n26293 ;
  assign li1398 = ~new_n26310 ;
  assign li1399 = ~new_n26320 ;
  assign li1400 = ~new_n26332 ;
  assign li1401 = ~new_n26349 ;
  assign li1402 = ~new_n26359 ;
  assign li1403 = ~new_n26371 ;
  assign li1404 = ~new_n26388 ;
  assign li1405 = ~new_n26398 ;
  assign li1406 = ~new_n26410 ;
  assign li1407 = ~new_n26427 ;
  assign li1408 = ~new_n26439 ;
  assign li1409 = ~new_n26451 ;
  assign li1410 = ~new_n26467 ;
  assign li1411 = ~new_n26484 ;
  assign li1412 = ~new_n26496 ;
  assign li1413 = ~new_n26513 ;
  assign li1414 = ~new_n26523 ;
  assign li1415 = ~new_n26535 ;
  assign li1416 = ~new_n26552 ;
  assign li1417 = ~new_n26562 ;
  assign li1418 = ~new_n26574 ;
  assign li1419 = ~new_n26591 ;
  assign li1420 = ~new_n26597 ;
  assign li1421 = ~new_n26603 ;
  assign li1422 = ~new_n26609 ;
  assign li1423 = ~new_n26615 ;
  assign li1424 = ~new_n26621 ;
  assign li1425 = ~new_n26628 ;
  assign li1426 = new_n26633 ;
  assign li1427 = new_n26638 ;
  assign li1428 = ~new_n26644 ;
  assign li1429 = new_n26654 ;
  assign li1430 = new_n26661 ;
  assign li1431 = ~new_n26701 ;
  assign li1432 = ~new_n26712 ;
  assign li1433 = ~new_n26718 ;
  assign li1434 = new_n26731 ;
  assign li1435 = ~new_n26742 ;
  assign li1436 = ~new_n26758 ;
  assign li1437 = ~new_n26764 ;
  assign li1438 = ~new_n26770 ;
  assign li1439 = ~new_n26776 ;
  assign li1440 = ~new_n26782 ;
  assign li1441 = ~new_n26789 ;
  assign li1442 = ~new_n26795 ;
  assign li1443 = ~new_n26801 ;
  assign li1444 = ~new_n26812 ;
  assign li1445 = ~new_n26823 ;
  assign li1446 = ~new_n26834 ;
  assign li1447 = ~new_n26841 ;
  assign li1448 = new_n26848 ;
  assign li1449 = ~new_n26855 ;
  assign li1450 = new_n26860 ;
  assign li1451 = ~new_n26866 ;
  assign li1452 = new_n26872 ;
  assign li1453 = new_n26882 ;
  assign li1454 = new_n26886 ;
  assign li1455 = new_n26890 ;
  assign li1456 = new_n26894 ;
  assign li1457 = new_n26898 ;
  assign li1458 = new_n26902 ;
  assign li1459 = new_n26906 ;
  assign li1460 = new_n26911 ;
  assign li1461 = new_n26921 ;
  assign li1462 = new_n26922 ;
  assign li1463 = new_n26926 ;
  assign li1464 = new_n26930 ;
  assign li1465 = new_n26934 ;
  assign li1466 = new_n26938 ;
  assign li1467 = new_n26942 ;
  assign li1468 = new_n26951 ;
  assign li1469 = ~new_n26957 ;
  assign li1470 = ~new_n26963 ;
  assign li1471 = ~new_n26969 ;
  assign li1472 = ~new_n26975 ;
  assign li1473 = ~new_n26981 ;
  assign li1474 = ~new_n26987 ;
  assign li1475 = ~new_n26993 ;
  assign li1476 = ~new_n26999 ;
 always @ (posedge ) begin
    lo0000 <= li0000 ;
 end
 always @ (posedge ) begin
    lo0001 <= li0001 ;
 end
 always @ (posedge ) begin
    lo0002 <= li0002 ;
 end
 always @ (posedge ) begin
    lo0003 <= li0003 ;
 end
 always @ (posedge ) begin
    lo0004 <= li0004 ;
 end
 always @ (posedge ) begin
    lo0005 <= li0005 ;
 end
 always @ (posedge ) begin
    lo0006 <= li0006 ;
 end
 always @ (posedge ) begin
    lo0007 <= li0007 ;
 end
 always @ (posedge ) begin
    lo0008 <= li0008 ;
 end
 always @ (posedge ) begin
    lo0009 <= li0009 ;
 end
 always @ (posedge ) begin
    lo0010 <= li0010 ;
 end
 always @ (posedge ) begin
    lo0011 <= li0011 ;
 end
 always @ (posedge ) begin
    lo0012 <= li0012 ;
 end
 always @ (posedge ) begin
    lo0013 <= li0013 ;
 end
 always @ (posedge ) begin
    lo0014 <= li0014 ;
 end
 always @ (posedge ) begin
    lo0015 <= li0015 ;
 end
 always @ (posedge ) begin
    lo0016 <= li0016 ;
 end
 always @ (posedge ) begin
    lo0017 <= li0017 ;
 end
 always @ (posedge ) begin
    lo0018 <= li0018 ;
 end
 always @ (posedge ) begin
    lo0019 <= li0019 ;
 end
 always @ (posedge ) begin
    lo0020 <= li0020 ;
 end
 always @ (posedge ) begin
    lo0021 <= li0021 ;
 end
 always @ (posedge ) begin
    lo0022 <= li0022 ;
 end
 always @ (posedge ) begin
    lo0023 <= li0023 ;
 end
 always @ (posedge ) begin
    lo0024 <= li0024 ;
 end
 always @ (posedge ) begin
    lo0025 <= li0025 ;
 end
 always @ (posedge ) begin
    lo0026 <= li0026 ;
 end
 always @ (posedge ) begin
    lo0027 <= li0027 ;
 end
 always @ (posedge ) begin
    lo0028 <= li0028 ;
 end
 always @ (posedge ) begin
    lo0029 <= li0029 ;
 end
 always @ (posedge ) begin
    lo0030 <= li0030 ;
 end
 always @ (posedge ) begin
    lo0031 <= li0031 ;
 end
 always @ (posedge ) begin
    lo0032 <= li0032 ;
 end
 always @ (posedge ) begin
    lo0033 <= li0033 ;
 end
 always @ (posedge ) begin
    lo0034 <= li0034 ;
 end
 always @ (posedge ) begin
    lo0035 <= li0035 ;
 end
 always @ (posedge ) begin
    lo0036 <= li0036 ;
 end
 always @ (posedge ) begin
    lo0037 <= li0037 ;
 end
 always @ (posedge ) begin
    lo0038 <= li0038 ;
 end
 always @ (posedge ) begin
    lo0039 <= li0039 ;
 end
 always @ (posedge ) begin
    lo0040 <= li0040 ;
 end
 always @ (posedge ) begin
    lo0041 <= li0041 ;
 end
 always @ (posedge ) begin
    lo0042 <= li0042 ;
 end
 always @ (posedge ) begin
    lo0043 <= li0043 ;
 end
 always @ (posedge ) begin
    lo0044 <= li0044 ;
 end
 always @ (posedge ) begin
    lo0045 <= li0045 ;
 end
 always @ (posedge ) begin
    lo0046 <= li0046 ;
 end
 always @ (posedge ) begin
    lo0047 <= li0047 ;
 end
 always @ (posedge ) begin
    lo0048 <= li0048 ;
 end
 always @ (posedge ) begin
    lo0049 <= li0049 ;
 end
 always @ (posedge ) begin
    lo0050 <= li0050 ;
 end
 always @ (posedge ) begin
    lo0051 <= li0051 ;
 end
 always @ (posedge ) begin
    lo0052 <= li0052 ;
 end
 always @ (posedge ) begin
    lo0053 <= li0053 ;
 end
 always @ (posedge ) begin
    lo0054 <= li0054 ;
 end
 always @ (posedge ) begin
    lo0055 <= li0055 ;
 end
 always @ (posedge ) begin
    lo0056 <= li0056 ;
 end
 always @ (posedge ) begin
    lo0057 <= li0057 ;
 end
 always @ (posedge ) begin
    lo0058 <= li0058 ;
 end
 always @ (posedge ) begin
    lo0059 <= li0059 ;
 end
 always @ (posedge ) begin
    lo0060 <= li0060 ;
 end
 always @ (posedge ) begin
    lo0061 <= li0061 ;
 end
 always @ (posedge ) begin
    lo0062 <= li0062 ;
 end
 always @ (posedge ) begin
    lo0063 <= li0063 ;
 end
 always @ (posedge ) begin
    lo0064 <= li0064 ;
 end
 always @ (posedge ) begin
    lo0065 <= li0065 ;
 end
 always @ (posedge ) begin
    lo0066 <= li0066 ;
 end
 always @ (posedge ) begin
    lo0067 <= li0067 ;
 end
 always @ (posedge ) begin
    lo0068 <= li0068 ;
 end
 always @ (posedge ) begin
    lo0069 <= li0069 ;
 end
 always @ (posedge ) begin
    lo0070 <= li0070 ;
 end
 always @ (posedge ) begin
    lo0071 <= li0071 ;
 end
 always @ (posedge ) begin
    lo0072 <= li0072 ;
 end
 always @ (posedge ) begin
    lo0073 <= li0073 ;
 end
 always @ (posedge ) begin
    lo0074 <= li0074 ;
 end
 always @ (posedge ) begin
    lo0075 <= li0075 ;
 end
 always @ (posedge ) begin
    lo0076 <= li0076 ;
 end
 always @ (posedge ) begin
    lo0077 <= li0077 ;
 end
 always @ (posedge ) begin
    lo0078 <= li0078 ;
 end
 always @ (posedge ) begin
    lo0079 <= li0079 ;
 end
 always @ (posedge ) begin
    lo0080 <= li0080 ;
 end
 always @ (posedge ) begin
    lo0081 <= li0081 ;
 end
 always @ (posedge ) begin
    lo0082 <= li0082 ;
 end
 always @ (posedge ) begin
    lo0083 <= li0083 ;
 end
 always @ (posedge ) begin
    lo0084 <= li0084 ;
 end
 always @ (posedge ) begin
    lo0085 <= li0085 ;
 end
 always @ (posedge ) begin
    lo0086 <= li0086 ;
 end
 always @ (posedge ) begin
    lo0087 <= li0087 ;
 end
 always @ (posedge ) begin
    lo0088 <= li0088 ;
 end
 always @ (posedge ) begin
    lo0089 <= li0089 ;
 end
 always @ (posedge ) begin
    lo0090 <= li0090 ;
 end
 always @ (posedge ) begin
    lo0091 <= li0091 ;
 end
 always @ (posedge ) begin
    lo0092 <= li0092 ;
 end
 always @ (posedge ) begin
    lo0093 <= li0093 ;
 end
 always @ (posedge ) begin
    lo0094 <= li0094 ;
 end
 always @ (posedge ) begin
    lo0095 <= li0095 ;
 end
 always @ (posedge ) begin
    lo0096 <= li0096 ;
 end
 always @ (posedge ) begin
    lo0097 <= li0097 ;
 end
 always @ (posedge ) begin
    lo0098 <= li0098 ;
 end
 always @ (posedge ) begin
    lo0099 <= li0099 ;
 end
 always @ (posedge ) begin
    lo0100 <= li0100 ;
 end
 always @ (posedge ) begin
    lo0101 <= li0101 ;
 end
 always @ (posedge ) begin
    lo0102 <= li0102 ;
 end
 always @ (posedge ) begin
    lo0103 <= li0103 ;
 end
 always @ (posedge ) begin
    lo0104 <= li0104 ;
 end
 always @ (posedge ) begin
    lo0105 <= li0105 ;
 end
 always @ (posedge ) begin
    lo0106 <= li0106 ;
 end
 always @ (posedge ) begin
    lo0107 <= li0107 ;
 end
 always @ (posedge ) begin
    lo0108 <= li0108 ;
 end
 always @ (posedge ) begin
    lo0109 <= li0109 ;
 end
 always @ (posedge ) begin
    lo0110 <= li0110 ;
 end
 always @ (posedge ) begin
    lo0111 <= li0111 ;
 end
 always @ (posedge ) begin
    lo0112 <= li0112 ;
 end
 always @ (posedge ) begin
    lo0113 <= li0113 ;
 end
 always @ (posedge ) begin
    lo0114 <= li0114 ;
 end
 always @ (posedge ) begin
    lo0115 <= li0115 ;
 end
 always @ (posedge ) begin
    lo0116 <= li0116 ;
 end
 always @ (posedge ) begin
    lo0117 <= li0117 ;
 end
 always @ (posedge ) begin
    lo0118 <= li0118 ;
 end
 always @ (posedge ) begin
    lo0119 <= li0119 ;
 end
 always @ (posedge ) begin
    lo0120 <= li0120 ;
 end
 always @ (posedge ) begin
    lo0121 <= li0121 ;
 end
 always @ (posedge ) begin
    lo0122 <= li0122 ;
 end
 always @ (posedge ) begin
    lo0123 <= li0123 ;
 end
 always @ (posedge ) begin
    lo0124 <= li0124 ;
 end
 always @ (posedge ) begin
    lo0125 <= li0125 ;
 end
 always @ (posedge ) begin
    lo0126 <= li0126 ;
 end
 always @ (posedge ) begin
    lo0127 <= li0127 ;
 end
 always @ (posedge ) begin
    lo0128 <= li0128 ;
 end
 always @ (posedge ) begin
    lo0129 <= li0129 ;
 end
 always @ (posedge ) begin
    lo0130 <= li0130 ;
 end
 always @ (posedge ) begin
    lo0131 <= li0131 ;
 end
 always @ (posedge ) begin
    lo0132 <= li0132 ;
 end
 always @ (posedge ) begin
    lo0133 <= li0133 ;
 end
 always @ (posedge ) begin
    lo0134 <= li0134 ;
 end
 always @ (posedge ) begin
    lo0135 <= li0135 ;
 end
 always @ (posedge ) begin
    lo0136 <= li0136 ;
 end
 always @ (posedge ) begin
    lo0137 <= li0137 ;
 end
 always @ (posedge ) begin
    lo0138 <= li0138 ;
 end
 always @ (posedge ) begin
    lo0139 <= li0139 ;
 end
 always @ (posedge ) begin
    lo0140 <= li0140 ;
 end
 always @ (posedge ) begin
    lo0141 <= li0141 ;
 end
 always @ (posedge ) begin
    lo0142 <= li0142 ;
 end
 always @ (posedge ) begin
    lo0143 <= li0143 ;
 end
 always @ (posedge ) begin
    lo0144 <= li0144 ;
 end
 always @ (posedge ) begin
    lo0145 <= li0145 ;
 end
 always @ (posedge ) begin
    lo0146 <= li0146 ;
 end
 always @ (posedge ) begin
    lo0147 <= li0147 ;
 end
 always @ (posedge ) begin
    lo0148 <= li0148 ;
 end
 always @ (posedge ) begin
    lo0149 <= li0149 ;
 end
 always @ (posedge ) begin
    lo0150 <= li0150 ;
 end
 always @ (posedge ) begin
    lo0151 <= li0151 ;
 end
 always @ (posedge ) begin
    lo0152 <= li0152 ;
 end
 always @ (posedge ) begin
    lo0153 <= li0153 ;
 end
 always @ (posedge ) begin
    lo0154 <= li0154 ;
 end
 always @ (posedge ) begin
    lo0155 <= li0155 ;
 end
 always @ (posedge ) begin
    lo0156 <= li0156 ;
 end
 always @ (posedge ) begin
    lo0157 <= li0157 ;
 end
 always @ (posedge ) begin
    lo0158 <= li0158 ;
 end
 always @ (posedge ) begin
    lo0159 <= li0159 ;
 end
 always @ (posedge ) begin
    lo0160 <= li0160 ;
 end
 always @ (posedge ) begin
    lo0161 <= li0161 ;
 end
 always @ (posedge ) begin
    lo0162 <= li0162 ;
 end
 always @ (posedge ) begin
    lo0163 <= li0163 ;
 end
 always @ (posedge ) begin
    lo0164 <= li0164 ;
 end
 always @ (posedge ) begin
    lo0165 <= li0165 ;
 end
 always @ (posedge ) begin
    lo0166 <= li0166 ;
 end
 always @ (posedge ) begin
    lo0167 <= li0167 ;
 end
 always @ (posedge ) begin
    lo0168 <= li0168 ;
 end
 always @ (posedge ) begin
    lo0169 <= li0169 ;
 end
 always @ (posedge ) begin
    lo0170 <= li0170 ;
 end
 always @ (posedge ) begin
    lo0171 <= li0171 ;
 end
 always @ (posedge ) begin
    lo0172 <= li0172 ;
 end
 always @ (posedge ) begin
    lo0173 <= li0173 ;
 end
 always @ (posedge ) begin
    lo0174 <= li0174 ;
 end
 always @ (posedge ) begin
    lo0175 <= li0175 ;
 end
 always @ (posedge ) begin
    lo0176 <= li0176 ;
 end
 always @ (posedge ) begin
    lo0177 <= li0177 ;
 end
 always @ (posedge ) begin
    lo0178 <= li0178 ;
 end
 always @ (posedge ) begin
    lo0179 <= li0179 ;
 end
 always @ (posedge ) begin
    lo0180 <= li0180 ;
 end
 always @ (posedge ) begin
    lo0181 <= li0181 ;
 end
 always @ (posedge ) begin
    lo0182 <= li0182 ;
 end
 always @ (posedge ) begin
    lo0183 <= li0183 ;
 end
 always @ (posedge ) begin
    lo0184 <= li0184 ;
 end
 always @ (posedge ) begin
    lo0185 <= li0185 ;
 end
 always @ (posedge ) begin
    lo0186 <= li0186 ;
 end
 always @ (posedge ) begin
    lo0187 <= li0187 ;
 end
 always @ (posedge ) begin
    lo0188 <= li0188 ;
 end
 always @ (posedge ) begin
    lo0189 <= li0189 ;
 end
 always @ (posedge ) begin
    lo0190 <= li0190 ;
 end
 always @ (posedge ) begin
    lo0191 <= li0191 ;
 end
 always @ (posedge ) begin
    lo0192 <= li0192 ;
 end
 always @ (posedge ) begin
    lo0193 <= li0193 ;
 end
 always @ (posedge ) begin
    lo0194 <= li0194 ;
 end
 always @ (posedge ) begin
    lo0195 <= li0195 ;
 end
 always @ (posedge ) begin
    lo0196 <= li0196 ;
 end
 always @ (posedge ) begin
    lo0197 <= li0197 ;
 end
 always @ (posedge ) begin
    lo0198 <= li0198 ;
 end
 always @ (posedge ) begin
    lo0199 <= li0199 ;
 end
 always @ (posedge ) begin
    lo0200 <= li0200 ;
 end
 always @ (posedge ) begin
    lo0201 <= li0201 ;
 end
 always @ (posedge ) begin
    lo0202 <= li0202 ;
 end
 always @ (posedge ) begin
    lo0203 <= li0203 ;
 end
 always @ (posedge ) begin
    lo0204 <= li0204 ;
 end
 always @ (posedge ) begin
    lo0205 <= li0205 ;
 end
 always @ (posedge ) begin
    lo0206 <= li0206 ;
 end
 always @ (posedge ) begin
    lo0207 <= li0207 ;
 end
 always @ (posedge ) begin
    lo0208 <= li0208 ;
 end
 always @ (posedge ) begin
    lo0209 <= li0209 ;
 end
 always @ (posedge ) begin
    lo0210 <= li0210 ;
 end
 always @ (posedge ) begin
    lo0211 <= li0211 ;
 end
 always @ (posedge ) begin
    lo0212 <= li0212 ;
 end
 always @ (posedge ) begin
    lo0213 <= li0213 ;
 end
 always @ (posedge ) begin
    lo0214 <= li0214 ;
 end
 always @ (posedge ) begin
    lo0215 <= li0215 ;
 end
 always @ (posedge ) begin
    lo0216 <= li0216 ;
 end
 always @ (posedge ) begin
    lo0217 <= li0217 ;
 end
 always @ (posedge ) begin
    lo0218 <= li0218 ;
 end
 always @ (posedge ) begin
    lo0219 <= li0219 ;
 end
 always @ (posedge ) begin
    lo0220 <= li0220 ;
 end
 always @ (posedge ) begin
    lo0221 <= li0221 ;
 end
 always @ (posedge ) begin
    lo0222 <= li0222 ;
 end
 always @ (posedge ) begin
    lo0223 <= li0223 ;
 end
 always @ (posedge ) begin
    lo0224 <= li0224 ;
 end
 always @ (posedge ) begin
    lo0225 <= li0225 ;
 end
 always @ (posedge ) begin
    lo0226 <= li0226 ;
 end
 always @ (posedge ) begin
    lo0227 <= li0227 ;
 end
 always @ (posedge ) begin
    lo0228 <= li0228 ;
 end
 always @ (posedge ) begin
    lo0229 <= li0229 ;
 end
 always @ (posedge ) begin
    lo0230 <= li0230 ;
 end
 always @ (posedge ) begin
    lo0231 <= li0231 ;
 end
 always @ (posedge ) begin
    lo0232 <= li0232 ;
 end
 always @ (posedge ) begin
    lo0233 <= li0233 ;
 end
 always @ (posedge ) begin
    lo0234 <= li0234 ;
 end
 always @ (posedge ) begin
    lo0235 <= li0235 ;
 end
 always @ (posedge ) begin
    lo0236 <= li0236 ;
 end
 always @ (posedge ) begin
    lo0237 <= li0237 ;
 end
 always @ (posedge ) begin
    lo0238 <= li0238 ;
 end
 always @ (posedge ) begin
    lo0239 <= li0239 ;
 end
 always @ (posedge ) begin
    lo0240 <= li0240 ;
 end
 always @ (posedge ) begin
    lo0241 <= li0241 ;
 end
 always @ (posedge ) begin
    lo0242 <= li0242 ;
 end
 always @ (posedge ) begin
    lo0243 <= li0243 ;
 end
 always @ (posedge ) begin
    lo0244 <= li0244 ;
 end
 always @ (posedge ) begin
    lo0245 <= li0245 ;
 end
 always @ (posedge ) begin
    lo0246 <= li0246 ;
 end
 always @ (posedge ) begin
    lo0247 <= li0247 ;
 end
 always @ (posedge ) begin
    lo0248 <= li0248 ;
 end
 always @ (posedge ) begin
    lo0249 <= li0249 ;
 end
 always @ (posedge ) begin
    lo0250 <= li0250 ;
 end
 always @ (posedge ) begin
    lo0251 <= li0251 ;
 end
 always @ (posedge ) begin
    lo0252 <= li0252 ;
 end
 always @ (posedge ) begin
    lo0253 <= li0253 ;
 end
 always @ (posedge ) begin
    lo0254 <= li0254 ;
 end
 always @ (posedge ) begin
    lo0255 <= li0255 ;
 end
 always @ (posedge ) begin
    lo0256 <= li0256 ;
 end
 always @ (posedge ) begin
    lo0257 <= li0257 ;
 end
 always @ (posedge ) begin
    lo0258 <= li0258 ;
 end
 always @ (posedge ) begin
    lo0259 <= li0259 ;
 end
 always @ (posedge ) begin
    lo0260 <= li0260 ;
 end
 always @ (posedge ) begin
    lo0261 <= li0261 ;
 end
 always @ (posedge ) begin
    lo0262 <= li0262 ;
 end
 always @ (posedge ) begin
    lo0263 <= li0263 ;
 end
 always @ (posedge ) begin
    lo0264 <= li0264 ;
 end
 always @ (posedge ) begin
    lo0265 <= li0265 ;
 end
 always @ (posedge ) begin
    lo0266 <= li0266 ;
 end
 always @ (posedge ) begin
    lo0267 <= li0267 ;
 end
 always @ (posedge ) begin
    lo0268 <= li0268 ;
 end
 always @ (posedge ) begin
    lo0269 <= li0269 ;
 end
 always @ (posedge ) begin
    lo0270 <= li0270 ;
 end
 always @ (posedge ) begin
    lo0271 <= li0271 ;
 end
 always @ (posedge ) begin
    lo0272 <= li0272 ;
 end
 always @ (posedge ) begin
    lo0273 <= li0273 ;
 end
 always @ (posedge ) begin
    lo0274 <= li0274 ;
 end
 always @ (posedge ) begin
    lo0275 <= li0275 ;
 end
 always @ (posedge ) begin
    lo0276 <= li0276 ;
 end
 always @ (posedge ) begin
    lo0277 <= li0277 ;
 end
 always @ (posedge ) begin
    lo0278 <= li0278 ;
 end
 always @ (posedge ) begin
    lo0279 <= li0279 ;
 end
 always @ (posedge ) begin
    lo0280 <= li0280 ;
 end
 always @ (posedge ) begin
    lo0281 <= li0281 ;
 end
 always @ (posedge ) begin
    lo0282 <= li0282 ;
 end
 always @ (posedge ) begin
    lo0283 <= li0283 ;
 end
 always @ (posedge ) begin
    lo0284 <= li0284 ;
 end
 always @ (posedge ) begin
    lo0285 <= li0285 ;
 end
 always @ (posedge ) begin
    lo0286 <= li0286 ;
 end
 always @ (posedge ) begin
    lo0287 <= li0287 ;
 end
 always @ (posedge ) begin
    lo0288 <= li0288 ;
 end
 always @ (posedge ) begin
    lo0289 <= li0289 ;
 end
 always @ (posedge ) begin
    lo0290 <= li0290 ;
 end
 always @ (posedge ) begin
    lo0291 <= li0291 ;
 end
 always @ (posedge ) begin
    lo0292 <= li0292 ;
 end
 always @ (posedge ) begin
    lo0293 <= li0293 ;
 end
 always @ (posedge ) begin
    lo0294 <= li0294 ;
 end
 always @ (posedge ) begin
    lo0295 <= li0295 ;
 end
 always @ (posedge ) begin
    lo0296 <= li0296 ;
 end
 always @ (posedge ) begin
    lo0297 <= li0297 ;
 end
 always @ (posedge ) begin
    lo0298 <= li0298 ;
 end
 always @ (posedge ) begin
    lo0299 <= li0299 ;
 end
 always @ (posedge ) begin
    lo0300 <= li0300 ;
 end
 always @ (posedge ) begin
    lo0301 <= li0301 ;
 end
 always @ (posedge ) begin
    lo0302 <= li0302 ;
 end
 always @ (posedge ) begin
    lo0303 <= li0303 ;
 end
 always @ (posedge ) begin
    lo0304 <= li0304 ;
 end
 always @ (posedge ) begin
    lo0305 <= li0305 ;
 end
 always @ (posedge ) begin
    lo0306 <= li0306 ;
 end
 always @ (posedge ) begin
    lo0307 <= li0307 ;
 end
 always @ (posedge ) begin
    lo0308 <= li0308 ;
 end
 always @ (posedge ) begin
    lo0309 <= li0309 ;
 end
 always @ (posedge ) begin
    lo0310 <= li0310 ;
 end
 always @ (posedge ) begin
    lo0311 <= li0311 ;
 end
 always @ (posedge ) begin
    lo0312 <= li0312 ;
 end
 always @ (posedge ) begin
    lo0313 <= li0313 ;
 end
 always @ (posedge ) begin
    lo0314 <= li0314 ;
 end
 always @ (posedge ) begin
    lo0315 <= li0315 ;
 end
 always @ (posedge ) begin
    lo0316 <= li0316 ;
 end
 always @ (posedge ) begin
    lo0317 <= li0317 ;
 end
 always @ (posedge ) begin
    lo0318 <= li0318 ;
 end
 always @ (posedge ) begin
    lo0319 <= li0319 ;
 end
 always @ (posedge ) begin
    lo0320 <= li0320 ;
 end
 always @ (posedge ) begin
    lo0321 <= li0321 ;
 end
 always @ (posedge ) begin
    lo0322 <= li0322 ;
 end
 always @ (posedge ) begin
    lo0323 <= li0323 ;
 end
 always @ (posedge ) begin
    lo0324 <= li0324 ;
 end
 always @ (posedge ) begin
    lo0325 <= li0325 ;
 end
 always @ (posedge ) begin
    lo0326 <= li0326 ;
 end
 always @ (posedge ) begin
    lo0327 <= li0327 ;
 end
 always @ (posedge ) begin
    lo0328 <= li0328 ;
 end
 always @ (posedge ) begin
    lo0329 <= li0329 ;
 end
 always @ (posedge ) begin
    lo0330 <= li0330 ;
 end
 always @ (posedge ) begin
    lo0331 <= li0331 ;
 end
 always @ (posedge ) begin
    lo0332 <= li0332 ;
 end
 always @ (posedge ) begin
    lo0333 <= li0333 ;
 end
 always @ (posedge ) begin
    lo0334 <= li0334 ;
 end
 always @ (posedge ) begin
    lo0335 <= li0335 ;
 end
 always @ (posedge ) begin
    lo0336 <= li0336 ;
 end
 always @ (posedge ) begin
    lo0337 <= li0337 ;
 end
 always @ (posedge ) begin
    lo0338 <= li0338 ;
 end
 always @ (posedge ) begin
    lo0339 <= li0339 ;
 end
 always @ (posedge ) begin
    lo0340 <= li0340 ;
 end
 always @ (posedge ) begin
    lo0341 <= li0341 ;
 end
 always @ (posedge ) begin
    lo0342 <= li0342 ;
 end
 always @ (posedge ) begin
    lo0343 <= li0343 ;
 end
 always @ (posedge ) begin
    lo0344 <= li0344 ;
 end
 always @ (posedge ) begin
    lo0345 <= li0345 ;
 end
 always @ (posedge ) begin
    lo0346 <= li0346 ;
 end
 always @ (posedge ) begin
    lo0347 <= li0347 ;
 end
 always @ (posedge ) begin
    lo0348 <= li0348 ;
 end
 always @ (posedge ) begin
    lo0349 <= li0349 ;
 end
 always @ (posedge ) begin
    lo0350 <= li0350 ;
 end
 always @ (posedge ) begin
    lo0351 <= li0351 ;
 end
 always @ (posedge ) begin
    lo0352 <= li0352 ;
 end
 always @ (posedge ) begin
    lo0353 <= li0353 ;
 end
 always @ (posedge ) begin
    lo0354 <= li0354 ;
 end
 always @ (posedge ) begin
    lo0355 <= li0355 ;
 end
 always @ (posedge ) begin
    lo0356 <= li0356 ;
 end
 always @ (posedge ) begin
    lo0357 <= li0357 ;
 end
 always @ (posedge ) begin
    lo0358 <= li0358 ;
 end
 always @ (posedge ) begin
    lo0359 <= li0359 ;
 end
 always @ (posedge ) begin
    lo0360 <= li0360 ;
 end
 always @ (posedge ) begin
    lo0361 <= li0361 ;
 end
 always @ (posedge ) begin
    lo0362 <= li0362 ;
 end
 always @ (posedge ) begin
    lo0363 <= li0363 ;
 end
 always @ (posedge ) begin
    lo0364 <= li0364 ;
 end
 always @ (posedge ) begin
    lo0365 <= li0365 ;
 end
 always @ (posedge ) begin
    lo0366 <= li0366 ;
 end
 always @ (posedge ) begin
    lo0367 <= li0367 ;
 end
 always @ (posedge ) begin
    lo0368 <= li0368 ;
 end
 always @ (posedge ) begin
    lo0369 <= li0369 ;
 end
 always @ (posedge ) begin
    lo0370 <= li0370 ;
 end
 always @ (posedge ) begin
    lo0371 <= li0371 ;
 end
 always @ (posedge ) begin
    lo0372 <= li0372 ;
 end
 always @ (posedge ) begin
    lo0373 <= li0373 ;
 end
 always @ (posedge ) begin
    lo0374 <= li0374 ;
 end
 always @ (posedge ) begin
    lo0375 <= li0375 ;
 end
 always @ (posedge ) begin
    lo0376 <= li0376 ;
 end
 always @ (posedge ) begin
    lo0377 <= li0377 ;
 end
 always @ (posedge ) begin
    lo0378 <= li0378 ;
 end
 always @ (posedge ) begin
    lo0379 <= li0379 ;
 end
 always @ (posedge ) begin
    lo0380 <= li0380 ;
 end
 always @ (posedge ) begin
    lo0381 <= li0381 ;
 end
 always @ (posedge ) begin
    lo0382 <= li0382 ;
 end
 always @ (posedge ) begin
    lo0383 <= li0383 ;
 end
 always @ (posedge ) begin
    lo0384 <= li0384 ;
 end
 always @ (posedge ) begin
    lo0385 <= li0385 ;
 end
 always @ (posedge ) begin
    lo0386 <= li0386 ;
 end
 always @ (posedge ) begin
    lo0387 <= li0387 ;
 end
 always @ (posedge ) begin
    lo0388 <= li0388 ;
 end
 always @ (posedge ) begin
    lo0389 <= li0389 ;
 end
 always @ (posedge ) begin
    lo0390 <= li0390 ;
 end
 always @ (posedge ) begin
    lo0391 <= li0391 ;
 end
 always @ (posedge ) begin
    lo0392 <= li0392 ;
 end
 always @ (posedge ) begin
    lo0393 <= li0393 ;
 end
 always @ (posedge ) begin
    lo0394 <= li0394 ;
 end
 always @ (posedge ) begin
    lo0395 <= li0395 ;
 end
 always @ (posedge ) begin
    lo0396 <= li0396 ;
 end
 always @ (posedge ) begin
    lo0397 <= li0397 ;
 end
 always @ (posedge ) begin
    lo0398 <= li0398 ;
 end
 always @ (posedge ) begin
    lo0399 <= li0399 ;
 end
 always @ (posedge ) begin
    lo0400 <= li0400 ;
 end
 always @ (posedge ) begin
    lo0401 <= li0401 ;
 end
 always @ (posedge ) begin
    lo0402 <= li0402 ;
 end
 always @ (posedge ) begin
    lo0403 <= li0403 ;
 end
 always @ (posedge ) begin
    lo0404 <= li0404 ;
 end
 always @ (posedge ) begin
    lo0405 <= li0405 ;
 end
 always @ (posedge ) begin
    lo0406 <= li0406 ;
 end
 always @ (posedge ) begin
    lo0407 <= li0407 ;
 end
 always @ (posedge ) begin
    lo0408 <= li0408 ;
 end
 always @ (posedge ) begin
    lo0409 <= li0409 ;
 end
 always @ (posedge ) begin
    lo0410 <= li0410 ;
 end
 always @ (posedge ) begin
    lo0411 <= li0411 ;
 end
 always @ (posedge ) begin
    lo0412 <= li0412 ;
 end
 always @ (posedge ) begin
    lo0413 <= li0413 ;
 end
 always @ (posedge ) begin
    lo0414 <= li0414 ;
 end
 always @ (posedge ) begin
    lo0415 <= li0415 ;
 end
 always @ (posedge ) begin
    lo0416 <= li0416 ;
 end
 always @ (posedge ) begin
    lo0417 <= li0417 ;
 end
 always @ (posedge ) begin
    lo0418 <= li0418 ;
 end
 always @ (posedge ) begin
    lo0419 <= li0419 ;
 end
 always @ (posedge ) begin
    lo0420 <= li0420 ;
 end
 always @ (posedge ) begin
    lo0421 <= li0421 ;
 end
 always @ (posedge ) begin
    lo0422 <= li0422 ;
 end
 always @ (posedge ) begin
    lo0423 <= li0423 ;
 end
 always @ (posedge ) begin
    lo0424 <= li0424 ;
 end
 always @ (posedge ) begin
    lo0425 <= li0425 ;
 end
 always @ (posedge ) begin
    lo0426 <= li0426 ;
 end
 always @ (posedge ) begin
    lo0427 <= li0427 ;
 end
 always @ (posedge ) begin
    lo0428 <= li0428 ;
 end
 always @ (posedge ) begin
    lo0429 <= li0429 ;
 end
 always @ (posedge ) begin
    lo0430 <= li0430 ;
 end
 always @ (posedge ) begin
    lo0431 <= li0431 ;
 end
 always @ (posedge ) begin
    lo0432 <= li0432 ;
 end
 always @ (posedge ) begin
    lo0433 <= li0433 ;
 end
 always @ (posedge ) begin
    lo0434 <= li0434 ;
 end
 always @ (posedge ) begin
    lo0435 <= li0435 ;
 end
 always @ (posedge ) begin
    lo0436 <= li0436 ;
 end
 always @ (posedge ) begin
    lo0437 <= li0437 ;
 end
 always @ (posedge ) begin
    lo0438 <= li0438 ;
 end
 always @ (posedge ) begin
    lo0439 <= li0439 ;
 end
 always @ (posedge ) begin
    lo0440 <= li0440 ;
 end
 always @ (posedge ) begin
    lo0441 <= li0441 ;
 end
 always @ (posedge ) begin
    lo0442 <= li0442 ;
 end
 always @ (posedge ) begin
    lo0443 <= li0443 ;
 end
 always @ (posedge ) begin
    lo0444 <= li0444 ;
 end
 always @ (posedge ) begin
    lo0445 <= li0445 ;
 end
 always @ (posedge ) begin
    lo0446 <= li0446 ;
 end
 always @ (posedge ) begin
    lo0447 <= li0447 ;
 end
 always @ (posedge ) begin
    lo0448 <= li0448 ;
 end
 always @ (posedge ) begin
    lo0449 <= li0449 ;
 end
 always @ (posedge ) begin
    lo0450 <= li0450 ;
 end
 always @ (posedge ) begin
    lo0451 <= li0451 ;
 end
 always @ (posedge ) begin
    lo0452 <= li0452 ;
 end
 always @ (posedge ) begin
    lo0453 <= li0453 ;
 end
 always @ (posedge ) begin
    lo0454 <= li0454 ;
 end
 always @ (posedge ) begin
    lo0455 <= li0455 ;
 end
 always @ (posedge ) begin
    lo0456 <= li0456 ;
 end
 always @ (posedge ) begin
    lo0457 <= li0457 ;
 end
 always @ (posedge ) begin
    lo0458 <= li0458 ;
 end
 always @ (posedge ) begin
    lo0459 <= li0459 ;
 end
 always @ (posedge ) begin
    lo0460 <= li0460 ;
 end
 always @ (posedge ) begin
    lo0461 <= li0461 ;
 end
 always @ (posedge ) begin
    lo0462 <= li0462 ;
 end
 always @ (posedge ) begin
    lo0463 <= li0463 ;
 end
 always @ (posedge ) begin
    lo0464 <= li0464 ;
 end
 always @ (posedge ) begin
    lo0465 <= li0465 ;
 end
 always @ (posedge ) begin
    lo0466 <= li0466 ;
 end
 always @ (posedge ) begin
    lo0467 <= li0467 ;
 end
 always @ (posedge ) begin
    lo0468 <= li0468 ;
 end
 always @ (posedge ) begin
    lo0469 <= li0469 ;
 end
 always @ (posedge ) begin
    lo0470 <= li0470 ;
 end
 always @ (posedge ) begin
    lo0471 <= li0471 ;
 end
 always @ (posedge ) begin
    lo0472 <= li0472 ;
 end
 always @ (posedge ) begin
    lo0473 <= li0473 ;
 end
 always @ (posedge ) begin
    lo0474 <= li0474 ;
 end
 always @ (posedge ) begin
    lo0475 <= li0475 ;
 end
 always @ (posedge ) begin
    lo0476 <= li0476 ;
 end
 always @ (posedge ) begin
    lo0477 <= li0477 ;
 end
 always @ (posedge ) begin
    lo0478 <= li0478 ;
 end
 always @ (posedge ) begin
    lo0479 <= li0479 ;
 end
 always @ (posedge ) begin
    lo0480 <= li0480 ;
 end
 always @ (posedge ) begin
    lo0481 <= li0481 ;
 end
 always @ (posedge ) begin
    lo0482 <= li0482 ;
 end
 always @ (posedge ) begin
    lo0483 <= li0483 ;
 end
 always @ (posedge ) begin
    lo0484 <= li0484 ;
 end
 always @ (posedge ) begin
    lo0485 <= li0485 ;
 end
 always @ (posedge ) begin
    lo0486 <= li0486 ;
 end
 always @ (posedge ) begin
    lo0487 <= li0487 ;
 end
 always @ (posedge ) begin
    lo0488 <= li0488 ;
 end
 always @ (posedge ) begin
    lo0489 <= li0489 ;
 end
 always @ (posedge ) begin
    lo0490 <= li0490 ;
 end
 always @ (posedge ) begin
    lo0491 <= li0491 ;
 end
 always @ (posedge ) begin
    lo0492 <= li0492 ;
 end
 always @ (posedge ) begin
    lo0493 <= li0493 ;
 end
 always @ (posedge ) begin
    lo0494 <= li0494 ;
 end
 always @ (posedge ) begin
    lo0495 <= li0495 ;
 end
 always @ (posedge ) begin
    lo0496 <= li0496 ;
 end
 always @ (posedge ) begin
    lo0497 <= li0497 ;
 end
 always @ (posedge ) begin
    lo0498 <= li0498 ;
 end
 always @ (posedge ) begin
    lo0499 <= li0499 ;
 end
 always @ (posedge ) begin
    lo0500 <= li0500 ;
 end
 always @ (posedge ) begin
    lo0501 <= li0501 ;
 end
 always @ (posedge ) begin
    lo0502 <= li0502 ;
 end
 always @ (posedge ) begin
    lo0503 <= li0503 ;
 end
 always @ (posedge ) begin
    lo0504 <= li0504 ;
 end
 always @ (posedge ) begin
    lo0505 <= li0505 ;
 end
 always @ (posedge ) begin
    lo0506 <= li0506 ;
 end
 always @ (posedge ) begin
    lo0507 <= li0507 ;
 end
 always @ (posedge ) begin
    lo0508 <= li0508 ;
 end
 always @ (posedge ) begin
    lo0509 <= li0509 ;
 end
 always @ (posedge ) begin
    lo0510 <= li0510 ;
 end
 always @ (posedge ) begin
    lo0511 <= li0511 ;
 end
 always @ (posedge ) begin
    lo0512 <= li0512 ;
 end
 always @ (posedge ) begin
    lo0513 <= li0513 ;
 end
 always @ (posedge ) begin
    lo0514 <= li0514 ;
 end
 always @ (posedge ) begin
    lo0515 <= li0515 ;
 end
 always @ (posedge ) begin
    lo0516 <= li0516 ;
 end
 always @ (posedge ) begin
    lo0517 <= li0517 ;
 end
 always @ (posedge ) begin
    lo0518 <= li0518 ;
 end
 always @ (posedge ) begin
    lo0519 <= li0519 ;
 end
 always @ (posedge ) begin
    lo0520 <= li0520 ;
 end
 always @ (posedge ) begin
    lo0521 <= li0521 ;
 end
 always @ (posedge ) begin
    lo0522 <= li0522 ;
 end
 always @ (posedge ) begin
    lo0523 <= li0523 ;
 end
 always @ (posedge ) begin
    lo0524 <= li0524 ;
 end
 always @ (posedge ) begin
    lo0525 <= li0525 ;
 end
 always @ (posedge ) begin
    lo0526 <= li0526 ;
 end
 always @ (posedge ) begin
    lo0527 <= li0527 ;
 end
 always @ (posedge ) begin
    lo0528 <= li0528 ;
 end
 always @ (posedge ) begin
    lo0529 <= li0529 ;
 end
 always @ (posedge ) begin
    lo0530 <= li0530 ;
 end
 always @ (posedge ) begin
    lo0531 <= li0531 ;
 end
 always @ (posedge ) begin
    lo0532 <= li0532 ;
 end
 always @ (posedge ) begin
    lo0533 <= li0533 ;
 end
 always @ (posedge ) begin
    lo0534 <= li0534 ;
 end
 always @ (posedge ) begin
    lo0535 <= li0535 ;
 end
 always @ (posedge ) begin
    lo0536 <= li0536 ;
 end
 always @ (posedge ) begin
    lo0537 <= li0537 ;
 end
 always @ (posedge ) begin
    lo0538 <= li0538 ;
 end
 always @ (posedge ) begin
    lo0539 <= li0539 ;
 end
 always @ (posedge ) begin
    lo0540 <= li0540 ;
 end
 always @ (posedge ) begin
    lo0541 <= li0541 ;
 end
 always @ (posedge ) begin
    lo0542 <= li0542 ;
 end
 always @ (posedge ) begin
    lo0543 <= li0543 ;
 end
 always @ (posedge ) begin
    lo0544 <= li0544 ;
 end
 always @ (posedge ) begin
    lo0545 <= li0545 ;
 end
 always @ (posedge ) begin
    lo0546 <= li0546 ;
 end
 always @ (posedge ) begin
    lo0547 <= li0547 ;
 end
 always @ (posedge ) begin
    lo0548 <= li0548 ;
 end
 always @ (posedge ) begin
    lo0549 <= li0549 ;
 end
 always @ (posedge ) begin
    lo0550 <= li0550 ;
 end
 always @ (posedge ) begin
    lo0551 <= li0551 ;
 end
 always @ (posedge ) begin
    lo0552 <= li0552 ;
 end
 always @ (posedge ) begin
    lo0553 <= li0553 ;
 end
 always @ (posedge ) begin
    lo0554 <= li0554 ;
 end
 always @ (posedge ) begin
    lo0555 <= li0555 ;
 end
 always @ (posedge ) begin
    lo0556 <= li0556 ;
 end
 always @ (posedge ) begin
    lo0557 <= li0557 ;
 end
 always @ (posedge ) begin
    lo0558 <= li0558 ;
 end
 always @ (posedge ) begin
    lo0559 <= li0559 ;
 end
 always @ (posedge ) begin
    lo0560 <= li0560 ;
 end
 always @ (posedge ) begin
    lo0561 <= li0561 ;
 end
 always @ (posedge ) begin
    lo0562 <= li0562 ;
 end
 always @ (posedge ) begin
    lo0563 <= li0563 ;
 end
 always @ (posedge ) begin
    lo0564 <= li0564 ;
 end
 always @ (posedge ) begin
    lo0565 <= li0565 ;
 end
 always @ (posedge ) begin
    lo0566 <= li0566 ;
 end
 always @ (posedge ) begin
    lo0567 <= li0567 ;
 end
 always @ (posedge ) begin
    lo0568 <= li0568 ;
 end
 always @ (posedge ) begin
    lo0569 <= li0569 ;
 end
 always @ (posedge ) begin
    lo0570 <= li0570 ;
 end
 always @ (posedge ) begin
    lo0571 <= li0571 ;
 end
 always @ (posedge ) begin
    lo0572 <= li0572 ;
 end
 always @ (posedge ) begin
    lo0573 <= li0573 ;
 end
 always @ (posedge ) begin
    lo0574 <= li0574 ;
 end
 always @ (posedge ) begin
    lo0575 <= li0575 ;
 end
 always @ (posedge ) begin
    lo0576 <= li0576 ;
 end
 always @ (posedge ) begin
    lo0577 <= li0577 ;
 end
 always @ (posedge ) begin
    lo0578 <= li0578 ;
 end
 always @ (posedge ) begin
    lo0579 <= li0579 ;
 end
 always @ (posedge ) begin
    lo0580 <= li0580 ;
 end
 always @ (posedge ) begin
    lo0581 <= li0581 ;
 end
 always @ (posedge ) begin
    lo0582 <= li0582 ;
 end
 always @ (posedge ) begin
    lo0583 <= li0583 ;
 end
 always @ (posedge ) begin
    lo0584 <= li0584 ;
 end
 always @ (posedge ) begin
    lo0585 <= li0585 ;
 end
 always @ (posedge ) begin
    lo0586 <= li0586 ;
 end
 always @ (posedge ) begin
    lo0587 <= li0587 ;
 end
 always @ (posedge ) begin
    lo0588 <= li0588 ;
 end
 always @ (posedge ) begin
    lo0589 <= li0589 ;
 end
 always @ (posedge ) begin
    lo0590 <= li0590 ;
 end
 always @ (posedge ) begin
    lo0591 <= li0591 ;
 end
 always @ (posedge ) begin
    lo0592 <= li0592 ;
 end
 always @ (posedge ) begin
    lo0593 <= li0593 ;
 end
 always @ (posedge ) begin
    lo0594 <= li0594 ;
 end
 always @ (posedge ) begin
    lo0595 <= li0595 ;
 end
 always @ (posedge ) begin
    lo0596 <= li0596 ;
 end
 always @ (posedge ) begin
    lo0597 <= li0597 ;
 end
 always @ (posedge ) begin
    lo0598 <= li0598 ;
 end
 always @ (posedge ) begin
    lo0599 <= li0599 ;
 end
 always @ (posedge ) begin
    lo0600 <= li0600 ;
 end
 always @ (posedge ) begin
    lo0601 <= li0601 ;
 end
 always @ (posedge ) begin
    lo0602 <= li0602 ;
 end
 always @ (posedge ) begin
    lo0603 <= li0603 ;
 end
 always @ (posedge ) begin
    lo0604 <= li0604 ;
 end
 always @ (posedge ) begin
    lo0605 <= li0605 ;
 end
 always @ (posedge ) begin
    lo0606 <= li0606 ;
 end
 always @ (posedge ) begin
    lo0607 <= li0607 ;
 end
 always @ (posedge ) begin
    lo0608 <= li0608 ;
 end
 always @ (posedge ) begin
    lo0609 <= li0609 ;
 end
 always @ (posedge ) begin
    lo0610 <= li0610 ;
 end
 always @ (posedge ) begin
    lo0611 <= li0611 ;
 end
 always @ (posedge ) begin
    lo0612 <= li0612 ;
 end
 always @ (posedge ) begin
    lo0613 <= li0613 ;
 end
 always @ (posedge ) begin
    lo0614 <= li0614 ;
 end
 always @ (posedge ) begin
    lo0615 <= li0615 ;
 end
 always @ (posedge ) begin
    lo0616 <= li0616 ;
 end
 always @ (posedge ) begin
    lo0617 <= li0617 ;
 end
 always @ (posedge ) begin
    lo0618 <= li0618 ;
 end
 always @ (posedge ) begin
    lo0619 <= li0619 ;
 end
 always @ (posedge ) begin
    lo0620 <= li0620 ;
 end
 always @ (posedge ) begin
    lo0621 <= li0621 ;
 end
 always @ (posedge ) begin
    lo0622 <= li0622 ;
 end
 always @ (posedge ) begin
    lo0623 <= li0623 ;
 end
 always @ (posedge ) begin
    lo0624 <= li0624 ;
 end
 always @ (posedge ) begin
    lo0625 <= li0625 ;
 end
 always @ (posedge ) begin
    lo0626 <= li0626 ;
 end
 always @ (posedge ) begin
    lo0627 <= li0627 ;
 end
 always @ (posedge ) begin
    lo0628 <= li0628 ;
 end
 always @ (posedge ) begin
    lo0629 <= li0629 ;
 end
 always @ (posedge ) begin
    lo0630 <= li0630 ;
 end
 always @ (posedge ) begin
    lo0631 <= li0631 ;
 end
 always @ (posedge ) begin
    lo0632 <= li0632 ;
 end
 always @ (posedge ) begin
    lo0633 <= li0633 ;
 end
 always @ (posedge ) begin
    lo0634 <= li0634 ;
 end
 always @ (posedge ) begin
    lo0635 <= li0635 ;
 end
 always @ (posedge ) begin
    lo0636 <= li0636 ;
 end
 always @ (posedge ) begin
    lo0637 <= li0637 ;
 end
 always @ (posedge ) begin
    lo0638 <= li0638 ;
 end
 always @ (posedge ) begin
    lo0639 <= li0639 ;
 end
 always @ (posedge ) begin
    lo0640 <= li0640 ;
 end
 always @ (posedge ) begin
    lo0641 <= li0641 ;
 end
 always @ (posedge ) begin
    lo0642 <= li0642 ;
 end
 always @ (posedge ) begin
    lo0643 <= li0643 ;
 end
 always @ (posedge ) begin
    lo0644 <= li0644 ;
 end
 always @ (posedge ) begin
    lo0645 <= li0645 ;
 end
 always @ (posedge ) begin
    lo0646 <= li0646 ;
 end
 always @ (posedge ) begin
    lo0647 <= li0647 ;
 end
 always @ (posedge ) begin
    lo0648 <= li0648 ;
 end
 always @ (posedge ) begin
    lo0649 <= li0649 ;
 end
 always @ (posedge ) begin
    lo0650 <= li0650 ;
 end
 always @ (posedge ) begin
    lo0651 <= li0651 ;
 end
 always @ (posedge ) begin
    lo0652 <= li0652 ;
 end
 always @ (posedge ) begin
    lo0653 <= li0653 ;
 end
 always @ (posedge ) begin
    lo0654 <= li0654 ;
 end
 always @ (posedge ) begin
    lo0655 <= li0655 ;
 end
 always @ (posedge ) begin
    lo0656 <= li0656 ;
 end
 always @ (posedge ) begin
    lo0657 <= li0657 ;
 end
 always @ (posedge ) begin
    lo0658 <= li0658 ;
 end
 always @ (posedge ) begin
    lo0659 <= li0659 ;
 end
 always @ (posedge ) begin
    lo0660 <= li0660 ;
 end
 always @ (posedge ) begin
    lo0661 <= li0661 ;
 end
 always @ (posedge ) begin
    lo0662 <= li0662 ;
 end
 always @ (posedge ) begin
    lo0663 <= li0663 ;
 end
 always @ (posedge ) begin
    lo0664 <= li0664 ;
 end
 always @ (posedge ) begin
    lo0665 <= li0665 ;
 end
 always @ (posedge ) begin
    lo0666 <= li0666 ;
 end
 always @ (posedge ) begin
    lo0667 <= li0667 ;
 end
 always @ (posedge ) begin
    lo0668 <= li0668 ;
 end
 always @ (posedge ) begin
    lo0669 <= li0669 ;
 end
 always @ (posedge ) begin
    lo0670 <= li0670 ;
 end
 always @ (posedge ) begin
    lo0671 <= li0671 ;
 end
 always @ (posedge ) begin
    lo0672 <= li0672 ;
 end
 always @ (posedge ) begin
    lo0673 <= li0673 ;
 end
 always @ (posedge ) begin
    lo0674 <= li0674 ;
 end
 always @ (posedge ) begin
    lo0675 <= li0675 ;
 end
 always @ (posedge ) begin
    lo0676 <= li0676 ;
 end
 always @ (posedge ) begin
    lo0677 <= li0677 ;
 end
 always @ (posedge ) begin
    lo0678 <= li0678 ;
 end
 always @ (posedge ) begin
    lo0679 <= li0679 ;
 end
 always @ (posedge ) begin
    lo0680 <= li0680 ;
 end
 always @ (posedge ) begin
    lo0681 <= li0681 ;
 end
 always @ (posedge ) begin
    lo0682 <= li0682 ;
 end
 always @ (posedge ) begin
    lo0683 <= li0683 ;
 end
 always @ (posedge ) begin
    lo0684 <= li0684 ;
 end
 always @ (posedge ) begin
    lo0685 <= li0685 ;
 end
 always @ (posedge ) begin
    lo0686 <= li0686 ;
 end
 always @ (posedge ) begin
    lo0687 <= li0687 ;
 end
 always @ (posedge ) begin
    lo0688 <= li0688 ;
 end
 always @ (posedge ) begin
    lo0689 <= li0689 ;
 end
 always @ (posedge ) begin
    lo0690 <= li0690 ;
 end
 always @ (posedge ) begin
    lo0691 <= li0691 ;
 end
 always @ (posedge ) begin
    lo0692 <= li0692 ;
 end
 always @ (posedge ) begin
    lo0693 <= li0693 ;
 end
 always @ (posedge ) begin
    lo0694 <= li0694 ;
 end
 always @ (posedge ) begin
    lo0695 <= li0695 ;
 end
 always @ (posedge ) begin
    lo0696 <= li0696 ;
 end
 always @ (posedge ) begin
    lo0697 <= li0697 ;
 end
 always @ (posedge ) begin
    lo0698 <= li0698 ;
 end
 always @ (posedge ) begin
    lo0699 <= li0699 ;
 end
 always @ (posedge ) begin
    lo0700 <= li0700 ;
 end
 always @ (posedge ) begin
    lo0701 <= li0701 ;
 end
 always @ (posedge ) begin
    lo0702 <= li0702 ;
 end
 always @ (posedge ) begin
    lo0703 <= li0703 ;
 end
 always @ (posedge ) begin
    lo0704 <= li0704 ;
 end
 always @ (posedge ) begin
    lo0705 <= li0705 ;
 end
 always @ (posedge ) begin
    lo0706 <= li0706 ;
 end
 always @ (posedge ) begin
    lo0707 <= li0707 ;
 end
 always @ (posedge ) begin
    lo0708 <= li0708 ;
 end
 always @ (posedge ) begin
    lo0709 <= li0709 ;
 end
 always @ (posedge ) begin
    lo0710 <= li0710 ;
 end
 always @ (posedge ) begin
    lo0711 <= li0711 ;
 end
 always @ (posedge ) begin
    lo0712 <= li0712 ;
 end
 always @ (posedge ) begin
    lo0713 <= li0713 ;
 end
 always @ (posedge ) begin
    lo0714 <= li0714 ;
 end
 always @ (posedge ) begin
    lo0715 <= li0715 ;
 end
 always @ (posedge ) begin
    lo0716 <= li0716 ;
 end
 always @ (posedge ) begin
    lo0717 <= li0717 ;
 end
 always @ (posedge ) begin
    lo0718 <= li0718 ;
 end
 always @ (posedge ) begin
    lo0719 <= li0719 ;
 end
 always @ (posedge ) begin
    lo0720 <= li0720 ;
 end
 always @ (posedge ) begin
    lo0721 <= li0721 ;
 end
 always @ (posedge ) begin
    lo0722 <= li0722 ;
 end
 always @ (posedge ) begin
    lo0723 <= li0723 ;
 end
 always @ (posedge ) begin
    lo0724 <= li0724 ;
 end
 always @ (posedge ) begin
    lo0725 <= li0725 ;
 end
 always @ (posedge ) begin
    lo0726 <= li0726 ;
 end
 always @ (posedge ) begin
    lo0727 <= li0727 ;
 end
 always @ (posedge ) begin
    lo0728 <= li0728 ;
 end
 always @ (posedge ) begin
    lo0729 <= li0729 ;
 end
 always @ (posedge ) begin
    lo0730 <= li0730 ;
 end
 always @ (posedge ) begin
    lo0731 <= li0731 ;
 end
 always @ (posedge ) begin
    lo0732 <= li0732 ;
 end
 always @ (posedge ) begin
    lo0733 <= li0733 ;
 end
 always @ (posedge ) begin
    lo0734 <= li0734 ;
 end
 always @ (posedge ) begin
    lo0735 <= li0735 ;
 end
 always @ (posedge ) begin
    lo0736 <= li0736 ;
 end
 always @ (posedge ) begin
    lo0737 <= li0737 ;
 end
 always @ (posedge ) begin
    lo0738 <= li0738 ;
 end
 always @ (posedge ) begin
    lo0739 <= li0739 ;
 end
 always @ (posedge ) begin
    lo0740 <= li0740 ;
 end
 always @ (posedge ) begin
    lo0741 <= li0741 ;
 end
 always @ (posedge ) begin
    lo0742 <= li0742 ;
 end
 always @ (posedge ) begin
    lo0743 <= li0743 ;
 end
 always @ (posedge ) begin
    lo0744 <= li0744 ;
 end
 always @ (posedge ) begin
    lo0745 <= li0745 ;
 end
 always @ (posedge ) begin
    lo0746 <= li0746 ;
 end
 always @ (posedge ) begin
    lo0747 <= li0747 ;
 end
 always @ (posedge ) begin
    lo0748 <= li0748 ;
 end
 always @ (posedge ) begin
    lo0749 <= li0749 ;
 end
 always @ (posedge ) begin
    lo0750 <= li0750 ;
 end
 always @ (posedge ) begin
    lo0751 <= li0751 ;
 end
 always @ (posedge ) begin
    lo0752 <= li0752 ;
 end
 always @ (posedge ) begin
    lo0753 <= li0753 ;
 end
 always @ (posedge ) begin
    lo0754 <= li0754 ;
 end
 always @ (posedge ) begin
    lo0755 <= li0755 ;
 end
 always @ (posedge ) begin
    lo0756 <= li0756 ;
 end
 always @ (posedge ) begin
    lo0757 <= li0757 ;
 end
 always @ (posedge ) begin
    lo0758 <= li0758 ;
 end
 always @ (posedge ) begin
    lo0759 <= li0759 ;
 end
 always @ (posedge ) begin
    lo0760 <= li0760 ;
 end
 always @ (posedge ) begin
    lo0761 <= li0761 ;
 end
 always @ (posedge ) begin
    lo0762 <= li0762 ;
 end
 always @ (posedge ) begin
    lo0763 <= li0763 ;
 end
 always @ (posedge ) begin
    lo0764 <= li0764 ;
 end
 always @ (posedge ) begin
    lo0765 <= li0765 ;
 end
 always @ (posedge ) begin
    lo0766 <= li0766 ;
 end
 always @ (posedge ) begin
    lo0767 <= li0767 ;
 end
 always @ (posedge ) begin
    lo0768 <= li0768 ;
 end
 always @ (posedge ) begin
    lo0769 <= li0769 ;
 end
 always @ (posedge ) begin
    lo0770 <= li0770 ;
 end
 always @ (posedge ) begin
    lo0771 <= li0771 ;
 end
 always @ (posedge ) begin
    lo0772 <= li0772 ;
 end
 always @ (posedge ) begin
    lo0773 <= li0773 ;
 end
 always @ (posedge ) begin
    lo0774 <= li0774 ;
 end
 always @ (posedge ) begin
    lo0775 <= li0775 ;
 end
 always @ (posedge ) begin
    lo0776 <= li0776 ;
 end
 always @ (posedge ) begin
    lo0777 <= li0777 ;
 end
 always @ (posedge ) begin
    lo0778 <= li0778 ;
 end
 always @ (posedge ) begin
    lo0779 <= li0779 ;
 end
 always @ (posedge ) begin
    lo0780 <= li0780 ;
 end
 always @ (posedge ) begin
    lo0781 <= li0781 ;
 end
 always @ (posedge ) begin
    lo0782 <= li0782 ;
 end
 always @ (posedge ) begin
    lo0783 <= li0783 ;
 end
 always @ (posedge ) begin
    lo0784 <= li0784 ;
 end
 always @ (posedge ) begin
    lo0785 <= li0785 ;
 end
 always @ (posedge ) begin
    lo0786 <= li0786 ;
 end
 always @ (posedge ) begin
    lo0787 <= li0787 ;
 end
 always @ (posedge ) begin
    lo0788 <= li0788 ;
 end
 always @ (posedge ) begin
    lo0789 <= li0789 ;
 end
 always @ (posedge ) begin
    lo0790 <= li0790 ;
 end
 always @ (posedge ) begin
    lo0791 <= li0791 ;
 end
 always @ (posedge ) begin
    lo0792 <= li0792 ;
 end
 always @ (posedge ) begin
    lo0793 <= li0793 ;
 end
 always @ (posedge ) begin
    lo0794 <= li0794 ;
 end
 always @ (posedge ) begin
    lo0795 <= li0795 ;
 end
 always @ (posedge ) begin
    lo0796 <= li0796 ;
 end
 always @ (posedge ) begin
    lo0797 <= li0797 ;
 end
 always @ (posedge ) begin
    lo0798 <= li0798 ;
 end
 always @ (posedge ) begin
    lo0799 <= li0799 ;
 end
 always @ (posedge ) begin
    lo0800 <= li0800 ;
 end
 always @ (posedge ) begin
    lo0801 <= li0801 ;
 end
 always @ (posedge ) begin
    lo0802 <= li0802 ;
 end
 always @ (posedge ) begin
    lo0803 <= li0803 ;
 end
 always @ (posedge ) begin
    lo0804 <= li0804 ;
 end
 always @ (posedge ) begin
    lo0805 <= li0805 ;
 end
 always @ (posedge ) begin
    lo0806 <= li0806 ;
 end
 always @ (posedge ) begin
    lo0807 <= li0807 ;
 end
 always @ (posedge ) begin
    lo0808 <= li0808 ;
 end
 always @ (posedge ) begin
    lo0809 <= li0809 ;
 end
 always @ (posedge ) begin
    lo0810 <= li0810 ;
 end
 always @ (posedge ) begin
    lo0811 <= li0811 ;
 end
 always @ (posedge ) begin
    lo0812 <= li0812 ;
 end
 always @ (posedge ) begin
    lo0813 <= li0813 ;
 end
 always @ (posedge ) begin
    lo0814 <= li0814 ;
 end
 always @ (posedge ) begin
    lo0815 <= li0815 ;
 end
 always @ (posedge ) begin
    lo0816 <= li0816 ;
 end
 always @ (posedge ) begin
    lo0817 <= li0817 ;
 end
 always @ (posedge ) begin
    lo0818 <= li0818 ;
 end
 always @ (posedge ) begin
    lo0819 <= li0819 ;
 end
 always @ (posedge ) begin
    lo0820 <= li0820 ;
 end
 always @ (posedge ) begin
    lo0821 <= li0821 ;
 end
 always @ (posedge ) begin
    lo0822 <= li0822 ;
 end
 always @ (posedge ) begin
    lo0823 <= li0823 ;
 end
 always @ (posedge ) begin
    lo0824 <= li0824 ;
 end
 always @ (posedge ) begin
    lo0825 <= li0825 ;
 end
 always @ (posedge ) begin
    lo0826 <= li0826 ;
 end
 always @ (posedge ) begin
    lo0827 <= li0827 ;
 end
 always @ (posedge ) begin
    lo0828 <= li0828 ;
 end
 always @ (posedge ) begin
    lo0829 <= li0829 ;
 end
 always @ (posedge ) begin
    lo0830 <= li0830 ;
 end
 always @ (posedge ) begin
    lo0831 <= li0831 ;
 end
 always @ (posedge ) begin
    lo0832 <= li0832 ;
 end
 always @ (posedge ) begin
    lo0833 <= li0833 ;
 end
 always @ (posedge ) begin
    lo0834 <= li0834 ;
 end
 always @ (posedge ) begin
    lo0835 <= li0835 ;
 end
 always @ (posedge ) begin
    lo0836 <= li0836 ;
 end
 always @ (posedge ) begin
    lo0837 <= li0837 ;
 end
 always @ (posedge ) begin
    lo0838 <= li0838 ;
 end
 always @ (posedge ) begin
    lo0839 <= li0839 ;
 end
 always @ (posedge ) begin
    lo0840 <= li0840 ;
 end
 always @ (posedge ) begin
    lo0841 <= li0841 ;
 end
 always @ (posedge ) begin
    lo0842 <= li0842 ;
 end
 always @ (posedge ) begin
    lo0843 <= li0843 ;
 end
 always @ (posedge ) begin
    lo0844 <= li0844 ;
 end
 always @ (posedge ) begin
    lo0845 <= li0845 ;
 end
 always @ (posedge ) begin
    lo0846 <= li0846 ;
 end
 always @ (posedge ) begin
    lo0847 <= li0847 ;
 end
 always @ (posedge ) begin
    lo0848 <= li0848 ;
 end
 always @ (posedge ) begin
    lo0849 <= li0849 ;
 end
 always @ (posedge ) begin
    lo0850 <= li0850 ;
 end
 always @ (posedge ) begin
    lo0851 <= li0851 ;
 end
 always @ (posedge ) begin
    lo0852 <= li0852 ;
 end
 always @ (posedge ) begin
    lo0853 <= li0853 ;
 end
 always @ (posedge ) begin
    lo0854 <= li0854 ;
 end
 always @ (posedge ) begin
    lo0855 <= li0855 ;
 end
 always @ (posedge ) begin
    lo0856 <= li0856 ;
 end
 always @ (posedge ) begin
    lo0857 <= li0857 ;
 end
 always @ (posedge ) begin
    lo0858 <= li0858 ;
 end
 always @ (posedge ) begin
    lo0859 <= li0859 ;
 end
 always @ (posedge ) begin
    lo0860 <= li0860 ;
 end
 always @ (posedge ) begin
    lo0861 <= li0861 ;
 end
 always @ (posedge ) begin
    lo0862 <= li0862 ;
 end
 always @ (posedge ) begin
    lo0863 <= li0863 ;
 end
 always @ (posedge ) begin
    lo0864 <= li0864 ;
 end
 always @ (posedge ) begin
    lo0865 <= li0865 ;
 end
 always @ (posedge ) begin
    lo0866 <= li0866 ;
 end
 always @ (posedge ) begin
    lo0867 <= li0867 ;
 end
 always @ (posedge ) begin
    lo0868 <= li0868 ;
 end
 always @ (posedge ) begin
    lo0869 <= li0869 ;
 end
 always @ (posedge ) begin
    lo0870 <= li0870 ;
 end
 always @ (posedge ) begin
    lo0871 <= li0871 ;
 end
 always @ (posedge ) begin
    lo0872 <= li0872 ;
 end
 always @ (posedge ) begin
    lo0873 <= li0873 ;
 end
 always @ (posedge ) begin
    lo0874 <= li0874 ;
 end
 always @ (posedge ) begin
    lo0875 <= li0875 ;
 end
 always @ (posedge ) begin
    lo0876 <= li0876 ;
 end
 always @ (posedge ) begin
    lo0877 <= li0877 ;
 end
 always @ (posedge ) begin
    lo0878 <= li0878 ;
 end
 always @ (posedge ) begin
    lo0879 <= li0879 ;
 end
 always @ (posedge ) begin
    lo0880 <= li0880 ;
 end
 always @ (posedge ) begin
    lo0881 <= li0881 ;
 end
 always @ (posedge ) begin
    lo0882 <= li0882 ;
 end
 always @ (posedge ) begin
    lo0883 <= li0883 ;
 end
 always @ (posedge ) begin
    lo0884 <= li0884 ;
 end
 always @ (posedge ) begin
    lo0885 <= li0885 ;
 end
 always @ (posedge ) begin
    lo0886 <= li0886 ;
 end
 always @ (posedge ) begin
    lo0887 <= li0887 ;
 end
 always @ (posedge ) begin
    lo0888 <= li0888 ;
 end
 always @ (posedge ) begin
    lo0889 <= li0889 ;
 end
 always @ (posedge ) begin
    lo0890 <= li0890 ;
 end
 always @ (posedge ) begin
    lo0891 <= li0891 ;
 end
 always @ (posedge ) begin
    lo0892 <= li0892 ;
 end
 always @ (posedge ) begin
    lo0893 <= li0893 ;
 end
 always @ (posedge ) begin
    lo0894 <= li0894 ;
 end
 always @ (posedge ) begin
    lo0895 <= li0895 ;
 end
 always @ (posedge ) begin
    lo0896 <= li0896 ;
 end
 always @ (posedge ) begin
    lo0897 <= li0897 ;
 end
 always @ (posedge ) begin
    lo0898 <= li0898 ;
 end
 always @ (posedge ) begin
    lo0899 <= li0899 ;
 end
 always @ (posedge ) begin
    lo0900 <= li0900 ;
 end
 always @ (posedge ) begin
    lo0901 <= li0901 ;
 end
 always @ (posedge ) begin
    lo0902 <= li0902 ;
 end
 always @ (posedge ) begin
    lo0903 <= li0903 ;
 end
 always @ (posedge ) begin
    lo0904 <= li0904 ;
 end
 always @ (posedge ) begin
    lo0905 <= li0905 ;
 end
 always @ (posedge ) begin
    lo0906 <= li0906 ;
 end
 always @ (posedge ) begin
    lo0907 <= li0907 ;
 end
 always @ (posedge ) begin
    lo0908 <= li0908 ;
 end
 always @ (posedge ) begin
    lo0909 <= li0909 ;
 end
 always @ (posedge ) begin
    lo0910 <= li0910 ;
 end
 always @ (posedge ) begin
    lo0911 <= li0911 ;
 end
 always @ (posedge ) begin
    lo0912 <= li0912 ;
 end
 always @ (posedge ) begin
    lo0913 <= li0913 ;
 end
 always @ (posedge ) begin
    lo0914 <= li0914 ;
 end
 always @ (posedge ) begin
    lo0915 <= li0915 ;
 end
 always @ (posedge ) begin
    lo0916 <= li0916 ;
 end
 always @ (posedge ) begin
    lo0917 <= li0917 ;
 end
 always @ (posedge ) begin
    lo0918 <= li0918 ;
 end
 always @ (posedge ) begin
    lo0919 <= li0919 ;
 end
 always @ (posedge ) begin
    lo0920 <= li0920 ;
 end
 always @ (posedge ) begin
    lo0921 <= li0921 ;
 end
 always @ (posedge ) begin
    lo0922 <= li0922 ;
 end
 always @ (posedge ) begin
    lo0923 <= li0923 ;
 end
 always @ (posedge ) begin
    lo0924 <= li0924 ;
 end
 always @ (posedge ) begin
    lo0925 <= li0925 ;
 end
 always @ (posedge ) begin
    lo0926 <= li0926 ;
 end
 always @ (posedge ) begin
    lo0927 <= li0927 ;
 end
 always @ (posedge ) begin
    lo0928 <= li0928 ;
 end
 always @ (posedge ) begin
    lo0929 <= li0929 ;
 end
 always @ (posedge ) begin
    lo0930 <= li0930 ;
 end
 always @ (posedge ) begin
    lo0931 <= li0931 ;
 end
 always @ (posedge ) begin
    lo0932 <= li0932 ;
 end
 always @ (posedge ) begin
    lo0933 <= li0933 ;
 end
 always @ (posedge ) begin
    lo0934 <= li0934 ;
 end
 always @ (posedge ) begin
    lo0935 <= li0935 ;
 end
 always @ (posedge ) begin
    lo0936 <= li0936 ;
 end
 always @ (posedge ) begin
    lo0937 <= li0937 ;
 end
 always @ (posedge ) begin
    lo0938 <= li0938 ;
 end
 always @ (posedge ) begin
    lo0939 <= li0939 ;
 end
 always @ (posedge ) begin
    lo0940 <= li0940 ;
 end
 always @ (posedge ) begin
    lo0941 <= li0941 ;
 end
 always @ (posedge ) begin
    lo0942 <= li0942 ;
 end
 always @ (posedge ) begin
    lo0943 <= li0943 ;
 end
 always @ (posedge ) begin
    lo0944 <= li0944 ;
 end
 always @ (posedge ) begin
    lo0945 <= li0945 ;
 end
 always @ (posedge ) begin
    lo0946 <= li0946 ;
 end
 always @ (posedge ) begin
    lo0947 <= li0947 ;
 end
 always @ (posedge ) begin
    lo0948 <= li0948 ;
 end
 always @ (posedge ) begin
    lo0949 <= li0949 ;
 end
 always @ (posedge ) begin
    lo0950 <= li0950 ;
 end
 always @ (posedge ) begin
    lo0951 <= li0951 ;
 end
 always @ (posedge ) begin
    lo0952 <= li0952 ;
 end
 always @ (posedge ) begin
    lo0953 <= li0953 ;
 end
 always @ (posedge ) begin
    lo0954 <= li0954 ;
 end
 always @ (posedge ) begin
    lo0955 <= li0955 ;
 end
 always @ (posedge ) begin
    lo0956 <= li0956 ;
 end
 always @ (posedge ) begin
    lo0957 <= li0957 ;
 end
 always @ (posedge ) begin
    lo0958 <= li0958 ;
 end
 always @ (posedge ) begin
    lo0959 <= li0959 ;
 end
 always @ (posedge ) begin
    lo0960 <= li0960 ;
 end
 always @ (posedge ) begin
    lo0961 <= li0961 ;
 end
 always @ (posedge ) begin
    lo0962 <= li0962 ;
 end
 always @ (posedge ) begin
    lo0963 <= li0963 ;
 end
 always @ (posedge ) begin
    lo0964 <= li0964 ;
 end
 always @ (posedge ) begin
    lo0965 <= li0965 ;
 end
 always @ (posedge ) begin
    lo0966 <= li0966 ;
 end
 always @ (posedge ) begin
    lo0967 <= li0967 ;
 end
 always @ (posedge ) begin
    lo0968 <= li0968 ;
 end
 always @ (posedge ) begin
    lo0969 <= li0969 ;
 end
 always @ (posedge ) begin
    lo0970 <= li0970 ;
 end
 always @ (posedge ) begin
    lo0971 <= li0971 ;
 end
 always @ (posedge ) begin
    lo0972 <= li0972 ;
 end
 always @ (posedge ) begin
    lo0973 <= li0973 ;
 end
 always @ (posedge ) begin
    lo0974 <= li0974 ;
 end
 always @ (posedge ) begin
    lo0975 <= li0975 ;
 end
 always @ (posedge ) begin
    lo0976 <= li0976 ;
 end
 always @ (posedge ) begin
    lo0977 <= li0977 ;
 end
 always @ (posedge ) begin
    lo0978 <= li0978 ;
 end
 always @ (posedge ) begin
    lo0979 <= li0979 ;
 end
 always @ (posedge ) begin
    lo0980 <= li0980 ;
 end
 always @ (posedge ) begin
    lo0981 <= li0981 ;
 end
 always @ (posedge ) begin
    lo0982 <= li0982 ;
 end
 always @ (posedge ) begin
    lo0983 <= li0983 ;
 end
 always @ (posedge ) begin
    lo0984 <= li0984 ;
 end
 always @ (posedge ) begin
    lo0985 <= li0985 ;
 end
 always @ (posedge ) begin
    lo0986 <= li0986 ;
 end
 always @ (posedge ) begin
    lo0987 <= li0987 ;
 end
 always @ (posedge ) begin
    lo0988 <= li0988 ;
 end
 always @ (posedge ) begin
    lo0989 <= li0989 ;
 end
 always @ (posedge ) begin
    lo0990 <= li0990 ;
 end
 always @ (posedge ) begin
    lo0991 <= li0991 ;
 end
 always @ (posedge ) begin
    lo0992 <= li0992 ;
 end
 always @ (posedge ) begin
    lo0993 <= li0993 ;
 end
 always @ (posedge ) begin
    lo0994 <= li0994 ;
 end
 always @ (posedge ) begin
    lo0995 <= li0995 ;
 end
 always @ (posedge ) begin
    lo0996 <= li0996 ;
 end
 always @ (posedge ) begin
    lo0997 <= li0997 ;
 end
 always @ (posedge ) begin
    lo0998 <= li0998 ;
 end
 always @ (posedge ) begin
    lo0999 <= li0999 ;
 end
 always @ (posedge ) begin
    lo1000 <= li1000 ;
 end
 always @ (posedge ) begin
    lo1001 <= li1001 ;
 end
 always @ (posedge ) begin
    lo1002 <= li1002 ;
 end
 always @ (posedge ) begin
    lo1003 <= li1003 ;
 end
 always @ (posedge ) begin
    lo1004 <= li1004 ;
 end
 always @ (posedge ) begin
    lo1005 <= li1005 ;
 end
 always @ (posedge ) begin
    lo1006 <= li1006 ;
 end
 always @ (posedge ) begin
    lo1007 <= li1007 ;
 end
 always @ (posedge ) begin
    lo1008 <= li1008 ;
 end
 always @ (posedge ) begin
    lo1009 <= li1009 ;
 end
 always @ (posedge ) begin
    lo1010 <= li1010 ;
 end
 always @ (posedge ) begin
    lo1011 <= li1011 ;
 end
 always @ (posedge ) begin
    lo1012 <= li1012 ;
 end
 always @ (posedge ) begin
    lo1013 <= li1013 ;
 end
 always @ (posedge ) begin
    lo1014 <= li1014 ;
 end
 always @ (posedge ) begin
    lo1015 <= li1015 ;
 end
 always @ (posedge ) begin
    lo1016 <= li1016 ;
 end
 always @ (posedge ) begin
    lo1017 <= li1017 ;
 end
 always @ (posedge ) begin
    lo1018 <= li1018 ;
 end
 always @ (posedge ) begin
    lo1019 <= li1019 ;
 end
 always @ (posedge ) begin
    lo1020 <= li1020 ;
 end
 always @ (posedge ) begin
    lo1021 <= li1021 ;
 end
 always @ (posedge ) begin
    lo1022 <= li1022 ;
 end
 always @ (posedge ) begin
    lo1023 <= li1023 ;
 end
 always @ (posedge ) begin
    lo1024 <= li1024 ;
 end
 always @ (posedge ) begin
    lo1025 <= li1025 ;
 end
 always @ (posedge ) begin
    lo1026 <= li1026 ;
 end
 always @ (posedge ) begin
    lo1027 <= li1027 ;
 end
 always @ (posedge ) begin
    lo1028 <= li1028 ;
 end
 always @ (posedge ) begin
    lo1029 <= li1029 ;
 end
 always @ (posedge ) begin
    lo1030 <= li1030 ;
 end
 always @ (posedge ) begin
    lo1031 <= li1031 ;
 end
 always @ (posedge ) begin
    lo1032 <= li1032 ;
 end
 always @ (posedge ) begin
    lo1033 <= li1033 ;
 end
 always @ (posedge ) begin
    lo1034 <= li1034 ;
 end
 always @ (posedge ) begin
    lo1035 <= li1035 ;
 end
 always @ (posedge ) begin
    lo1036 <= li1036 ;
 end
 always @ (posedge ) begin
    lo1037 <= li1037 ;
 end
 always @ (posedge ) begin
    lo1038 <= li1038 ;
 end
 always @ (posedge ) begin
    lo1039 <= li1039 ;
 end
 always @ (posedge ) begin
    lo1040 <= li1040 ;
 end
 always @ (posedge ) begin
    lo1041 <= li1041 ;
 end
 always @ (posedge ) begin
    lo1042 <= li1042 ;
 end
 always @ (posedge ) begin
    lo1043 <= li1043 ;
 end
 always @ (posedge ) begin
    lo1044 <= li1044 ;
 end
 always @ (posedge ) begin
    lo1045 <= li1045 ;
 end
 always @ (posedge ) begin
    lo1046 <= li1046 ;
 end
 always @ (posedge ) begin
    lo1047 <= li1047 ;
 end
 always @ (posedge ) begin
    lo1048 <= li1048 ;
 end
 always @ (posedge ) begin
    lo1049 <= li1049 ;
 end
 always @ (posedge ) begin
    lo1050 <= li1050 ;
 end
 always @ (posedge ) begin
    lo1051 <= li1051 ;
 end
 always @ (posedge ) begin
    lo1052 <= li1052 ;
 end
 always @ (posedge ) begin
    lo1053 <= li1053 ;
 end
 always @ (posedge ) begin
    lo1054 <= li1054 ;
 end
 always @ (posedge ) begin
    lo1055 <= li1055 ;
 end
 always @ (posedge ) begin
    lo1056 <= li1056 ;
 end
 always @ (posedge ) begin
    lo1057 <= li1057 ;
 end
 always @ (posedge ) begin
    lo1058 <= li1058 ;
 end
 always @ (posedge ) begin
    lo1059 <= li1059 ;
 end
 always @ (posedge ) begin
    lo1060 <= li1060 ;
 end
 always @ (posedge ) begin
    lo1061 <= li1061 ;
 end
 always @ (posedge ) begin
    lo1062 <= li1062 ;
 end
 always @ (posedge ) begin
    lo1063 <= li1063 ;
 end
 always @ (posedge ) begin
    lo1064 <= li1064 ;
 end
 always @ (posedge ) begin
    lo1065 <= li1065 ;
 end
 always @ (posedge ) begin
    lo1066 <= li1066 ;
 end
 always @ (posedge ) begin
    lo1067 <= li1067 ;
 end
 always @ (posedge ) begin
    lo1068 <= li1068 ;
 end
 always @ (posedge ) begin
    lo1069 <= li1069 ;
 end
 always @ (posedge ) begin
    lo1070 <= li1070 ;
 end
 always @ (posedge ) begin
    lo1071 <= li1071 ;
 end
 always @ (posedge ) begin
    lo1072 <= li1072 ;
 end
 always @ (posedge ) begin
    lo1073 <= li1073 ;
 end
 always @ (posedge ) begin
    lo1074 <= li1074 ;
 end
 always @ (posedge ) begin
    lo1075 <= li1075 ;
 end
 always @ (posedge ) begin
    lo1076 <= li1076 ;
 end
 always @ (posedge ) begin
    lo1077 <= li1077 ;
 end
 always @ (posedge ) begin
    lo1078 <= li1078 ;
 end
 always @ (posedge ) begin
    lo1079 <= li1079 ;
 end
 always @ (posedge ) begin
    lo1080 <= li1080 ;
 end
 always @ (posedge ) begin
    lo1081 <= li1081 ;
 end
 always @ (posedge ) begin
    lo1082 <= li1082 ;
 end
 always @ (posedge ) begin
    lo1083 <= li1083 ;
 end
 always @ (posedge ) begin
    lo1084 <= li1084 ;
 end
 always @ (posedge ) begin
    lo1085 <= li1085 ;
 end
 always @ (posedge ) begin
    lo1086 <= li1086 ;
 end
 always @ (posedge ) begin
    lo1087 <= li1087 ;
 end
 always @ (posedge ) begin
    lo1088 <= li1088 ;
 end
 always @ (posedge ) begin
    lo1089 <= li1089 ;
 end
 always @ (posedge ) begin
    lo1090 <= li1090 ;
 end
 always @ (posedge ) begin
    lo1091 <= li1091 ;
 end
 always @ (posedge ) begin
    lo1092 <= li1092 ;
 end
 always @ (posedge ) begin
    lo1093 <= li1093 ;
 end
 always @ (posedge ) begin
    lo1094 <= li1094 ;
 end
 always @ (posedge ) begin
    lo1095 <= li1095 ;
 end
 always @ (posedge ) begin
    lo1096 <= li1096 ;
 end
 always @ (posedge ) begin
    lo1097 <= li1097 ;
 end
 always @ (posedge ) begin
    lo1098 <= li1098 ;
 end
 always @ (posedge ) begin
    lo1099 <= li1099 ;
 end
 always @ (posedge ) begin
    lo1100 <= li1100 ;
 end
 always @ (posedge ) begin
    lo1101 <= li1101 ;
 end
 always @ (posedge ) begin
    lo1102 <= li1102 ;
 end
 always @ (posedge ) begin
    lo1103 <= li1103 ;
 end
 always @ (posedge ) begin
    lo1104 <= li1104 ;
 end
 always @ (posedge ) begin
    lo1105 <= li1105 ;
 end
 always @ (posedge ) begin
    lo1106 <= li1106 ;
 end
 always @ (posedge ) begin
    lo1107 <= li1107 ;
 end
 always @ (posedge ) begin
    lo1108 <= li1108 ;
 end
 always @ (posedge ) begin
    lo1109 <= li1109 ;
 end
 always @ (posedge ) begin
    lo1110 <= li1110 ;
 end
 always @ (posedge ) begin
    lo1111 <= li1111 ;
 end
 always @ (posedge ) begin
    lo1112 <= li1112 ;
 end
 always @ (posedge ) begin
    lo1113 <= li1113 ;
 end
 always @ (posedge ) begin
    lo1114 <= li1114 ;
 end
 always @ (posedge ) begin
    lo1115 <= li1115 ;
 end
 always @ (posedge ) begin
    lo1116 <= li1116 ;
 end
 always @ (posedge ) begin
    lo1117 <= li1117 ;
 end
 always @ (posedge ) begin
    lo1118 <= li1118 ;
 end
 always @ (posedge ) begin
    lo1119 <= li1119 ;
 end
 always @ (posedge ) begin
    lo1120 <= li1120 ;
 end
 always @ (posedge ) begin
    lo1121 <= li1121 ;
 end
 always @ (posedge ) begin
    lo1122 <= li1122 ;
 end
 always @ (posedge ) begin
    lo1123 <= li1123 ;
 end
 always @ (posedge ) begin
    lo1124 <= li1124 ;
 end
 always @ (posedge ) begin
    lo1125 <= li1125 ;
 end
 always @ (posedge ) begin
    lo1126 <= li1126 ;
 end
 always @ (posedge ) begin
    lo1127 <= li1127 ;
 end
 always @ (posedge ) begin
    lo1128 <= li1128 ;
 end
 always @ (posedge ) begin
    lo1129 <= li1129 ;
 end
 always @ (posedge ) begin
    lo1130 <= li1130 ;
 end
 always @ (posedge ) begin
    lo1131 <= li1131 ;
 end
 always @ (posedge ) begin
    lo1132 <= li1132 ;
 end
 always @ (posedge ) begin
    lo1133 <= li1133 ;
 end
 always @ (posedge ) begin
    lo1134 <= li1134 ;
 end
 always @ (posedge ) begin
    lo1135 <= li1135 ;
 end
 always @ (posedge ) begin
    lo1136 <= li1136 ;
 end
 always @ (posedge ) begin
    lo1137 <= li1137 ;
 end
 always @ (posedge ) begin
    lo1138 <= li1138 ;
 end
 always @ (posedge ) begin
    lo1139 <= li1139 ;
 end
 always @ (posedge ) begin
    lo1140 <= li1140 ;
 end
 always @ (posedge ) begin
    lo1141 <= li1141 ;
 end
 always @ (posedge ) begin
    lo1142 <= li1142 ;
 end
 always @ (posedge ) begin
    lo1143 <= li1143 ;
 end
 always @ (posedge ) begin
    lo1144 <= li1144 ;
 end
 always @ (posedge ) begin
    lo1145 <= li1145 ;
 end
 always @ (posedge ) begin
    lo1146 <= li1146 ;
 end
 always @ (posedge ) begin
    lo1147 <= li1147 ;
 end
 always @ (posedge ) begin
    lo1148 <= li1148 ;
 end
 always @ (posedge ) begin
    lo1149 <= li1149 ;
 end
 always @ (posedge ) begin
    lo1150 <= li1150 ;
 end
 always @ (posedge ) begin
    lo1151 <= li1151 ;
 end
 always @ (posedge ) begin
    lo1152 <= li1152 ;
 end
 always @ (posedge ) begin
    lo1153 <= li1153 ;
 end
 always @ (posedge ) begin
    lo1154 <= li1154 ;
 end
 always @ (posedge ) begin
    lo1155 <= li1155 ;
 end
 always @ (posedge ) begin
    lo1156 <= li1156 ;
 end
 always @ (posedge ) begin
    lo1157 <= li1157 ;
 end
 always @ (posedge ) begin
    lo1158 <= li1158 ;
 end
 always @ (posedge ) begin
    lo1159 <= li1159 ;
 end
 always @ (posedge ) begin
    lo1160 <= li1160 ;
 end
 always @ (posedge ) begin
    lo1161 <= li1161 ;
 end
 always @ (posedge ) begin
    lo1162 <= li1162 ;
 end
 always @ (posedge ) begin
    lo1163 <= li1163 ;
 end
 always @ (posedge ) begin
    lo1164 <= li1164 ;
 end
 always @ (posedge ) begin
    lo1165 <= li1165 ;
 end
 always @ (posedge ) begin
    lo1166 <= li1166 ;
 end
 always @ (posedge ) begin
    lo1167 <= li1167 ;
 end
 always @ (posedge ) begin
    lo1168 <= li1168 ;
 end
 always @ (posedge ) begin
    lo1169 <= li1169 ;
 end
 always @ (posedge ) begin
    lo1170 <= li1170 ;
 end
 always @ (posedge ) begin
    lo1171 <= li1171 ;
 end
 always @ (posedge ) begin
    lo1172 <= li1172 ;
 end
 always @ (posedge ) begin
    lo1173 <= li1173 ;
 end
 always @ (posedge ) begin
    lo1174 <= li1174 ;
 end
 always @ (posedge ) begin
    lo1175 <= li1175 ;
 end
 always @ (posedge ) begin
    lo1176 <= li1176 ;
 end
 always @ (posedge ) begin
    lo1177 <= li1177 ;
 end
 always @ (posedge ) begin
    lo1178 <= li1178 ;
 end
 always @ (posedge ) begin
    lo1179 <= li1179 ;
 end
 always @ (posedge ) begin
    lo1180 <= li1180 ;
 end
 always @ (posedge ) begin
    lo1181 <= li1181 ;
 end
 always @ (posedge ) begin
    lo1182 <= li1182 ;
 end
 always @ (posedge ) begin
    lo1183 <= li1183 ;
 end
 always @ (posedge ) begin
    lo1184 <= li1184 ;
 end
 always @ (posedge ) begin
    lo1185 <= li1185 ;
 end
 always @ (posedge ) begin
    lo1186 <= li1186 ;
 end
 always @ (posedge ) begin
    lo1187 <= li1187 ;
 end
 always @ (posedge ) begin
    lo1188 <= li1188 ;
 end
 always @ (posedge ) begin
    lo1189 <= li1189 ;
 end
 always @ (posedge ) begin
    lo1190 <= li1190 ;
 end
 always @ (posedge ) begin
    lo1191 <= li1191 ;
 end
 always @ (posedge ) begin
    lo1192 <= li1192 ;
 end
 always @ (posedge ) begin
    lo1193 <= li1193 ;
 end
 always @ (posedge ) begin
    lo1194 <= li1194 ;
 end
 always @ (posedge ) begin
    lo1195 <= li1195 ;
 end
 always @ (posedge ) begin
    lo1196 <= li1196 ;
 end
 always @ (posedge ) begin
    lo1197 <= li1197 ;
 end
 always @ (posedge ) begin
    lo1198 <= li1198 ;
 end
 always @ (posedge ) begin
    lo1199 <= li1199 ;
 end
 always @ (posedge ) begin
    lo1200 <= li1200 ;
 end
 always @ (posedge ) begin
    lo1201 <= li1201 ;
 end
 always @ (posedge ) begin
    lo1202 <= li1202 ;
 end
 always @ (posedge ) begin
    lo1203 <= li1203 ;
 end
 always @ (posedge ) begin
    lo1204 <= li1204 ;
 end
 always @ (posedge ) begin
    lo1205 <= li1205 ;
 end
 always @ (posedge ) begin
    lo1206 <= li1206 ;
 end
 always @ (posedge ) begin
    lo1207 <= li1207 ;
 end
 always @ (posedge ) begin
    lo1208 <= li1208 ;
 end
 always @ (posedge ) begin
    lo1209 <= li1209 ;
 end
 always @ (posedge ) begin
    lo1210 <= li1210 ;
 end
 always @ (posedge ) begin
    lo1211 <= li1211 ;
 end
 always @ (posedge ) begin
    lo1212 <= li1212 ;
 end
 always @ (posedge ) begin
    lo1213 <= li1213 ;
 end
 always @ (posedge ) begin
    lo1214 <= li1214 ;
 end
 always @ (posedge ) begin
    lo1215 <= li1215 ;
 end
 always @ (posedge ) begin
    lo1216 <= li1216 ;
 end
 always @ (posedge ) begin
    lo1217 <= li1217 ;
 end
 always @ (posedge ) begin
    lo1218 <= li1218 ;
 end
 always @ (posedge ) begin
    lo1219 <= li1219 ;
 end
 always @ (posedge ) begin
    lo1220 <= li1220 ;
 end
 always @ (posedge ) begin
    lo1221 <= li1221 ;
 end
 always @ (posedge ) begin
    lo1222 <= li1222 ;
 end
 always @ (posedge ) begin
    lo1223 <= li1223 ;
 end
 always @ (posedge ) begin
    lo1224 <= li1224 ;
 end
 always @ (posedge ) begin
    lo1225 <= li1225 ;
 end
 always @ (posedge ) begin
    lo1226 <= li1226 ;
 end
 always @ (posedge ) begin
    lo1227 <= li1227 ;
 end
 always @ (posedge ) begin
    lo1228 <= li1228 ;
 end
 always @ (posedge ) begin
    lo1229 <= li1229 ;
 end
 always @ (posedge ) begin
    lo1230 <= li1230 ;
 end
 always @ (posedge ) begin
    lo1231 <= li1231 ;
 end
 always @ (posedge ) begin
    lo1232 <= li1232 ;
 end
 always @ (posedge ) begin
    lo1233 <= li1233 ;
 end
 always @ (posedge ) begin
    lo1234 <= li1234 ;
 end
 always @ (posedge ) begin
    lo1235 <= li1235 ;
 end
 always @ (posedge ) begin
    lo1236 <= li1236 ;
 end
 always @ (posedge ) begin
    lo1237 <= li1237 ;
 end
 always @ (posedge ) begin
    lo1238 <= li1238 ;
 end
 always @ (posedge ) begin
    lo1239 <= li1239 ;
 end
 always @ (posedge ) begin
    lo1240 <= li1240 ;
 end
 always @ (posedge ) begin
    lo1241 <= li1241 ;
 end
 always @ (posedge ) begin
    lo1242 <= li1242 ;
 end
 always @ (posedge ) begin
    lo1243 <= li1243 ;
 end
 always @ (posedge ) begin
    lo1244 <= li1244 ;
 end
 always @ (posedge ) begin
    lo1245 <= li1245 ;
 end
 always @ (posedge ) begin
    lo1246 <= li1246 ;
 end
 always @ (posedge ) begin
    lo1247 <= li1247 ;
 end
 always @ (posedge ) begin
    lo1248 <= li1248 ;
 end
 always @ (posedge ) begin
    lo1249 <= li1249 ;
 end
 always @ (posedge ) begin
    lo1250 <= li1250 ;
 end
 always @ (posedge ) begin
    lo1251 <= li1251 ;
 end
 always @ (posedge ) begin
    lo1252 <= li1252 ;
 end
 always @ (posedge ) begin
    lo1253 <= li1253 ;
 end
 always @ (posedge ) begin
    lo1254 <= li1254 ;
 end
 always @ (posedge ) begin
    lo1255 <= li1255 ;
 end
 always @ (posedge ) begin
    lo1256 <= li1256 ;
 end
 always @ (posedge ) begin
    lo1257 <= li1257 ;
 end
 always @ (posedge ) begin
    lo1258 <= li1258 ;
 end
 always @ (posedge ) begin
    lo1259 <= li1259 ;
 end
 always @ (posedge ) begin
    lo1260 <= li1260 ;
 end
 always @ (posedge ) begin
    lo1261 <= li1261 ;
 end
 always @ (posedge ) begin
    lo1262 <= li1262 ;
 end
 always @ (posedge ) begin
    lo1263 <= li1263 ;
 end
 always @ (posedge ) begin
    lo1264 <= li1264 ;
 end
 always @ (posedge ) begin
    lo1265 <= li1265 ;
 end
 always @ (posedge ) begin
    lo1266 <= li1266 ;
 end
 always @ (posedge ) begin
    lo1267 <= li1267 ;
 end
 always @ (posedge ) begin
    lo1268 <= li1268 ;
 end
 always @ (posedge ) begin
    lo1269 <= li1269 ;
 end
 always @ (posedge ) begin
    lo1270 <= li1270 ;
 end
 always @ (posedge ) begin
    lo1271 <= li1271 ;
 end
 always @ (posedge ) begin
    lo1272 <= li1272 ;
 end
 always @ (posedge ) begin
    lo1273 <= li1273 ;
 end
 always @ (posedge ) begin
    lo1274 <= li1274 ;
 end
 always @ (posedge ) begin
    lo1275 <= li1275 ;
 end
 always @ (posedge ) begin
    lo1276 <= li1276 ;
 end
 always @ (posedge ) begin
    lo1277 <= li1277 ;
 end
 always @ (posedge ) begin
    lo1278 <= li1278 ;
 end
 always @ (posedge ) begin
    lo1279 <= li1279 ;
 end
 always @ (posedge ) begin
    lo1280 <= li1280 ;
 end
 always @ (posedge ) begin
    lo1281 <= li1281 ;
 end
 always @ (posedge ) begin
    lo1282 <= li1282 ;
 end
 always @ (posedge ) begin
    lo1283 <= li1283 ;
 end
 always @ (posedge ) begin
    lo1284 <= li1284 ;
 end
 always @ (posedge ) begin
    lo1285 <= li1285 ;
 end
 always @ (posedge ) begin
    lo1286 <= li1286 ;
 end
 always @ (posedge ) begin
    lo1287 <= li1287 ;
 end
 always @ (posedge ) begin
    lo1288 <= li1288 ;
 end
 always @ (posedge ) begin
    lo1289 <= li1289 ;
 end
 always @ (posedge ) begin
    lo1290 <= li1290 ;
 end
 always @ (posedge ) begin
    lo1291 <= li1291 ;
 end
 always @ (posedge ) begin
    lo1292 <= li1292 ;
 end
 always @ (posedge ) begin
    lo1293 <= li1293 ;
 end
 always @ (posedge ) begin
    lo1294 <= li1294 ;
 end
 always @ (posedge ) begin
    lo1295 <= li1295 ;
 end
 always @ (posedge ) begin
    lo1296 <= li1296 ;
 end
 always @ (posedge ) begin
    lo1297 <= li1297 ;
 end
 always @ (posedge ) begin
    lo1298 <= li1298 ;
 end
 always @ (posedge ) begin
    lo1299 <= li1299 ;
 end
 always @ (posedge ) begin
    lo1300 <= li1300 ;
 end
 always @ (posedge ) begin
    lo1301 <= li1301 ;
 end
 always @ (posedge ) begin
    lo1302 <= li1302 ;
 end
 always @ (posedge ) begin
    lo1303 <= li1303 ;
 end
 always @ (posedge ) begin
    lo1304 <= li1304 ;
 end
 always @ (posedge ) begin
    lo1305 <= li1305 ;
 end
 always @ (posedge ) begin
    lo1306 <= li1306 ;
 end
 always @ (posedge ) begin
    lo1307 <= li1307 ;
 end
 always @ (posedge ) begin
    lo1308 <= li1308 ;
 end
 always @ (posedge ) begin
    lo1309 <= li1309 ;
 end
 always @ (posedge ) begin
    lo1310 <= li1310 ;
 end
 always @ (posedge ) begin
    lo1311 <= li1311 ;
 end
 always @ (posedge ) begin
    lo1312 <= li1312 ;
 end
 always @ (posedge ) begin
    lo1313 <= li1313 ;
 end
 always @ (posedge ) begin
    lo1314 <= li1314 ;
 end
 always @ (posedge ) begin
    lo1315 <= li1315 ;
 end
 always @ (posedge ) begin
    lo1316 <= li1316 ;
 end
 always @ (posedge ) begin
    lo1317 <= li1317 ;
 end
 always @ (posedge ) begin
    lo1318 <= li1318 ;
 end
 always @ (posedge ) begin
    lo1319 <= li1319 ;
 end
 always @ (posedge ) begin
    lo1320 <= li1320 ;
 end
 always @ (posedge ) begin
    lo1321 <= li1321 ;
 end
 always @ (posedge ) begin
    lo1322 <= li1322 ;
 end
 always @ (posedge ) begin
    lo1323 <= li1323 ;
 end
 always @ (posedge ) begin
    lo1324 <= li1324 ;
 end
 always @ (posedge ) begin
    lo1325 <= li1325 ;
 end
 always @ (posedge ) begin
    lo1326 <= li1326 ;
 end
 always @ (posedge ) begin
    lo1327 <= li1327 ;
 end
 always @ (posedge ) begin
    lo1328 <= li1328 ;
 end
 always @ (posedge ) begin
    lo1329 <= li1329 ;
 end
 always @ (posedge ) begin
    lo1330 <= li1330 ;
 end
 always @ (posedge ) begin
    lo1331 <= li1331 ;
 end
 always @ (posedge ) begin
    lo1332 <= li1332 ;
 end
 always @ (posedge ) begin
    lo1333 <= li1333 ;
 end
 always @ (posedge ) begin
    lo1334 <= li1334 ;
 end
 always @ (posedge ) begin
    lo1335 <= li1335 ;
 end
 always @ (posedge ) begin
    lo1336 <= li1336 ;
 end
 always @ (posedge ) begin
    lo1337 <= li1337 ;
 end
 always @ (posedge ) begin
    lo1338 <= li1338 ;
 end
 always @ (posedge ) begin
    lo1339 <= li1339 ;
 end
 always @ (posedge ) begin
    lo1340 <= li1340 ;
 end
 always @ (posedge ) begin
    lo1341 <= li1341 ;
 end
 always @ (posedge ) begin
    lo1342 <= li1342 ;
 end
 always @ (posedge ) begin
    lo1343 <= li1343 ;
 end
 always @ (posedge ) begin
    lo1344 <= li1344 ;
 end
 always @ (posedge ) begin
    lo1345 <= li1345 ;
 end
 always @ (posedge ) begin
    lo1346 <= li1346 ;
 end
 always @ (posedge ) begin
    lo1347 <= li1347 ;
 end
 always @ (posedge ) begin
    lo1348 <= li1348 ;
 end
 always @ (posedge ) begin
    lo1349 <= li1349 ;
 end
 always @ (posedge ) begin
    lo1350 <= li1350 ;
 end
 always @ (posedge ) begin
    lo1351 <= li1351 ;
 end
 always @ (posedge ) begin
    lo1352 <= li1352 ;
 end
 always @ (posedge ) begin
    lo1353 <= li1353 ;
 end
 always @ (posedge ) begin
    lo1354 <= li1354 ;
 end
 always @ (posedge ) begin
    lo1355 <= li1355 ;
 end
 always @ (posedge ) begin
    lo1356 <= li1356 ;
 end
 always @ (posedge ) begin
    lo1357 <= li1357 ;
 end
 always @ (posedge ) begin
    lo1358 <= li1358 ;
 end
 always @ (posedge ) begin
    lo1359 <= li1359 ;
 end
 always @ (posedge ) begin
    lo1360 <= li1360 ;
 end
 always @ (posedge ) begin
    lo1361 <= li1361 ;
 end
 always @ (posedge ) begin
    lo1362 <= li1362 ;
 end
 always @ (posedge ) begin
    lo1363 <= li1363 ;
 end
 always @ (posedge ) begin
    lo1364 <= li1364 ;
 end
 always @ (posedge ) begin
    lo1365 <= li1365 ;
 end
 always @ (posedge ) begin
    lo1366 <= li1366 ;
 end
 always @ (posedge ) begin
    lo1367 <= li1367 ;
 end
 always @ (posedge ) begin
    lo1368 <= li1368 ;
 end
 always @ (posedge ) begin
    lo1369 <= li1369 ;
 end
 always @ (posedge ) begin
    lo1370 <= li1370 ;
 end
 always @ (posedge ) begin
    lo1371 <= li1371 ;
 end
 always @ (posedge ) begin
    lo1372 <= li1372 ;
 end
 always @ (posedge ) begin
    lo1373 <= li1373 ;
 end
 always @ (posedge ) begin
    lo1374 <= li1374 ;
 end
 always @ (posedge ) begin
    lo1375 <= li1375 ;
 end
 always @ (posedge ) begin
    lo1376 <= li1376 ;
 end
 always @ (posedge ) begin
    lo1377 <= li1377 ;
 end
 always @ (posedge ) begin
    lo1378 <= li1378 ;
 end
 always @ (posedge ) begin
    lo1379 <= li1379 ;
 end
 always @ (posedge ) begin
    lo1380 <= li1380 ;
 end
 always @ (posedge ) begin
    lo1381 <= li1381 ;
 end
 always @ (posedge ) begin
    lo1382 <= li1382 ;
 end
 always @ (posedge ) begin
    lo1383 <= li1383 ;
 end
 always @ (posedge ) begin
    lo1384 <= li1384 ;
 end
 always @ (posedge ) begin
    lo1385 <= li1385 ;
 end
 always @ (posedge ) begin
    lo1386 <= li1386 ;
 end
 always @ (posedge ) begin
    lo1387 <= li1387 ;
 end
 always @ (posedge ) begin
    lo1388 <= li1388 ;
 end
 always @ (posedge ) begin
    lo1389 <= li1389 ;
 end
 always @ (posedge ) begin
    lo1390 <= li1390 ;
 end
 always @ (posedge ) begin
    lo1391 <= li1391 ;
 end
 always @ (posedge ) begin
    lo1392 <= li1392 ;
 end
 always @ (posedge ) begin
    lo1393 <= li1393 ;
 end
 always @ (posedge ) begin
    lo1394 <= li1394 ;
 end
 always @ (posedge ) begin
    lo1395 <= li1395 ;
 end
 always @ (posedge ) begin
    lo1396 <= li1396 ;
 end
 always @ (posedge ) begin
    lo1397 <= li1397 ;
 end
 always @ (posedge ) begin
    lo1398 <= li1398 ;
 end
 always @ (posedge ) begin
    lo1399 <= li1399 ;
 end
 always @ (posedge ) begin
    lo1400 <= li1400 ;
 end
 always @ (posedge ) begin
    lo1401 <= li1401 ;
 end
 always @ (posedge ) begin
    lo1402 <= li1402 ;
 end
 always @ (posedge ) begin
    lo1403 <= li1403 ;
 end
 always @ (posedge ) begin
    lo1404 <= li1404 ;
 end
 always @ (posedge ) begin
    lo1405 <= li1405 ;
 end
 always @ (posedge ) begin
    lo1406 <= li1406 ;
 end
 always @ (posedge ) begin
    lo1407 <= li1407 ;
 end
 always @ (posedge ) begin
    lo1408 <= li1408 ;
 end
 always @ (posedge ) begin
    lo1409 <= li1409 ;
 end
 always @ (posedge ) begin
    lo1410 <= li1410 ;
 end
 always @ (posedge ) begin
    lo1411 <= li1411 ;
 end
 always @ (posedge ) begin
    lo1412 <= li1412 ;
 end
 always @ (posedge ) begin
    lo1413 <= li1413 ;
 end
 always @ (posedge ) begin
    lo1414 <= li1414 ;
 end
 always @ (posedge ) begin
    lo1415 <= li1415 ;
 end
 always @ (posedge ) begin
    lo1416 <= li1416 ;
 end
 always @ (posedge ) begin
    lo1417 <= li1417 ;
 end
 always @ (posedge ) begin
    lo1418 <= li1418 ;
 end
 always @ (posedge ) begin
    lo1419 <= li1419 ;
 end
 always @ (posedge ) begin
    lo1420 <= li1420 ;
 end
 always @ (posedge ) begin
    lo1421 <= li1421 ;
 end
 always @ (posedge ) begin
    lo1422 <= li1422 ;
 end
 always @ (posedge ) begin
    lo1423 <= li1423 ;
 end
 always @ (posedge ) begin
    lo1424 <= li1424 ;
 end
 always @ (posedge ) begin
    lo1425 <= li1425 ;
 end
 always @ (posedge ) begin
    lo1426 <= li1426 ;
 end
 always @ (posedge ) begin
    lo1427 <= li1427 ;
 end
 always @ (posedge ) begin
    lo1428 <= li1428 ;
 end
 always @ (posedge ) begin
    lo1429 <= li1429 ;
 end
 always @ (posedge ) begin
    lo1430 <= li1430 ;
 end
 always @ (posedge ) begin
    lo1431 <= li1431 ;
 end
 always @ (posedge ) begin
    lo1432 <= li1432 ;
 end
 always @ (posedge ) begin
    lo1433 <= li1433 ;
 end
 always @ (posedge ) begin
    lo1434 <= li1434 ;
 end
 always @ (posedge ) begin
    lo1435 <= li1435 ;
 end
 always @ (posedge ) begin
    lo1436 <= li1436 ;
 end
 always @ (posedge ) begin
    lo1437 <= li1437 ;
 end
 always @ (posedge ) begin
    lo1438 <= li1438 ;
 end
 always @ (posedge ) begin
    lo1439 <= li1439 ;
 end
 always @ (posedge ) begin
    lo1440 <= li1440 ;
 end
 always @ (posedge ) begin
    lo1441 <= li1441 ;
 end
 always @ (posedge ) begin
    lo1442 <= li1442 ;
 end
 always @ (posedge ) begin
    lo1443 <= li1443 ;
 end
 always @ (posedge ) begin
    lo1444 <= li1444 ;
 end
 always @ (posedge ) begin
    lo1445 <= li1445 ;
 end
 always @ (posedge ) begin
    lo1446 <= li1446 ;
 end
 always @ (posedge ) begin
    lo1447 <= li1447 ;
 end
 always @ (posedge ) begin
    lo1448 <= li1448 ;
 end
 always @ (posedge ) begin
    lo1449 <= li1449 ;
 end
 always @ (posedge ) begin
    lo1450 <= li1450 ;
 end
 always @ (posedge ) begin
    lo1451 <= li1451 ;
 end
 always @ (posedge ) begin
    lo1452 <= li1452 ;
 end
 always @ (posedge ) begin
    lo1453 <= li1453 ;
 end
 always @ (posedge ) begin
    lo1454 <= li1454 ;
 end
 always @ (posedge ) begin
    lo1455 <= li1455 ;
 end
 always @ (posedge ) begin
    lo1456 <= li1456 ;
 end
 always @ (posedge ) begin
    lo1457 <= li1457 ;
 end
 always @ (posedge ) begin
    lo1458 <= li1458 ;
 end
 always @ (posedge ) begin
    lo1459 <= li1459 ;
 end
 always @ (posedge ) begin
    lo1460 <= li1460 ;
 end
 always @ (posedge ) begin
    lo1461 <= li1461 ;
 end
 always @ (posedge ) begin
    lo1462 <= li1462 ;
 end
 always @ (posedge ) begin
    lo1463 <= li1463 ;
 end
 always @ (posedge ) begin
    lo1464 <= li1464 ;
 end
 always @ (posedge ) begin
    lo1465 <= li1465 ;
 end
 always @ (posedge ) begin
    lo1466 <= li1466 ;
 end
 always @ (posedge ) begin
    lo1467 <= li1467 ;
 end
 always @ (posedge ) begin
    lo1468 <= li1468 ;
 end
 always @ (posedge ) begin
    lo1469 <= li1469 ;
 end
 always @ (posedge ) begin
    lo1470 <= li1470 ;
 end
 always @ (posedge ) begin
    lo1471 <= li1471 ;
 end
 always @ (posedge ) begin
    lo1472 <= li1472 ;
 end
 always @ (posedge ) begin
    lo1473 <= li1473 ;
 end
 always @ (posedge ) begin
    lo1474 <= li1474 ;
 end
 always @ (posedge ) begin
    lo1475 <= li1475 ;
 end
 always @ (posedge ) begin
    lo1476 <= li1476 ;
 end
 initial begin
    lo0000 <= 1'b0;
    lo0001 <= 1'b0;
    lo0002 <= 1'b0;
    lo0003 <= 1'b0;
    lo0004 <= 1'b0;
    lo0005 <= 1'b0;
    lo0006 <= 1'b0;
    lo0007 <= 1'b0;
    lo0008 <= 1'b0;
    lo0009 <= 1'b0;
    lo0010 <= 1'b0;
    lo0011 <= 1'b0;
    lo0012 <= 1'b0;
    lo0013 <= 1'b0;
    lo0014 <= 1'b0;
    lo0015 <= 1'b0;
    lo0016 <= 1'b0;
    lo0017 <= 1'b0;
    lo0018 <= 1'b0;
    lo0019 <= 1'b0;
    lo0020 <= 1'b0;
    lo0021 <= 1'b0;
    lo0022 <= 1'b0;
    lo0023 <= 1'b0;
    lo0024 <= 1'b0;
    lo0025 <= 1'b0;
    lo0026 <= 1'b0;
    lo0027 <= 1'b0;
    lo0028 <= 1'b0;
    lo0029 <= 1'b0;
    lo0030 <= 1'b0;
    lo0031 <= 1'b0;
    lo0032 <= 1'b0;
    lo0033 <= 1'b0;
    lo0034 <= 1'b0;
    lo0035 <= 1'b0;
    lo0036 <= 1'b0;
    lo0037 <= 1'b0;
    lo0038 <= 1'b0;
    lo0039 <= 1'b0;
    lo0040 <= 1'b0;
    lo0041 <= 1'b0;
    lo0042 <= 1'b0;
    lo0043 <= 1'b0;
    lo0044 <= 1'b0;
    lo0045 <= 1'b0;
    lo0046 <= 1'b0;
    lo0047 <= 1'b0;
    lo0048 <= 1'b0;
    lo0049 <= 1'b0;
    lo0050 <= 1'b0;
    lo0051 <= 1'b0;
    lo0052 <= 1'b0;
    lo0053 <= 1'b0;
    lo0054 <= 1'b0;
    lo0055 <= 1'b0;
    lo0056 <= 1'b0;
    lo0057 <= 1'b0;
    lo0058 <= 1'b0;
    lo0059 <= 1'b0;
    lo0060 <= 1'b0;
    lo0061 <= 1'b0;
    lo0062 <= 1'b0;
    lo0063 <= 1'b0;
    lo0064 <= 1'b0;
    lo0065 <= 1'b0;
    lo0066 <= 1'b0;
    lo0067 <= 1'b0;
    lo0068 <= 1'b0;
    lo0069 <= 1'b0;
    lo0070 <= 1'b0;
    lo0071 <= 1'b0;
    lo0072 <= 1'b0;
    lo0073 <= 1'b0;
    lo0074 <= 1'b0;
    lo0075 <= 1'b0;
    lo0076 <= 1'b0;
    lo0077 <= 1'b0;
    lo0078 <= 1'b0;
    lo0079 <= 1'b0;
    lo0080 <= 1'b0;
    lo0081 <= 1'b0;
    lo0082 <= 1'b0;
    lo0083 <= 1'b0;
    lo0084 <= 1'b0;
    lo0085 <= 1'b0;
    lo0086 <= 1'b0;
    lo0087 <= 1'b0;
    lo0088 <= 1'b0;
    lo0089 <= 1'b0;
    lo0090 <= 1'b0;
    lo0091 <= 1'b0;
    lo0092 <= 1'b0;
    lo0093 <= 1'b0;
    lo0094 <= 1'b0;
    lo0095 <= 1'b0;
    lo0096 <= 1'b0;
    lo0097 <= 1'b0;
    lo0098 <= 1'b0;
    lo0099 <= 1'b0;
    lo0100 <= 1'b0;
    lo0101 <= 1'b0;
    lo0102 <= 1'b0;
    lo0103 <= 1'b0;
    lo0104 <= 1'b0;
    lo0105 <= 1'b0;
    lo0106 <= 1'b0;
    lo0107 <= 1'b0;
    lo0108 <= 1'b0;
    lo0109 <= 1'b0;
    lo0110 <= 1'b0;
    lo0111 <= 1'b0;
    lo0112 <= 1'b0;
    lo0113 <= 1'b0;
    lo0114 <= 1'b0;
    lo0115 <= 1'b0;
    lo0116 <= 1'b0;
    lo0117 <= 1'b0;
    lo0118 <= 1'b0;
    lo0119 <= 1'b0;
    lo0120 <= 1'b0;
    lo0121 <= 1'b0;
    lo0122 <= 1'b0;
    lo0123 <= 1'b0;
    lo0124 <= 1'b0;
    lo0125 <= 1'b0;
    lo0126 <= 1'b0;
    lo0127 <= 1'b0;
    lo0128 <= 1'b0;
    lo0129 <= 1'b0;
    lo0130 <= 1'b0;
    lo0131 <= 1'b0;
    lo0132 <= 1'b0;
    lo0133 <= 1'b0;
    lo0134 <= 1'b0;
    lo0135 <= 1'b0;
    lo0136 <= 1'b0;
    lo0137 <= 1'b0;
    lo0138 <= 1'b0;
    lo0139 <= 1'b0;
    lo0140 <= 1'b0;
    lo0141 <= 1'b0;
    lo0142 <= 1'b0;
    lo0143 <= 1'b0;
    lo0144 <= 1'b0;
    lo0145 <= 1'b0;
    lo0146 <= 1'b0;
    lo0147 <= 1'b0;
    lo0148 <= 1'b0;
    lo0149 <= 1'b0;
    lo0150 <= 1'b0;
    lo0151 <= 1'b0;
    lo0152 <= 1'b0;
    lo0153 <= 1'b0;
    lo0154 <= 1'b0;
    lo0155 <= 1'b0;
    lo0156 <= 1'b0;
    lo0157 <= 1'b0;
    lo0158 <= 1'b0;
    lo0159 <= 1'b0;
    lo0160 <= 1'b0;
    lo0161 <= 1'b0;
    lo0162 <= 1'b0;
    lo0163 <= 1'b0;
    lo0164 <= 1'b0;
    lo0165 <= 1'b0;
    lo0166 <= 1'b0;
    lo0167 <= 1'b0;
    lo0168 <= 1'b0;
    lo0169 <= 1'b0;
    lo0170 <= 1'b0;
    lo0171 <= 1'b0;
    lo0172 <= 1'b0;
    lo0173 <= 1'b0;
    lo0174 <= 1'b0;
    lo0175 <= 1'b0;
    lo0176 <= 1'b0;
    lo0177 <= 1'b0;
    lo0178 <= 1'b0;
    lo0179 <= 1'b0;
    lo0180 <= 1'b0;
    lo0181 <= 1'b0;
    lo0182 <= 1'b0;
    lo0183 <= 1'b0;
    lo0184 <= 1'b0;
    lo0185 <= 1'b0;
    lo0186 <= 1'b0;
    lo0187 <= 1'b0;
    lo0188 <= 1'b0;
    lo0189 <= 1'b0;
    lo0190 <= 1'b0;
    lo0191 <= 1'b0;
    lo0192 <= 1'b0;
    lo0193 <= 1'b0;
    lo0194 <= 1'b0;
    lo0195 <= 1'b0;
    lo0196 <= 1'b0;
    lo0197 <= 1'b0;
    lo0198 <= 1'b0;
    lo0199 <= 1'b0;
    lo0200 <= 1'b0;
    lo0201 <= 1'b0;
    lo0202 <= 1'b0;
    lo0203 <= 1'b0;
    lo0204 <= 1'b0;
    lo0205 <= 1'b0;
    lo0206 <= 1'b0;
    lo0207 <= 1'b0;
    lo0208 <= 1'b0;
    lo0209 <= 1'b0;
    lo0210 <= 1'b0;
    lo0211 <= 1'b0;
    lo0212 <= 1'b0;
    lo0213 <= 1'b0;
    lo0214 <= 1'b0;
    lo0215 <= 1'b0;
    lo0216 <= 1'b0;
    lo0217 <= 1'b0;
    lo0218 <= 1'b0;
    lo0219 <= 1'b0;
    lo0220 <= 1'b0;
    lo0221 <= 1'b0;
    lo0222 <= 1'b0;
    lo0223 <= 1'b0;
    lo0224 <= 1'b0;
    lo0225 <= 1'b0;
    lo0226 <= 1'b0;
    lo0227 <= 1'b0;
    lo0228 <= 1'b0;
    lo0229 <= 1'b0;
    lo0230 <= 1'b0;
    lo0231 <= 1'b0;
    lo0232 <= 1'b0;
    lo0233 <= 1'b0;
    lo0234 <= 1'b0;
    lo0235 <= 1'b0;
    lo0236 <= 1'b0;
    lo0237 <= 1'b0;
    lo0238 <= 1'b0;
    lo0239 <= 1'b0;
    lo0240 <= 1'b0;
    lo0241 <= 1'b0;
    lo0242 <= 1'b0;
    lo0243 <= 1'b0;
    lo0244 <= 1'b0;
    lo0245 <= 1'b0;
    lo0246 <= 1'b0;
    lo0247 <= 1'b0;
    lo0248 <= 1'b0;
    lo0249 <= 1'b0;
    lo0250 <= 1'b0;
    lo0251 <= 1'b0;
    lo0252 <= 1'b0;
    lo0253 <= 1'b0;
    lo0254 <= 1'b0;
    lo0255 <= 1'b0;
    lo0256 <= 1'b0;
    lo0257 <= 1'b0;
    lo0258 <= 1'b0;
    lo0259 <= 1'b0;
    lo0260 <= 1'b0;
    lo0261 <= 1'b0;
    lo0262 <= 1'b0;
    lo0263 <= 1'b0;
    lo0264 <= 1'b0;
    lo0265 <= 1'b0;
    lo0266 <= 1'b0;
    lo0267 <= 1'b0;
    lo0268 <= 1'b0;
    lo0269 <= 1'b0;
    lo0270 <= 1'b0;
    lo0271 <= 1'b0;
    lo0272 <= 1'b0;
    lo0273 <= 1'b0;
    lo0274 <= 1'b0;
    lo0275 <= 1'b0;
    lo0276 <= 1'b0;
    lo0277 <= 1'b0;
    lo0278 <= 1'b0;
    lo0279 <= 1'b0;
    lo0280 <= 1'b0;
    lo0281 <= 1'b0;
    lo0282 <= 1'b0;
    lo0283 <= 1'b0;
    lo0284 <= 1'b0;
    lo0285 <= 1'b0;
    lo0286 <= 1'b0;
    lo0287 <= 1'b0;
    lo0288 <= 1'b0;
    lo0289 <= 1'b0;
    lo0290 <= 1'b0;
    lo0291 <= 1'b0;
    lo0292 <= 1'b0;
    lo0293 <= 1'b0;
    lo0294 <= 1'b0;
    lo0295 <= 1'b0;
    lo0296 <= 1'b0;
    lo0297 <= 1'b0;
    lo0298 <= 1'b0;
    lo0299 <= 1'b0;
    lo0300 <= 1'b0;
    lo0301 <= 1'b0;
    lo0302 <= 1'b0;
    lo0303 <= 1'b0;
    lo0304 <= 1'b0;
    lo0305 <= 1'b0;
    lo0306 <= 1'b0;
    lo0307 <= 1'b0;
    lo0308 <= 1'b0;
    lo0309 <= 1'b0;
    lo0310 <= 1'b0;
    lo0311 <= 1'b0;
    lo0312 <= 1'b0;
    lo0313 <= 1'b0;
    lo0314 <= 1'b0;
    lo0315 <= 1'b0;
    lo0316 <= 1'b0;
    lo0317 <= 1'b0;
    lo0318 <= 1'b0;
    lo0319 <= 1'b0;
    lo0320 <= 1'b0;
    lo0321 <= 1'b0;
    lo0322 <= 1'b0;
    lo0323 <= 1'b0;
    lo0324 <= 1'b0;
    lo0325 <= 1'b0;
    lo0326 <= 1'b0;
    lo0327 <= 1'b0;
    lo0328 <= 1'b0;
    lo0329 <= 1'b0;
    lo0330 <= 1'b0;
    lo0331 <= 1'b0;
    lo0332 <= 1'b0;
    lo0333 <= 1'b0;
    lo0334 <= 1'b0;
    lo0335 <= 1'b0;
    lo0336 <= 1'b0;
    lo0337 <= 1'b0;
    lo0338 <= 1'b0;
    lo0339 <= 1'b0;
    lo0340 <= 1'b0;
    lo0341 <= 1'b0;
    lo0342 <= 1'b0;
    lo0343 <= 1'b0;
    lo0344 <= 1'b0;
    lo0345 <= 1'b0;
    lo0346 <= 1'b0;
    lo0347 <= 1'b0;
    lo0348 <= 1'b0;
    lo0349 <= 1'b0;
    lo0350 <= 1'b0;
    lo0351 <= 1'b0;
    lo0352 <= 1'b0;
    lo0353 <= 1'b0;
    lo0354 <= 1'b0;
    lo0355 <= 1'b0;
    lo0356 <= 1'b0;
    lo0357 <= 1'b0;
    lo0358 <= 1'b0;
    lo0359 <= 1'b0;
    lo0360 <= 1'b0;
    lo0361 <= 1'b0;
    lo0362 <= 1'b0;
    lo0363 <= 1'b0;
    lo0364 <= 1'b0;
    lo0365 <= 1'b0;
    lo0366 <= 1'b0;
    lo0367 <= 1'b0;
    lo0368 <= 1'b0;
    lo0369 <= 1'b0;
    lo0370 <= 1'b0;
    lo0371 <= 1'b0;
    lo0372 <= 1'b0;
    lo0373 <= 1'b0;
    lo0374 <= 1'b0;
    lo0375 <= 1'b0;
    lo0376 <= 1'b0;
    lo0377 <= 1'b0;
    lo0378 <= 1'b0;
    lo0379 <= 1'b0;
    lo0380 <= 1'b0;
    lo0381 <= 1'b0;
    lo0382 <= 1'b0;
    lo0383 <= 1'b0;
    lo0384 <= 1'b0;
    lo0385 <= 1'b0;
    lo0386 <= 1'b0;
    lo0387 <= 1'b0;
    lo0388 <= 1'b0;
    lo0389 <= 1'b0;
    lo0390 <= 1'b0;
    lo0391 <= 1'b0;
    lo0392 <= 1'b0;
    lo0393 <= 1'b0;
    lo0394 <= 1'b0;
    lo0395 <= 1'b0;
    lo0396 <= 1'b0;
    lo0397 <= 1'b0;
    lo0398 <= 1'b0;
    lo0399 <= 1'b0;
    lo0400 <= 1'b0;
    lo0401 <= 1'b0;
    lo0402 <= 1'b0;
    lo0403 <= 1'b0;
    lo0404 <= 1'b0;
    lo0405 <= 1'b0;
    lo0406 <= 1'b0;
    lo0407 <= 1'b0;
    lo0408 <= 1'b0;
    lo0409 <= 1'b0;
    lo0410 <= 1'b0;
    lo0411 <= 1'b0;
    lo0412 <= 1'b0;
    lo0413 <= 1'b0;
    lo0414 <= 1'b0;
    lo0415 <= 1'b0;
    lo0416 <= 1'b0;
    lo0417 <= 1'b0;
    lo0418 <= 1'b0;
    lo0419 <= 1'b0;
    lo0420 <= 1'b0;
    lo0421 <= 1'b0;
    lo0422 <= 1'b0;
    lo0423 <= 1'b0;
    lo0424 <= 1'b0;
    lo0425 <= 1'b0;
    lo0426 <= 1'b0;
    lo0427 <= 1'b0;
    lo0428 <= 1'b0;
    lo0429 <= 1'b0;
    lo0430 <= 1'b0;
    lo0431 <= 1'b0;
    lo0432 <= 1'b0;
    lo0433 <= 1'b0;
    lo0434 <= 1'b0;
    lo0435 <= 1'b0;
    lo0436 <= 1'b0;
    lo0437 <= 1'b0;
    lo0438 <= 1'b0;
    lo0439 <= 1'b0;
    lo0440 <= 1'b0;
    lo0441 <= 1'b0;
    lo0442 <= 1'b0;
    lo0443 <= 1'b0;
    lo0444 <= 1'b0;
    lo0445 <= 1'b0;
    lo0446 <= 1'b0;
    lo0447 <= 1'b0;
    lo0448 <= 1'b0;
    lo0449 <= 1'b0;
    lo0450 <= 1'b0;
    lo0451 <= 1'b0;
    lo0452 <= 1'b0;
    lo0453 <= 1'b0;
    lo0454 <= 1'b0;
    lo0455 <= 1'b0;
    lo0456 <= 1'b0;
    lo0457 <= 1'b0;
    lo0458 <= 1'b0;
    lo0459 <= 1'b0;
    lo0460 <= 1'b0;
    lo0461 <= 1'b0;
    lo0462 <= 1'b0;
    lo0463 <= 1'b0;
    lo0464 <= 1'b0;
    lo0465 <= 1'b0;
    lo0466 <= 1'b0;
    lo0467 <= 1'b0;
    lo0468 <= 1'b0;
    lo0469 <= 1'b0;
    lo0470 <= 1'b0;
    lo0471 <= 1'b0;
    lo0472 <= 1'b0;
    lo0473 <= 1'b0;
    lo0474 <= 1'b0;
    lo0475 <= 1'b0;
    lo0476 <= 1'b0;
    lo0477 <= 1'b0;
    lo0478 <= 1'b0;
    lo0479 <= 1'b0;
    lo0480 <= 1'b0;
    lo0481 <= 1'b0;
    lo0482 <= 1'b0;
    lo0483 <= 1'b0;
    lo0484 <= 1'b0;
    lo0485 <= 1'b0;
    lo0486 <= 1'b0;
    lo0487 <= 1'b0;
    lo0488 <= 1'b0;
    lo0489 <= 1'b0;
    lo0490 <= 1'b0;
    lo0491 <= 1'b0;
    lo0492 <= 1'b0;
    lo0493 <= 1'b0;
    lo0494 <= 1'b0;
    lo0495 <= 1'b0;
    lo0496 <= 1'b0;
    lo0497 <= 1'b0;
    lo0498 <= 1'b0;
    lo0499 <= 1'b0;
    lo0500 <= 1'b0;
    lo0501 <= 1'b0;
    lo0502 <= 1'b0;
    lo0503 <= 1'b0;
    lo0504 <= 1'b0;
    lo0505 <= 1'b0;
    lo0506 <= 1'b0;
    lo0507 <= 1'b0;
    lo0508 <= 1'b0;
    lo0509 <= 1'b0;
    lo0510 <= 1'b0;
    lo0511 <= 1'b0;
    lo0512 <= 1'b0;
    lo0513 <= 1'b0;
    lo0514 <= 1'b0;
    lo0515 <= 1'b0;
    lo0516 <= 1'b0;
    lo0517 <= 1'b0;
    lo0518 <= 1'b0;
    lo0519 <= 1'b0;
    lo0520 <= 1'b0;
    lo0521 <= 1'b0;
    lo0522 <= 1'b0;
    lo0523 <= 1'b0;
    lo0524 <= 1'b0;
    lo0525 <= 1'b0;
    lo0526 <= 1'b0;
    lo0527 <= 1'b0;
    lo0528 <= 1'b0;
    lo0529 <= 1'b0;
    lo0530 <= 1'b0;
    lo0531 <= 1'b0;
    lo0532 <= 1'b0;
    lo0533 <= 1'b0;
    lo0534 <= 1'b0;
    lo0535 <= 1'b0;
    lo0536 <= 1'b0;
    lo0537 <= 1'b0;
    lo0538 <= 1'b0;
    lo0539 <= 1'b0;
    lo0540 <= 1'b0;
    lo0541 <= 1'b0;
    lo0542 <= 1'b0;
    lo0543 <= 1'b0;
    lo0544 <= 1'b0;
    lo0545 <= 1'b0;
    lo0546 <= 1'b0;
    lo0547 <= 1'b0;
    lo0548 <= 1'b0;
    lo0549 <= 1'b0;
    lo0550 <= 1'b0;
    lo0551 <= 1'b0;
    lo0552 <= 1'b0;
    lo0553 <= 1'b0;
    lo0554 <= 1'b0;
    lo0555 <= 1'b0;
    lo0556 <= 1'b0;
    lo0557 <= 1'b0;
    lo0558 <= 1'b0;
    lo0559 <= 1'b0;
    lo0560 <= 1'b0;
    lo0561 <= 1'b0;
    lo0562 <= 1'b0;
    lo0563 <= 1'b0;
    lo0564 <= 1'b0;
    lo0565 <= 1'b0;
    lo0566 <= 1'b0;
    lo0567 <= 1'b0;
    lo0568 <= 1'b0;
    lo0569 <= 1'b0;
    lo0570 <= 1'b0;
    lo0571 <= 1'b0;
    lo0572 <= 1'b0;
    lo0573 <= 1'b0;
    lo0574 <= 1'b0;
    lo0575 <= 1'b0;
    lo0576 <= 1'b0;
    lo0577 <= 1'b0;
    lo0578 <= 1'b0;
    lo0579 <= 1'b0;
    lo0580 <= 1'b0;
    lo0581 <= 1'b0;
    lo0582 <= 1'b0;
    lo0583 <= 1'b0;
    lo0584 <= 1'b0;
    lo0585 <= 1'b0;
    lo0586 <= 1'b0;
    lo0587 <= 1'b0;
    lo0588 <= 1'b0;
    lo0589 <= 1'b0;
    lo0590 <= 1'b0;
    lo0591 <= 1'b0;
    lo0592 <= 1'b0;
    lo0593 <= 1'b0;
    lo0594 <= 1'b0;
    lo0595 <= 1'b0;
    lo0596 <= 1'b0;
    lo0597 <= 1'b0;
    lo0598 <= 1'b0;
    lo0599 <= 1'b0;
    lo0600 <= 1'b0;
    lo0601 <= 1'b0;
    lo0602 <= 1'b0;
    lo0603 <= 1'b0;
    lo0604 <= 1'b0;
    lo0605 <= 1'b0;
    lo0606 <= 1'b0;
    lo0607 <= 1'b0;
    lo0608 <= 1'b0;
    lo0609 <= 1'b0;
    lo0610 <= 1'b0;
    lo0611 <= 1'b0;
    lo0612 <= 1'b0;
    lo0613 <= 1'b0;
    lo0614 <= 1'b0;
    lo0615 <= 1'b0;
    lo0616 <= 1'b0;
    lo0617 <= 1'b0;
    lo0618 <= 1'b0;
    lo0619 <= 1'b0;
    lo0620 <= 1'b0;
    lo0621 <= 1'b0;
    lo0622 <= 1'b0;
    lo0623 <= 1'b0;
    lo0624 <= 1'b0;
    lo0625 <= 1'b0;
    lo0626 <= 1'b0;
    lo0627 <= 1'b0;
    lo0628 <= 1'b0;
    lo0629 <= 1'b0;
    lo0630 <= 1'b0;
    lo0631 <= 1'b0;
    lo0632 <= 1'b0;
    lo0633 <= 1'b0;
    lo0634 <= 1'b0;
    lo0635 <= 1'b0;
    lo0636 <= 1'b0;
    lo0637 <= 1'b0;
    lo0638 <= 1'b0;
    lo0639 <= 1'b0;
    lo0640 <= 1'b0;
    lo0641 <= 1'b0;
    lo0642 <= 1'b0;
    lo0643 <= 1'b0;
    lo0644 <= 1'b0;
    lo0645 <= 1'b0;
    lo0646 <= 1'b0;
    lo0647 <= 1'b0;
    lo0648 <= 1'b0;
    lo0649 <= 1'b0;
    lo0650 <= 1'b0;
    lo0651 <= 1'b0;
    lo0652 <= 1'b0;
    lo0653 <= 1'b0;
    lo0654 <= 1'b0;
    lo0655 <= 1'b0;
    lo0656 <= 1'b0;
    lo0657 <= 1'b0;
    lo0658 <= 1'b0;
    lo0659 <= 1'b0;
    lo0660 <= 1'b0;
    lo0661 <= 1'b0;
    lo0662 <= 1'b0;
    lo0663 <= 1'b0;
    lo0664 <= 1'b0;
    lo0665 <= 1'b0;
    lo0666 <= 1'b0;
    lo0667 <= 1'b0;
    lo0668 <= 1'b0;
    lo0669 <= 1'b0;
    lo0670 <= 1'b0;
    lo0671 <= 1'b0;
    lo0672 <= 1'b0;
    lo0673 <= 1'b0;
    lo0674 <= 1'b0;
    lo0675 <= 1'b0;
    lo0676 <= 1'b0;
    lo0677 <= 1'b0;
    lo0678 <= 1'b0;
    lo0679 <= 1'b0;
    lo0680 <= 1'b0;
    lo0681 <= 1'b0;
    lo0682 <= 1'b0;
    lo0683 <= 1'b0;
    lo0684 <= 1'b0;
    lo0685 <= 1'b0;
    lo0686 <= 1'b0;
    lo0687 <= 1'b0;
    lo0688 <= 1'b0;
    lo0689 <= 1'b0;
    lo0690 <= 1'b0;
    lo0691 <= 1'b0;
    lo0692 <= 1'b0;
    lo0693 <= 1'b0;
    lo0694 <= 1'b0;
    lo0695 <= 1'b0;
    lo0696 <= 1'b0;
    lo0697 <= 1'b0;
    lo0698 <= 1'b0;
    lo0699 <= 1'b0;
    lo0700 <= 1'b0;
    lo0701 <= 1'b0;
    lo0702 <= 1'b0;
    lo0703 <= 1'b0;
    lo0704 <= 1'b0;
    lo0705 <= 1'b0;
    lo0706 <= 1'b0;
    lo0707 <= 1'b0;
    lo0708 <= 1'b0;
    lo0709 <= 1'b0;
    lo0710 <= 1'b0;
    lo0711 <= 1'b0;
    lo0712 <= 1'b0;
    lo0713 <= 1'b0;
    lo0714 <= 1'b0;
    lo0715 <= 1'b0;
    lo0716 <= 1'b0;
    lo0717 <= 1'b0;
    lo0718 <= 1'b0;
    lo0719 <= 1'b0;
    lo0720 <= 1'b0;
    lo0721 <= 1'b0;
    lo0722 <= 1'b0;
    lo0723 <= 1'b0;
    lo0724 <= 1'b0;
    lo0725 <= 1'b0;
    lo0726 <= 1'b0;
    lo0727 <= 1'b0;
    lo0728 <= 1'b0;
    lo0729 <= 1'b0;
    lo0730 <= 1'b0;
    lo0731 <= 1'b0;
    lo0732 <= 1'b0;
    lo0733 <= 1'b0;
    lo0734 <= 1'b0;
    lo0735 <= 1'b0;
    lo0736 <= 1'b0;
    lo0737 <= 1'b0;
    lo0738 <= 1'b0;
    lo0739 <= 1'b0;
    lo0740 <= 1'b0;
    lo0741 <= 1'b0;
    lo0742 <= 1'b0;
    lo0743 <= 1'b0;
    lo0744 <= 1'b0;
    lo0745 <= 1'b0;
    lo0746 <= 1'b0;
    lo0747 <= 1'b0;
    lo0748 <= 1'b0;
    lo0749 <= 1'b0;
    lo0750 <= 1'b0;
    lo0751 <= 1'b0;
    lo0752 <= 1'b0;
    lo0753 <= 1'b0;
    lo0754 <= 1'b0;
    lo0755 <= 1'b0;
    lo0756 <= 1'b0;
    lo0757 <= 1'b0;
    lo0758 <= 1'b0;
    lo0759 <= 1'b0;
    lo0760 <= 1'b0;
    lo0761 <= 1'b0;
    lo0762 <= 1'b0;
    lo0763 <= 1'b0;
    lo0764 <= 1'b0;
    lo0765 <= 1'b0;
    lo0766 <= 1'b0;
    lo0767 <= 1'b0;
    lo0768 <= 1'b0;
    lo0769 <= 1'b0;
    lo0770 <= 1'b0;
    lo0771 <= 1'b0;
    lo0772 <= 1'b0;
    lo0773 <= 1'b0;
    lo0774 <= 1'b0;
    lo0775 <= 1'b0;
    lo0776 <= 1'b0;
    lo0777 <= 1'b0;
    lo0778 <= 1'b0;
    lo0779 <= 1'b0;
    lo0780 <= 1'b0;
    lo0781 <= 1'b0;
    lo0782 <= 1'b0;
    lo0783 <= 1'b0;
    lo0784 <= 1'b0;
    lo0785 <= 1'b0;
    lo0786 <= 1'b0;
    lo0787 <= 1'b0;
    lo0788 <= 1'b0;
    lo0789 <= 1'b0;
    lo0790 <= 1'b0;
    lo0791 <= 1'b0;
    lo0792 <= 1'b0;
    lo0793 <= 1'b0;
    lo0794 <= 1'b0;
    lo0795 <= 1'b0;
    lo0796 <= 1'b0;
    lo0797 <= 1'b0;
    lo0798 <= 1'b0;
    lo0799 <= 1'b0;
    lo0800 <= 1'b0;
    lo0801 <= 1'b0;
    lo0802 <= 1'b0;
    lo0803 <= 1'b0;
    lo0804 <= 1'b0;
    lo0805 <= 1'b0;
    lo0806 <= 1'b0;
    lo0807 <= 1'b0;
    lo0808 <= 1'b0;
    lo0809 <= 1'b0;
    lo0810 <= 1'b0;
    lo0811 <= 1'b0;
    lo0812 <= 1'b0;
    lo0813 <= 1'b0;
    lo0814 <= 1'b0;
    lo0815 <= 1'b0;
    lo0816 <= 1'b0;
    lo0817 <= 1'b0;
    lo0818 <= 1'b0;
    lo0819 <= 1'b0;
    lo0820 <= 1'b0;
    lo0821 <= 1'b0;
    lo0822 <= 1'b0;
    lo0823 <= 1'b0;
    lo0824 <= 1'b0;
    lo0825 <= 1'b0;
    lo0826 <= 1'b0;
    lo0827 <= 1'b0;
    lo0828 <= 1'b0;
    lo0829 <= 1'b0;
    lo0830 <= 1'b0;
    lo0831 <= 1'b0;
    lo0832 <= 1'b0;
    lo0833 <= 1'b0;
    lo0834 <= 1'b0;
    lo0835 <= 1'b0;
    lo0836 <= 1'b0;
    lo0837 <= 1'b0;
    lo0838 <= 1'b0;
    lo0839 <= 1'b0;
    lo0840 <= 1'b0;
    lo0841 <= 1'b0;
    lo0842 <= 1'b0;
    lo0843 <= 1'b0;
    lo0844 <= 1'b0;
    lo0845 <= 1'b0;
    lo0846 <= 1'b0;
    lo0847 <= 1'b0;
    lo0848 <= 1'b0;
    lo0849 <= 1'b0;
    lo0850 <= 1'b0;
    lo0851 <= 1'b0;
    lo0852 <= 1'b0;
    lo0853 <= 1'b0;
    lo0854 <= 1'b0;
    lo0855 <= 1'b0;
    lo0856 <= 1'b0;
    lo0857 <= 1'b0;
    lo0858 <= 1'b0;
    lo0859 <= 1'b0;
    lo0860 <= 1'b0;
    lo0861 <= 1'b0;
    lo0862 <= 1'b0;
    lo0863 <= 1'b0;
    lo0864 <= 1'b0;
    lo0865 <= 1'b0;
    lo0866 <= 1'b0;
    lo0867 <= 1'b0;
    lo0868 <= 1'b0;
    lo0869 <= 1'b0;
    lo0870 <= 1'b0;
    lo0871 <= 1'b0;
    lo0872 <= 1'b0;
    lo0873 <= 1'b0;
    lo0874 <= 1'b0;
    lo0875 <= 1'b0;
    lo0876 <= 1'b0;
    lo0877 <= 1'b0;
    lo0878 <= 1'b0;
    lo0879 <= 1'b0;
    lo0880 <= 1'b0;
    lo0881 <= 1'b0;
    lo0882 <= 1'b0;
    lo0883 <= 1'b0;
    lo0884 <= 1'b0;
    lo0885 <= 1'b0;
    lo0886 <= 1'b0;
    lo0887 <= 1'b0;
    lo0888 <= 1'b0;
    lo0889 <= 1'b0;
    lo0890 <= 1'b0;
    lo0891 <= 1'b0;
    lo0892 <= 1'b0;
    lo0893 <= 1'b0;
    lo0894 <= 1'b0;
    lo0895 <= 1'b0;
    lo0896 <= 1'b0;
    lo0897 <= 1'b0;
    lo0898 <= 1'b0;
    lo0899 <= 1'b0;
    lo0900 <= 1'b0;
    lo0901 <= 1'b0;
    lo0902 <= 1'b0;
    lo0903 <= 1'b0;
    lo0904 <= 1'b0;
    lo0905 <= 1'b0;
    lo0906 <= 1'b0;
    lo0907 <= 1'b0;
    lo0908 <= 1'b0;
    lo0909 <= 1'b0;
    lo0910 <= 1'b0;
    lo0911 <= 1'b0;
    lo0912 <= 1'b0;
    lo0913 <= 1'b0;
    lo0914 <= 1'b0;
    lo0915 <= 1'b0;
    lo0916 <= 1'b0;
    lo0917 <= 1'b0;
    lo0918 <= 1'b0;
    lo0919 <= 1'b0;
    lo0920 <= 1'b0;
    lo0921 <= 1'b0;
    lo0922 <= 1'b0;
    lo0923 <= 1'b0;
    lo0924 <= 1'b0;
    lo0925 <= 1'b0;
    lo0926 <= 1'b0;
    lo0927 <= 1'b0;
    lo0928 <= 1'b0;
    lo0929 <= 1'b0;
    lo0930 <= 1'b0;
    lo0931 <= 1'b0;
    lo0932 <= 1'b0;
    lo0933 <= 1'b0;
    lo0934 <= 1'b0;
    lo0935 <= 1'b0;
    lo0936 <= 1'b0;
    lo0937 <= 1'b0;
    lo0938 <= 1'b0;
    lo0939 <= 1'b0;
    lo0940 <= 1'b0;
    lo0941 <= 1'b0;
    lo0942 <= 1'b0;
    lo0943 <= 1'b0;
    lo0944 <= 1'b0;
    lo0945 <= 1'b0;
    lo0946 <= 1'b0;
    lo0947 <= 1'b0;
    lo0948 <= 1'b0;
    lo0949 <= 1'b0;
    lo0950 <= 1'b0;
    lo0951 <= 1'b0;
    lo0952 <= 1'b0;
    lo0953 <= 1'b0;
    lo0954 <= 1'b0;
    lo0955 <= 1'b0;
    lo0956 <= 1'b0;
    lo0957 <= 1'b0;
    lo0958 <= 1'b0;
    lo0959 <= 1'b0;
    lo0960 <= 1'b0;
    lo0961 <= 1'b0;
    lo0962 <= 1'b0;
    lo0963 <= 1'b0;
    lo0964 <= 1'b0;
    lo0965 <= 1'b0;
    lo0966 <= 1'b0;
    lo0967 <= 1'b0;
    lo0968 <= 1'b0;
    lo0969 <= 1'b0;
    lo0970 <= 1'b0;
    lo0971 <= 1'b0;
    lo0972 <= 1'b0;
    lo0973 <= 1'b0;
    lo0974 <= 1'b0;
    lo0975 <= 1'b0;
    lo0976 <= 1'b0;
    lo0977 <= 1'b0;
    lo0978 <= 1'b0;
    lo0979 <= 1'b0;
    lo0980 <= 1'b0;
    lo0981 <= 1'b0;
    lo0982 <= 1'b0;
    lo0983 <= 1'b0;
    lo0984 <= 1'b0;
    lo0985 <= 1'b0;
    lo0986 <= 1'b0;
    lo0987 <= 1'b0;
    lo0988 <= 1'b0;
    lo0989 <= 1'b0;
    lo0990 <= 1'b0;
    lo0991 <= 1'b0;
    lo0992 <= 1'b0;
    lo0993 <= 1'b0;
    lo0994 <= 1'b0;
    lo0995 <= 1'b0;
    lo0996 <= 1'b0;
    lo0997 <= 1'b0;
    lo0998 <= 1'b0;
    lo0999 <= 1'b0;
    lo1000 <= 1'b0;
    lo1001 <= 1'b0;
    lo1002 <= 1'b0;
    lo1003 <= 1'b0;
    lo1004 <= 1'b0;
    lo1005 <= 1'b0;
    lo1006 <= 1'b0;
    lo1007 <= 1'b0;
    lo1008 <= 1'b0;
    lo1009 <= 1'b0;
    lo1010 <= 1'b0;
    lo1011 <= 1'b0;
    lo1012 <= 1'b0;
    lo1013 <= 1'b0;
    lo1014 <= 1'b0;
    lo1015 <= 1'b0;
    lo1016 <= 1'b0;
    lo1017 <= 1'b0;
    lo1018 <= 1'b0;
    lo1019 <= 1'b0;
    lo1020 <= 1'b0;
    lo1021 <= 1'b0;
    lo1022 <= 1'b0;
    lo1023 <= 1'b0;
    lo1024 <= 1'b0;
    lo1025 <= 1'b0;
    lo1026 <= 1'b0;
    lo1027 <= 1'b0;
    lo1028 <= 1'b0;
    lo1029 <= 1'b0;
    lo1030 <= 1'b0;
    lo1031 <= 1'b0;
    lo1032 <= 1'b0;
    lo1033 <= 1'b0;
    lo1034 <= 1'b0;
    lo1035 <= 1'b0;
    lo1036 <= 1'b0;
    lo1037 <= 1'b0;
    lo1038 <= 1'b0;
    lo1039 <= 1'b0;
    lo1040 <= 1'b0;
    lo1041 <= 1'b0;
    lo1042 <= 1'b0;
    lo1043 <= 1'b0;
    lo1044 <= 1'b0;
    lo1045 <= 1'b0;
    lo1046 <= 1'b0;
    lo1047 <= 1'b0;
    lo1048 <= 1'b0;
    lo1049 <= 1'b0;
    lo1050 <= 1'b0;
    lo1051 <= 1'b0;
    lo1052 <= 1'b0;
    lo1053 <= 1'b0;
    lo1054 <= 1'b0;
    lo1055 <= 1'b0;
    lo1056 <= 1'b0;
    lo1057 <= 1'b0;
    lo1058 <= 1'b0;
    lo1059 <= 1'b0;
    lo1060 <= 1'b0;
    lo1061 <= 1'b0;
    lo1062 <= 1'b0;
    lo1063 <= 1'b0;
    lo1064 <= 1'b0;
    lo1065 <= 1'b0;
    lo1066 <= 1'b0;
    lo1067 <= 1'b0;
    lo1068 <= 1'b0;
    lo1069 <= 1'b0;
    lo1070 <= 1'b0;
    lo1071 <= 1'b0;
    lo1072 <= 1'b0;
    lo1073 <= 1'b0;
    lo1074 <= 1'b0;
    lo1075 <= 1'b0;
    lo1076 <= 1'b0;
    lo1077 <= 1'b0;
    lo1078 <= 1'b0;
    lo1079 <= 1'b0;
    lo1080 <= 1'b0;
    lo1081 <= 1'b0;
    lo1082 <= 1'b0;
    lo1083 <= 1'b0;
    lo1084 <= 1'b0;
    lo1085 <= 1'b0;
    lo1086 <= 1'b0;
    lo1087 <= 1'b0;
    lo1088 <= 1'b0;
    lo1089 <= 1'b0;
    lo1090 <= 1'b0;
    lo1091 <= 1'b0;
    lo1092 <= 1'b0;
    lo1093 <= 1'b0;
    lo1094 <= 1'b0;
    lo1095 <= 1'b0;
    lo1096 <= 1'b0;
    lo1097 <= 1'b0;
    lo1098 <= 1'b0;
    lo1099 <= 1'b0;
    lo1100 <= 1'b0;
    lo1101 <= 1'b0;
    lo1102 <= 1'b0;
    lo1103 <= 1'b0;
    lo1104 <= 1'b0;
    lo1105 <= 1'b0;
    lo1106 <= 1'b0;
    lo1107 <= 1'b0;
    lo1108 <= 1'b0;
    lo1109 <= 1'b0;
    lo1110 <= 1'b0;
    lo1111 <= 1'b0;
    lo1112 <= 1'b0;
    lo1113 <= 1'b0;
    lo1114 <= 1'b0;
    lo1115 <= 1'b0;
    lo1116 <= 1'b0;
    lo1117 <= 1'b0;
    lo1118 <= 1'b0;
    lo1119 <= 1'b0;
    lo1120 <= 1'b0;
    lo1121 <= 1'b0;
    lo1122 <= 1'b0;
    lo1123 <= 1'b0;
    lo1124 <= 1'b0;
    lo1125 <= 1'b0;
    lo1126 <= 1'b0;
    lo1127 <= 1'b0;
    lo1128 <= 1'b0;
    lo1129 <= 1'b0;
    lo1130 <= 1'b0;
    lo1131 <= 1'b0;
    lo1132 <= 1'b0;
    lo1133 <= 1'b0;
    lo1134 <= 1'b0;
    lo1135 <= 1'b0;
    lo1136 <= 1'b0;
    lo1137 <= 1'b0;
    lo1138 <= 1'b0;
    lo1139 <= 1'b0;
    lo1140 <= 1'b0;
    lo1141 <= 1'b0;
    lo1142 <= 1'b0;
    lo1143 <= 1'b0;
    lo1144 <= 1'b0;
    lo1145 <= 1'b0;
    lo1146 <= 1'b0;
    lo1147 <= 1'b0;
    lo1148 <= 1'b0;
    lo1149 <= 1'b0;
    lo1150 <= 1'b0;
    lo1151 <= 1'b0;
    lo1152 <= 1'b0;
    lo1153 <= 1'b0;
    lo1154 <= 1'b0;
    lo1155 <= 1'b0;
    lo1156 <= 1'b0;
    lo1157 <= 1'b0;
    lo1158 <= 1'b0;
    lo1159 <= 1'b0;
    lo1160 <= 1'b0;
    lo1161 <= 1'b0;
    lo1162 <= 1'b0;
    lo1163 <= 1'b0;
    lo1164 <= 1'b0;
    lo1165 <= 1'b0;
    lo1166 <= 1'b0;
    lo1167 <= 1'b0;
    lo1168 <= 1'b0;
    lo1169 <= 1'b0;
    lo1170 <= 1'b0;
    lo1171 <= 1'b0;
    lo1172 <= 1'b0;
    lo1173 <= 1'b0;
    lo1174 <= 1'b0;
    lo1175 <= 1'b0;
    lo1176 <= 1'b0;
    lo1177 <= 1'b0;
    lo1178 <= 1'b0;
    lo1179 <= 1'b0;
    lo1180 <= 1'b0;
    lo1181 <= 1'b0;
    lo1182 <= 1'b0;
    lo1183 <= 1'b0;
    lo1184 <= 1'b0;
    lo1185 <= 1'b0;
    lo1186 <= 1'b0;
    lo1187 <= 1'b0;
    lo1188 <= 1'b0;
    lo1189 <= 1'b0;
    lo1190 <= 1'b0;
    lo1191 <= 1'b0;
    lo1192 <= 1'b0;
    lo1193 <= 1'b0;
    lo1194 <= 1'b0;
    lo1195 <= 1'b0;
    lo1196 <= 1'b0;
    lo1197 <= 1'b0;
    lo1198 <= 1'b0;
    lo1199 <= 1'b0;
    lo1200 <= 1'b0;
    lo1201 <= 1'b0;
    lo1202 <= 1'b0;
    lo1203 <= 1'b0;
    lo1204 <= 1'b0;
    lo1205 <= 1'b0;
    lo1206 <= 1'b0;
    lo1207 <= 1'b0;
    lo1208 <= 1'b0;
    lo1209 <= 1'b0;
    lo1210 <= 1'b0;
    lo1211 <= 1'b0;
    lo1212 <= 1'b0;
    lo1213 <= 1'b0;
    lo1214 <= 1'b0;
    lo1215 <= 1'b0;
    lo1216 <= 1'b0;
    lo1217 <= 1'b0;
    lo1218 <= 1'b0;
    lo1219 <= 1'b0;
    lo1220 <= 1'b0;
    lo1221 <= 1'b0;
    lo1222 <= 1'b0;
    lo1223 <= 1'b0;
    lo1224 <= 1'b0;
    lo1225 <= 1'b0;
    lo1226 <= 1'b0;
    lo1227 <= 1'b0;
    lo1228 <= 1'b0;
    lo1229 <= 1'b0;
    lo1230 <= 1'b0;
    lo1231 <= 1'b0;
    lo1232 <= 1'b0;
    lo1233 <= 1'b0;
    lo1234 <= 1'b0;
    lo1235 <= 1'b0;
    lo1236 <= 1'b0;
    lo1237 <= 1'b0;
    lo1238 <= 1'b0;
    lo1239 <= 1'b0;
    lo1240 <= 1'b0;
    lo1241 <= 1'b0;
    lo1242 <= 1'b0;
    lo1243 <= 1'b0;
    lo1244 <= 1'b0;
    lo1245 <= 1'b0;
    lo1246 <= 1'b0;
    lo1247 <= 1'b0;
    lo1248 <= 1'b0;
    lo1249 <= 1'b0;
    lo1250 <= 1'b0;
    lo1251 <= 1'b0;
    lo1252 <= 1'b0;
    lo1253 <= 1'b0;
    lo1254 <= 1'b0;
    lo1255 <= 1'b0;
    lo1256 <= 1'b0;
    lo1257 <= 1'b0;
    lo1258 <= 1'b0;
    lo1259 <= 1'b0;
    lo1260 <= 1'b0;
    lo1261 <= 1'b0;
    lo1262 <= 1'b0;
    lo1263 <= 1'b0;
    lo1264 <= 1'b0;
    lo1265 <= 1'b0;
    lo1266 <= 1'b0;
    lo1267 <= 1'b0;
    lo1268 <= 1'b0;
    lo1269 <= 1'b0;
    lo1270 <= 1'b0;
    lo1271 <= 1'b0;
    lo1272 <= 1'b0;
    lo1273 <= 1'b0;
    lo1274 <= 1'b0;
    lo1275 <= 1'b0;
    lo1276 <= 1'b0;
    lo1277 <= 1'b0;
    lo1278 <= 1'b0;
    lo1279 <= 1'b0;
    lo1280 <= 1'b0;
    lo1281 <= 1'b0;
    lo1282 <= 1'b0;
    lo1283 <= 1'b0;
    lo1284 <= 1'b0;
    lo1285 <= 1'b0;
    lo1286 <= 1'b0;
    lo1287 <= 1'b0;
    lo1288 <= 1'b0;
    lo1289 <= 1'b0;
    lo1290 <= 1'b0;
    lo1291 <= 1'b0;
    lo1292 <= 1'b0;
    lo1293 <= 1'b0;
    lo1294 <= 1'b0;
    lo1295 <= 1'b0;
    lo1296 <= 1'b0;
    lo1297 <= 1'b0;
    lo1298 <= 1'b0;
    lo1299 <= 1'b0;
    lo1300 <= 1'b0;
    lo1301 <= 1'b0;
    lo1302 <= 1'b0;
    lo1303 <= 1'b0;
    lo1304 <= 1'b0;
    lo1305 <= 1'b0;
    lo1306 <= 1'b0;
    lo1307 <= 1'b0;
    lo1308 <= 1'b0;
    lo1309 <= 1'b0;
    lo1310 <= 1'b0;
    lo1311 <= 1'b0;
    lo1312 <= 1'b0;
    lo1313 <= 1'b0;
    lo1314 <= 1'b0;
    lo1315 <= 1'b0;
    lo1316 <= 1'b0;
    lo1317 <= 1'b0;
    lo1318 <= 1'b0;
    lo1319 <= 1'b0;
    lo1320 <= 1'b0;
    lo1321 <= 1'b0;
    lo1322 <= 1'b0;
    lo1323 <= 1'b0;
    lo1324 <= 1'b0;
    lo1325 <= 1'b0;
    lo1326 <= 1'b0;
    lo1327 <= 1'b0;
    lo1328 <= 1'b0;
    lo1329 <= 1'b0;
    lo1330 <= 1'b0;
    lo1331 <= 1'b0;
    lo1332 <= 1'b0;
    lo1333 <= 1'b0;
    lo1334 <= 1'b0;
    lo1335 <= 1'b0;
    lo1336 <= 1'b0;
    lo1337 <= 1'b0;
    lo1338 <= 1'b0;
    lo1339 <= 1'b0;
    lo1340 <= 1'b0;
    lo1341 <= 1'b0;
    lo1342 <= 1'b0;
    lo1343 <= 1'b0;
    lo1344 <= 1'b0;
    lo1345 <= 1'b0;
    lo1346 <= 1'b0;
    lo1347 <= 1'b0;
    lo1348 <= 1'b0;
    lo1349 <= 1'b0;
    lo1350 <= 1'b0;
    lo1351 <= 1'b0;
    lo1352 <= 1'b0;
    lo1353 <= 1'b0;
    lo1354 <= 1'b0;
    lo1355 <= 1'b0;
    lo1356 <= 1'b0;
    lo1357 <= 1'b0;
    lo1358 <= 1'b0;
    lo1359 <= 1'b0;
    lo1360 <= 1'b0;
    lo1361 <= 1'b0;
    lo1362 <= 1'b0;
    lo1363 <= 1'b0;
    lo1364 <= 1'b0;
    lo1365 <= 1'b0;
    lo1366 <= 1'b0;
    lo1367 <= 1'b0;
    lo1368 <= 1'b0;
    lo1369 <= 1'b0;
    lo1370 <= 1'b0;
    lo1371 <= 1'b0;
    lo1372 <= 1'b0;
    lo1373 <= 1'b0;
    lo1374 <= 1'b0;
    lo1375 <= 1'b0;
    lo1376 <= 1'b0;
    lo1377 <= 1'b0;
    lo1378 <= 1'b0;
    lo1379 <= 1'b0;
    lo1380 <= 1'b0;
    lo1381 <= 1'b0;
    lo1382 <= 1'b0;
    lo1383 <= 1'b0;
    lo1384 <= 1'b0;
    lo1385 <= 1'b0;
    lo1386 <= 1'b0;
    lo1387 <= 1'b0;
    lo1388 <= 1'b0;
    lo1389 <= 1'b0;
    lo1390 <= 1'b0;
    lo1391 <= 1'b0;
    lo1392 <= 1'b0;
    lo1393 <= 1'b0;
    lo1394 <= 1'b0;
    lo1395 <= 1'b0;
    lo1396 <= 1'b0;
    lo1397 <= 1'b0;
    lo1398 <= 1'b0;
    lo1399 <= 1'b0;
    lo1400 <= 1'b0;
    lo1401 <= 1'b0;
    lo1402 <= 1'b0;
    lo1403 <= 1'b0;
    lo1404 <= 1'b0;
    lo1405 <= 1'b0;
    lo1406 <= 1'b0;
    lo1407 <= 1'b0;
    lo1408 <= 1'b0;
    lo1409 <= 1'b0;
    lo1410 <= 1'b0;
    lo1411 <= 1'b0;
    lo1412 <= 1'b0;
    lo1413 <= 1'b0;
    lo1414 <= 1'b0;
    lo1415 <= 1'b0;
    lo1416 <= 1'b0;
    lo1417 <= 1'b0;
    lo1418 <= 1'b0;
    lo1419 <= 1'b0;
    lo1420 <= 1'b0;
    lo1421 <= 1'b0;
    lo1422 <= 1'b0;
    lo1423 <= 1'b0;
    lo1424 <= 1'b0;
    lo1425 <= 1'b0;
    lo1426 <= 1'b0;
    lo1427 <= 1'b0;
    lo1428 <= 1'b0;
    lo1429 <= 1'b0;
    lo1430 <= 1'b0;
    lo1431 <= 1'b0;
    lo1432 <= 1'b0;
    lo1433 <= 1'b0;
    lo1434 <= 1'b0;
    lo1435 <= 1'b0;
    lo1436 <= 1'b0;
    lo1437 <= 1'b0;
    lo1438 <= 1'b0;
    lo1439 <= 1'b0;
    lo1440 <= 1'b0;
    lo1441 <= 1'b0;
    lo1442 <= 1'b0;
    lo1443 <= 1'b0;
    lo1444 <= 1'b0;
    lo1445 <= 1'b0;
    lo1446 <= 1'b0;
    lo1447 <= 1'b0;
    lo1448 <= 1'b0;
    lo1449 <= 1'b0;
    lo1450 <= 1'b0;
    lo1451 <= 1'b0;
    lo1452 <= 1'b0;
    lo1453 <= 1'b0;
    lo1454 <= 1'b0;
    lo1455 <= 1'b0;
    lo1456 <= 1'b0;
    lo1457 <= 1'b0;
    lo1458 <= 1'b0;
    lo1459 <= 1'b0;
    lo1460 <= 1'b0;
    lo1461 <= 1'b0;
    lo1462 <= 1'b0;
    lo1463 <= 1'b0;
    lo1464 <= 1'b0;
    lo1465 <= 1'b0;
    lo1466 <= 1'b0;
    lo1467 <= 1'b0;
    lo1468 <= 1'b0;
    lo1469 <= 1'b0;
    lo1470 <= 1'b0;
    lo1471 <= 1'b0;
    lo1472 <= 1'b0;
    lo1473 <= 1'b0;
    lo1474 <= 1'b0;
    lo1475 <= 1'b0;
    lo1476 <= 1'b0;
 end
endmodule
